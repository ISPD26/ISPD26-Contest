module aes_cipher_top (SE,
    clk,
    done,
    ld,
    rst,
    key,
    text_in,
    text_out);
 input SE;
 input clk;
 output done;
 input ld;
 input rst;
 input [127:0] key;
 input [127:0] text_in;
 output [127:0] text_out;

 wire net259;
 wire n100;
 wire n1000;
 wire n1001;
 wire n1002;
 wire n1003;
 wire n1004;
 wire n1005;
 wire n1006;
 wire n1007;
 wire n1008;
 wire n1009;
 wire n101;
 wire n1010;
 wire n1011;
 wire n1012;
 wire n1013;
 wire n1014;
 wire n1015;
 wire n1016;
 wire n1017;
 wire n1018;
 wire n1019;
 wire n102;
 wire n1020;
 wire n1021;
 wire n1022;
 wire n1023;
 wire n1024;
 wire n1025;
 wire n1026;
 wire n1027;
 wire n1028;
 wire n1029;
 wire n103;
 wire n1030;
 wire n1031;
 wire n1032;
 wire n1033;
 wire n1034;
 wire n1035;
 wire n1036;
 wire n1037;
 wire n1038;
 wire n1039;
 wire n104;
 wire n1040;
 wire n1041;
 wire n1042;
 wire n1043;
 wire n1044;
 wire n1045;
 wire n1046;
 wire n1047;
 wire n1048;
 wire n1049;
 wire n105;
 wire n1050;
 wire n1051;
 wire n1052;
 wire n1053;
 wire n1054;
 wire n1055;
 wire n1056;
 wire n1057;
 wire n1058;
 wire n1059;
 wire n106;
 wire n1060;
 wire n1061;
 wire n1062;
 wire n1063;
 wire n1064;
 wire n1065;
 wire n1066;
 wire n1067;
 wire n1068;
 wire n1069;
 wire n107;
 wire n1070;
 wire n1071;
 wire n1072;
 wire n1073;
 wire n1074;
 wire n1075;
 wire n1076;
 wire n1077;
 wire n1078;
 wire n1079;
 wire n108;
 wire n1080;
 wire n1081;
 wire n1082;
 wire n1083;
 wire n1084;
 wire n1085;
 wire n1086;
 wire n1087;
 wire n1088;
 wire n1089;
 wire n109;
 wire n1090;
 wire n1091;
 wire n1092;
 wire n1093;
 wire n1094;
 wire n1095;
 wire n1096;
 wire n1097;
 wire n1098;
 wire n1099;
 wire n110;
 wire n1100;
 wire n1101;
 wire n1102;
 wire n1103;
 wire n1104;
 wire n1105;
 wire n1106;
 wire n1107;
 wire n1108;
 wire n1109;
 wire n111;
 wire n1110;
 wire n1111;
 wire n1112;
 wire n1113;
 wire n1114;
 wire n1115;
 wire n1116;
 wire n1117;
 wire n1118;
 wire n1119;
 wire n112;
 wire n1120;
 wire n1121;
 wire n1122;
 wire n1123;
 wire n1124;
 wire n1125;
 wire n1126;
 wire n1127;
 wire n1128;
 wire n1129;
 wire n113;
 wire n1130;
 wire n1131;
 wire n1132;
 wire n1133;
 wire n1134;
 wire n1135;
 wire n1136;
 wire n1137;
 wire n1138;
 wire n1139;
 wire n114;
 wire n1140;
 wire n1141;
 wire n1142;
 wire n1143;
 wire n1144;
 wire n1145;
 wire n1146;
 wire n1147;
 wire n1148;
 wire n1149;
 wire n115;
 wire n1150;
 wire n1151;
 wire n1152;
 wire n1153;
 wire n1154;
 wire n1155;
 wire n1156;
 wire n1157;
 wire n1158;
 wire n1159;
 wire n116;
 wire n1160;
 wire n1161;
 wire n1162;
 wire n1163;
 wire n1164;
 wire n1165;
 wire n1166;
 wire n1167;
 wire n1168;
 wire n1169;
 wire n117;
 wire n1170;
 wire n1171;
 wire n1172;
 wire n1173;
 wire n1174;
 wire n1175;
 wire n1176;
 wire n1177;
 wire n1178;
 wire n1179;
 wire n118;
 wire n1180;
 wire n1181;
 wire n1182;
 wire n1183;
 wire n1184;
 wire n1185;
 wire n1186;
 wire n1187;
 wire n1188;
 wire n1189;
 wire n119;
 wire n1190;
 wire n1191;
 wire n1192;
 wire n1193;
 wire n1194;
 wire n1195;
 wire n1196;
 wire n1197;
 wire n1198;
 wire n1199;
 wire n120;
 wire n1200;
 wire n1201;
 wire n1202;
 wire n1203;
 wire n1204;
 wire n1205;
 wire n1206;
 wire n1207;
 wire n1208;
 wire n1209;
 wire n121;
 wire n1210;
 wire n1211;
 wire n1212;
 wire n1213;
 wire n1214;
 wire n1215;
 wire n1216;
 wire n1217;
 wire n1218;
 wire n1219;
 wire n122;
 wire n1220;
 wire n1221;
 wire n1222;
 wire n1223;
 wire n1224;
 wire n1225;
 wire n1226;
 wire n1227;
 wire n1228;
 wire n1229;
 wire n123;
 wire n1230;
 wire n1231;
 wire n1232;
 wire n124;
 wire n125;
 wire n126;
 wire n127;
 wire n128;
 wire n129;
 wire n130;
 wire n131;
 wire n132;
 wire n133;
 wire n134;
 wire n135;
 wire n136;
 wire n137;
 wire n138;
 wire n139;
 wire n140;
 wire n141;
 wire n142;
 wire n143;
 wire n144;
 wire n145;
 wire n146;
 wire n147;
 wire n148;
 wire n149;
 wire n150;
 wire n151;
 wire n152;
 wire n153;
 wire n154;
 wire n155;
 wire n156;
 wire n157;
 wire n158;
 wire n159;
 wire n160;
 wire n161;
 wire n162;
 wire n163;
 wire n164;
 wire n165;
 wire n166;
 wire n167;
 wire n168;
 wire n169;
 wire n170;
 wire n171;
 wire n172;
 wire n173;
 wire n174;
 wire n175;
 wire n176;
 wire n177;
 wire n178;
 wire n179;
 wire n180;
 wire n181;
 wire n182;
 wire n183;
 wire n184;
 wire n185;
 wire n186;
 wire n187;
 wire n188;
 wire n189;
 wire n190;
 wire n191;
 wire n192;
 wire n193;
 wire n194;
 wire n195;
 wire n196;
 wire n197;
 wire n198;
 wire n199;
 wire n200;
 wire n201;
 wire n202;
 wire n203;
 wire n204;
 wire n205;
 wire n206;
 wire n207;
 wire n208;
 wire n209;
 wire n210;
 wire n211;
 wire n212;
 wire n213;
 wire n214;
 wire n215;
 wire n216;
 wire n217;
 wire n218;
 wire n219;
 wire n220;
 wire n221;
 wire n222;
 wire n223;
 wire n224;
 wire n225;
 wire n226;
 wire n227;
 wire n228;
 wire n229;
 wire n230;
 wire n231;
 wire n232;
 wire n233;
 wire n234;
 wire n235;
 wire n236;
 wire n237;
 wire n238;
 wire n239;
 wire n240;
 wire n241;
 wire n242;
 wire n243;
 wire n244;
 wire n245;
 wire n246;
 wire n247;
 wire n248;
 wire n249;
 wire n250;
 wire n251;
 wire n252;
 wire n253;
 wire n254;
 wire n255;
 wire n256;
 wire n257;
 wire n258;
 wire n259;
 wire n260;
 wire n261;
 wire n262;
 wire n263;
 wire n264;
 wire n265;
 wire n266;
 wire n267;
 wire n268;
 wire n269;
 wire n270;
 wire n271;
 wire n272;
 wire n273;
 wire n274;
 wire n275;
 wire n276;
 wire n277;
 wire n278;
 wire n279;
 wire n280;
 wire n281;
 wire n282;
 wire n283;
 wire n284;
 wire n285;
 wire n286;
 wire n287;
 wire n288;
 wire n289;
 wire n290;
 wire n291;
 wire n292;
 wire n293;
 wire n294;
 wire n295;
 wire n296;
 wire n297;
 wire n298;
 wire n299;
 wire n300;
 wire n301;
 wire n302;
 wire n303;
 wire n304;
 wire n305;
 wire n306;
 wire n307;
 wire n308;
 wire n309;
 wire n310;
 wire n311;
 wire n312;
 wire n313;
 wire n314;
 wire n315;
 wire n316;
 wire n317;
 wire n318;
 wire n319;
 wire n320;
 wire n321;
 wire n322;
 wire n323;
 wire n324;
 wire n325;
 wire n326;
 wire n327;
 wire n328;
 wire n329;
 wire n330;
 wire n331;
 wire n332;
 wire n333;
 wire n334;
 wire n335;
 wire n336;
 wire n337;
 wire n338;
 wire n339;
 wire n340;
 wire n341;
 wire n342;
 wire n343;
 wire n344;
 wire n345;
 wire n346;
 wire n347;
 wire n348;
 wire n349;
 wire n350;
 wire n351;
 wire n352;
 wire n353;
 wire n354;
 wire n355;
 wire n356;
 wire n357;
 wire n358;
 wire n359;
 wire n360;
 wire n361;
 wire n362;
 wire n363;
 wire n364;
 wire n365;
 wire n366;
 wire n367;
 wire n368;
 wire n369;
 wire n370;
 wire n371;
 wire n372;
 wire n373;
 wire n374;
 wire n375;
 wire n376;
 wire n377;
 wire n378;
 wire n379;
 wire n38;
 wire n380;
 wire n381;
 wire n382;
 wire n383;
 wire n384;
 wire n385;
 wire n386;
 wire n387;
 wire n388;
 wire n389;
 wire n39;
 wire n390;
 wire n391;
 wire n392;
 wire n393;
 wire n394;
 wire n395;
 wire n396;
 wire n397;
 wire n398;
 wire n399;
 wire n40;
 wire n400;
 wire n401;
 wire n402;
 wire n403;
 wire n404;
 wire n405;
 wire n406;
 wire n407;
 wire n408;
 wire n409;
 wire n41;
 wire n410;
 wire n411;
 wire n412;
 wire n413;
 wire n414;
 wire n415;
 wire n416;
 wire n417;
 wire n418;
 wire n419;
 wire n42;
 wire n420;
 wire n421;
 wire n422;
 wire n423;
 wire n424;
 wire n425;
 wire n426;
 wire n427;
 wire n428;
 wire n429;
 wire n43;
 wire n430;
 wire n431;
 wire n432;
 wire n433;
 wire n434;
 wire n435;
 wire n436;
 wire n437;
 wire n438;
 wire n439;
 wire n44;
 wire n440;
 wire n441;
 wire n442;
 wire n443;
 wire n444;
 wire n445;
 wire n446;
 wire n447;
 wire n448;
 wire n449;
 wire n45;
 wire n450;
 wire n451;
 wire n452;
 wire n453;
 wire n454;
 wire n455;
 wire n456;
 wire n457;
 wire n458;
 wire n459;
 wire n46;
 wire n460;
 wire n461;
 wire n462;
 wire n463;
 wire n464;
 wire n465;
 wire n466;
 wire n467;
 wire n468;
 wire n469;
 wire n47;
 wire n470;
 wire n471;
 wire n472;
 wire n473;
 wire n474;
 wire n475;
 wire n476;
 wire n477;
 wire n478;
 wire n479;
 wire n48;
 wire n480;
 wire n481;
 wire n482;
 wire n483;
 wire n484;
 wire n485;
 wire n486;
 wire n487;
 wire n488;
 wire n489;
 wire n49;
 wire n490;
 wire n491;
 wire n492;
 wire n493;
 wire n494;
 wire n495;
 wire n496;
 wire n497;
 wire n498;
 wire n499;
 wire n50;
 wire n500;
 wire n501;
 wire n502;
 wire n503;
 wire n504;
 wire n505;
 wire n506;
 wire n507;
 wire n508;
 wire n509;
 wire n51;
 wire n510;
 wire n511;
 wire n512;
 wire n513;
 wire n514;
 wire n515;
 wire n516;
 wire n517;
 wire n518;
 wire n519;
 wire n52;
 wire n520;
 wire n521;
 wire n522;
 wire n523;
 wire n524;
 wire n525;
 wire n526;
 wire n527;
 wire n528;
 wire n529;
 wire n53;
 wire n530;
 wire n531;
 wire n532;
 wire n533;
 wire n534;
 wire n535;
 wire n536;
 wire n537;
 wire n538;
 wire n539;
 wire n54;
 wire n540;
 wire n541;
 wire n542;
 wire n543;
 wire n544;
 wire n545;
 wire n546;
 wire n547;
 wire n548;
 wire n549;
 wire n55;
 wire n550;
 wire n551;
 wire n552;
 wire n553;
 wire n554;
 wire n555;
 wire n556;
 wire n557;
 wire n558;
 wire n559;
 wire n56;
 wire n560;
 wire n561;
 wire n562;
 wire n563;
 wire n564;
 wire n565;
 wire n566;
 wire n567;
 wire n568;
 wire n569;
 wire n57;
 wire n570;
 wire n571;
 wire n572;
 wire n573;
 wire n574;
 wire n575;
 wire n576;
 wire n577;
 wire n578;
 wire n579;
 wire n58;
 wire n580;
 wire n581;
 wire n582;
 wire n583;
 wire n584;
 wire n585;
 wire n586;
 wire n587;
 wire n588;
 wire n589;
 wire n59;
 wire n590;
 wire n591;
 wire n592;
 wire n593;
 wire n594;
 wire n595;
 wire n596;
 wire n597;
 wire n598;
 wire n599;
 wire n60;
 wire n600;
 wire n601;
 wire n602;
 wire n603;
 wire n604;
 wire n605;
 wire n606;
 wire n607;
 wire n608;
 wire n609;
 wire n61;
 wire n610;
 wire n611;
 wire n612;
 wire n613;
 wire n614;
 wire n615;
 wire n616;
 wire n617;
 wire n618;
 wire n619;
 wire n62;
 wire n620;
 wire n621;
 wire n622;
 wire n623;
 wire n624;
 wire n625;
 wire n626;
 wire n627;
 wire n628;
 wire n629;
 wire n63;
 wire n630;
 wire n631;
 wire n632;
 wire n633;
 wire n634;
 wire n635;
 wire n636;
 wire n637;
 wire n638;
 wire n639;
 wire n64;
 wire n640;
 wire n641;
 wire n642;
 wire n643;
 wire n644;
 wire n645;
 wire n646;
 wire n647;
 wire n648;
 wire n649;
 wire n65;
 wire n650;
 wire n651;
 wire n652;
 wire n653;
 wire n654;
 wire n655;
 wire n656;
 wire n657;
 wire n658;
 wire n659;
 wire n66;
 wire n660;
 wire n661;
 wire n662;
 wire n663;
 wire n664;
 wire n665;
 wire n666;
 wire n667;
 wire n668;
 wire n669;
 wire n67;
 wire n670;
 wire n671;
 wire n672;
 wire n673;
 wire n674;
 wire n675;
 wire n676;
 wire n677;
 wire n678;
 wire n679;
 wire n68;
 wire n680;
 wire n681;
 wire n682;
 wire n683;
 wire n684;
 wire n685;
 wire n686;
 wire n687;
 wire n688;
 wire n689;
 wire n69;
 wire n690;
 wire n691;
 wire n692;
 wire n693;
 wire n694;
 wire n695;
 wire n696;
 wire n697;
 wire n698;
 wire n699;
 wire n70;
 wire n700;
 wire n701;
 wire n702;
 wire n703;
 wire n704;
 wire n705;
 wire n706;
 wire n707;
 wire n708;
 wire n709;
 wire n71;
 wire n710;
 wire n711;
 wire n712;
 wire n713;
 wire n714;
 wire n715;
 wire n716;
 wire n717;
 wire n718;
 wire n719;
 wire n72;
 wire n720;
 wire n721;
 wire n722;
 wire n723;
 wire n724;
 wire n725;
 wire n726;
 wire n727;
 wire n728;
 wire n729;
 wire n73;
 wire n730;
 wire n731;
 wire n732;
 wire n733;
 wire n734;
 wire n735;
 wire n736;
 wire n737;
 wire n738;
 wire n739;
 wire n74;
 wire n740;
 wire n741;
 wire n742;
 wire n743;
 wire n744;
 wire n745;
 wire n746;
 wire n747;
 wire n748;
 wire n749;
 wire n75;
 wire n750;
 wire n751;
 wire n752;
 wire n753;
 wire n754;
 wire n755;
 wire n756;
 wire n757;
 wire n758;
 wire n759;
 wire n76;
 wire n760;
 wire n761;
 wire n762;
 wire n763;
 wire n764;
 wire n765;
 wire n766;
 wire n767;
 wire n768;
 wire n769;
 wire n77;
 wire n770;
 wire n771;
 wire n772;
 wire n773;
 wire n774;
 wire n775;
 wire n776;
 wire n777;
 wire n778;
 wire n779;
 wire n78;
 wire n780;
 wire n781;
 wire n782;
 wire n783;
 wire n784;
 wire n785;
 wire n786;
 wire n787;
 wire n788;
 wire n789;
 wire n79;
 wire n790;
 wire n791;
 wire n792;
 wire n793;
 wire n794;
 wire n795;
 wire n796;
 wire n797;
 wire n798;
 wire n799;
 wire n80;
 wire n800;
 wire n801;
 wire n802;
 wire n803;
 wire n804;
 wire n805;
 wire n806;
 wire n807;
 wire n808;
 wire n809;
 wire n81;
 wire n810;
 wire n811;
 wire n812;
 wire n813;
 wire n814;
 wire n815;
 wire n816;
 wire n817;
 wire n818;
 wire n819;
 wire n82;
 wire n820;
 wire n821;
 wire n822;
 wire n823;
 wire n824;
 wire n825;
 wire n826;
 wire n827;
 wire n828;
 wire n829;
 wire n83;
 wire n830;
 wire n831;
 wire n832;
 wire n833;
 wire n834;
 wire n835;
 wire n836;
 wire n837;
 wire n838;
 wire n839;
 wire n84;
 wire n840;
 wire n841;
 wire n842;
 wire n843;
 wire n844;
 wire n845;
 wire n846;
 wire n847;
 wire n848;
 wire n849;
 wire n85;
 wire n850;
 wire n851;
 wire n852;
 wire n853;
 wire n854;
 wire n855;
 wire n856;
 wire n857;
 wire n858;
 wire n859;
 wire n86;
 wire n860;
 wire n861;
 wire n862;
 wire n863;
 wire n864;
 wire n865;
 wire n866;
 wire n867;
 wire n868;
 wire n869;
 wire n87;
 wire n870;
 wire n871;
 wire n872;
 wire n873;
 wire n874;
 wire n875;
 wire n876;
 wire n877;
 wire n878;
 wire n879;
 wire n88;
 wire n880;
 wire n881;
 wire n882;
 wire n883;
 wire n884;
 wire n885;
 wire n886;
 wire n887;
 wire n888;
 wire n889;
 wire n89;
 wire n890;
 wire n891;
 wire n892;
 wire n893;
 wire n894;
 wire n895;
 wire n896;
 wire n897;
 wire n898;
 wire n899;
 wire n90;
 wire n900;
 wire n901;
 wire n902;
 wire n903;
 wire n904;
 wire n905;
 wire n906;
 wire n907;
 wire n908;
 wire n909;
 wire n91;
 wire n910;
 wire n911;
 wire n912;
 wire n913;
 wire n914;
 wire n915;
 wire n916;
 wire n917;
 wire n918;
 wire n919;
 wire n92;
 wire n920;
 wire n921;
 wire n922;
 wire n923;
 wire n924;
 wire n925;
 wire n926;
 wire n927;
 wire n928;
 wire n929;
 wire n93;
 wire n930;
 wire n931;
 wire n932;
 wire n933;
 wire n934;
 wire n935;
 wire n936;
 wire n937;
 wire n938;
 wire n939;
 wire n94;
 wire n940;
 wire n941;
 wire n942;
 wire n943;
 wire n944;
 wire n945;
 wire n946;
 wire n947;
 wire n948;
 wire n949;
 wire n95;
 wire n950;
 wire n951;
 wire n952;
 wire n953;
 wire n954;
 wire n955;
 wire n956;
 wire n957;
 wire n958;
 wire n959;
 wire n96;
 wire n960;
 wire n961;
 wire n962;
 wire n963;
 wire n964;
 wire n965;
 wire n966;
 wire n967;
 wire n968;
 wire n969;
 wire n97;
 wire n970;
 wire n971;
 wire n972;
 wire n973;
 wire n974;
 wire n975;
 wire n976;
 wire n977;
 wire n978;
 wire n979;
 wire n98;
 wire n980;
 wire n981;
 wire n982;
 wire n983;
 wire n984;
 wire n985;
 wire n986;
 wire n987;
 wire n988;
 wire n989;
 wire n99;
 wire n990;
 wire n991;
 wire n992;
 wire n993;
 wire n994;
 wire n995;
 wire n996;
 wire n997;
 wire n998;
 wire n999;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire \i43/n10 ;
 wire \i43/n100 ;
 wire \i43/n101 ;
 wire \i43/n102 ;
 wire \i43/n103 ;
 wire \i43/n104 ;
 wire \i43/n105 ;
 wire \i43/n106 ;
 wire \i43/n107 ;
 wire \i43/n108 ;
 wire \i43/n109 ;
 wire \i43/n11 ;
 wire \i43/n110 ;
 wire \i43/n111 ;
 wire \i43/n112 ;
 wire \i43/n113 ;
 wire \i43/n114 ;
 wire \i43/n115 ;
 wire \i43/n116 ;
 wire \i43/n117 ;
 wire \i43/n118 ;
 wire \i43/n119 ;
 wire \i43/n12 ;
 wire \i43/n120 ;
 wire \i43/n121 ;
 wire \i43/n122 ;
 wire \i43/n123 ;
 wire \i43/n124 ;
 wire \i43/n125 ;
 wire \i43/n126 ;
 wire \i43/n127 ;
 wire \i43/n128 ;
 wire \i43/n129 ;
 wire \i43/n13 ;
 wire \i43/n130 ;
 wire \i43/n131 ;
 wire \i43/n132 ;
 wire \i43/n133 ;
 wire \i43/n134 ;
 wire \i43/n135 ;
 wire \i43/n136 ;
 wire \i43/n137 ;
 wire \i43/n138 ;
 wire \i43/n139 ;
 wire \i43/n14 ;
 wire \i43/n140 ;
 wire \i43/n141 ;
 wire \i43/n142 ;
 wire \i43/n143 ;
 wire \i43/n144 ;
 wire \i43/n145 ;
 wire \i43/n146 ;
 wire \i43/n147 ;
 wire \i43/n148 ;
 wire \i43/n149 ;
 wire \i43/n15 ;
 wire \i43/n150 ;
 wire \i43/n151 ;
 wire \i43/n152 ;
 wire \i43/n153 ;
 wire \i43/n154 ;
 wire \i43/n155 ;
 wire \i43/n156 ;
 wire \i43/n157 ;
 wire \i43/n158 ;
 wire \i43/n159 ;
 wire \i43/n16 ;
 wire \i43/n160 ;
 wire \i43/n161 ;
 wire \i43/n162 ;
 wire \i43/n163 ;
 wire \i43/n164 ;
 wire \i43/n165 ;
 wire \i43/n166 ;
 wire \i43/n167 ;
 wire \i43/n168 ;
 wire \i43/n169 ;
 wire \i43/n17 ;
 wire \i43/n170 ;
 wire \i43/n171 ;
 wire \i43/n172 ;
 wire \i43/n173 ;
 wire \i43/n174 ;
 wire \i43/n175 ;
 wire \i43/n176 ;
 wire \i43/n177 ;
 wire \i43/n178 ;
 wire \i43/n179 ;
 wire \i43/n18 ;
 wire \i43/n180 ;
 wire \i43/n181 ;
 wire \i43/n182 ;
 wire \i43/n183 ;
 wire \i43/n184 ;
 wire \i43/n185 ;
 wire \i43/n186 ;
 wire \i43/n187 ;
 wire \i43/n188 ;
 wire \i43/n189 ;
 wire \i43/n19 ;
 wire \i43/n190 ;
 wire \i43/n191 ;
 wire \i43/n192 ;
 wire \i43/n193 ;
 wire \i43/n194 ;
 wire \i43/n195 ;
 wire \i43/n196 ;
 wire \i43/n197 ;
 wire \i43/n198 ;
 wire \i43/n199 ;
 wire \i43/n20 ;
 wire \i43/n200 ;
 wire \i43/n201 ;
 wire \i43/n202 ;
 wire \i43/n203 ;
 wire \i43/n204 ;
 wire \i43/n205 ;
 wire \i43/n206 ;
 wire \i43/n207 ;
 wire \i43/n208 ;
 wire \i43/n209 ;
 wire \i43/n21 ;
 wire \i43/n210 ;
 wire \i43/n211 ;
 wire \i43/n212 ;
 wire \i43/n213 ;
 wire \i43/n214 ;
 wire \i43/n215 ;
 wire \i43/n216 ;
 wire \i43/n217 ;
 wire \i43/n218 ;
 wire \i43/n219 ;
 wire \i43/n22 ;
 wire \i43/n220 ;
 wire \i43/n221 ;
 wire \i43/n222 ;
 wire \i43/n223 ;
 wire \i43/n224 ;
 wire \i43/n225 ;
 wire \i43/n226 ;
 wire \i43/n227 ;
 wire \i43/n228 ;
 wire \i43/n229 ;
 wire \i43/n23 ;
 wire \i43/n230 ;
 wire \i43/n231 ;
 wire \i43/n232 ;
 wire \i43/n233 ;
 wire \i43/n234 ;
 wire \i43/n235 ;
 wire \i43/n236 ;
 wire \i43/n237 ;
 wire \i43/n238 ;
 wire \i43/n239 ;
 wire \i43/n24 ;
 wire \i43/n240 ;
 wire \i43/n241 ;
 wire \i43/n242 ;
 wire \i43/n243 ;
 wire \i43/n244 ;
 wire \i43/n245 ;
 wire \i43/n246 ;
 wire \i43/n247 ;
 wire \i43/n248 ;
 wire \i43/n249 ;
 wire \i43/n25 ;
 wire \i43/n250 ;
 wire \i43/n251 ;
 wire \i43/n252 ;
 wire \i43/n253 ;
 wire \i43/n254 ;
 wire \i43/n255 ;
 wire \i43/n256 ;
 wire \i43/n257 ;
 wire \i43/n258 ;
 wire \i43/n259 ;
 wire \i43/n26 ;
 wire \i43/n260 ;
 wire \i43/n261 ;
 wire \i43/n262 ;
 wire \i43/n263 ;
 wire \i43/n264 ;
 wire \i43/n265 ;
 wire \i43/n266 ;
 wire \i43/n267 ;
 wire \i43/n268 ;
 wire \i43/n269 ;
 wire \i43/n27 ;
 wire \i43/n270 ;
 wire \i43/n271 ;
 wire \i43/n272 ;
 wire \i43/n273 ;
 wire \i43/n274 ;
 wire \i43/n275 ;
 wire \i43/n276 ;
 wire \i43/n277 ;
 wire \i43/n278 ;
 wire \i43/n279 ;
 wire \i43/n28 ;
 wire \i43/n280 ;
 wire \i43/n281 ;
 wire \i43/n282 ;
 wire \i43/n283 ;
 wire \i43/n284 ;
 wire \i43/n285 ;
 wire \i43/n286 ;
 wire \i43/n287 ;
 wire \i43/n288 ;
 wire \i43/n289 ;
 wire \i43/n29 ;
 wire \i43/n290 ;
 wire \i43/n291 ;
 wire \i43/n292 ;
 wire \i43/n293 ;
 wire \i43/n294 ;
 wire \i43/n295 ;
 wire \i43/n296 ;
 wire \i43/n297 ;
 wire \i43/n298 ;
 wire \i43/n299 ;
 wire \i43/n3 ;
 wire \i43/n30 ;
 wire \i43/n300 ;
 wire \i43/n301 ;
 wire \i43/n302 ;
 wire \i43/n303 ;
 wire \i43/n304 ;
 wire \i43/n305 ;
 wire \i43/n306 ;
 wire \i43/n307 ;
 wire \i43/n308 ;
 wire \i43/n309 ;
 wire \i43/n31 ;
 wire \i43/n310 ;
 wire \i43/n311 ;
 wire \i43/n312 ;
 wire \i43/n313 ;
 wire \i43/n314 ;
 wire \i43/n315 ;
 wire \i43/n316 ;
 wire \i43/n317 ;
 wire \i43/n318 ;
 wire \i43/n319 ;
 wire \i43/n32 ;
 wire \i43/n320 ;
 wire \i43/n321 ;
 wire \i43/n322 ;
 wire \i43/n323 ;
 wire \i43/n324 ;
 wire \i43/n325 ;
 wire \i43/n326 ;
 wire \i43/n327 ;
 wire \i43/n328 ;
 wire \i43/n329 ;
 wire \i43/n33 ;
 wire \i43/n330 ;
 wire \i43/n331 ;
 wire \i43/n332 ;
 wire \i43/n333 ;
 wire \i43/n334 ;
 wire \i43/n335 ;
 wire \i43/n336 ;
 wire \i43/n337 ;
 wire \i43/n338 ;
 wire \i43/n339 ;
 wire \i43/n34 ;
 wire \i43/n340 ;
 wire \i43/n341 ;
 wire \i43/n342 ;
 wire \i43/n343 ;
 wire \i43/n344 ;
 wire \i43/n345 ;
 wire \i43/n346 ;
 wire \i43/n347 ;
 wire \i43/n348 ;
 wire \i43/n349 ;
 wire \i43/n35 ;
 wire \i43/n350 ;
 wire \i43/n351 ;
 wire \i43/n352 ;
 wire \i43/n353 ;
 wire \i43/n354 ;
 wire \i43/n355 ;
 wire \i43/n356 ;
 wire \i43/n357 ;
 wire \i43/n358 ;
 wire \i43/n359 ;
 wire \i43/n36 ;
 wire \i43/n360 ;
 wire \i43/n361 ;
 wire \i43/n362 ;
 wire \i43/n363 ;
 wire \i43/n364 ;
 wire \i43/n365 ;
 wire \i43/n366 ;
 wire \i43/n367 ;
 wire \i43/n368 ;
 wire \i43/n369 ;
 wire \i43/n37 ;
 wire \i43/n370 ;
 wire \i43/n371 ;
 wire \i43/n372 ;
 wire \i43/n373 ;
 wire \i43/n374 ;
 wire \i43/n375 ;
 wire \i43/n376 ;
 wire \i43/n377 ;
 wire \i43/n378 ;
 wire \i43/n379 ;
 wire \i43/n38 ;
 wire \i43/n380 ;
 wire \i43/n381 ;
 wire \i43/n382 ;
 wire \i43/n383 ;
 wire \i43/n384 ;
 wire \i43/n385 ;
 wire \i43/n386 ;
 wire \i43/n387 ;
 wire \i43/n388 ;
 wire \i43/n389 ;
 wire \i43/n39 ;
 wire \i43/n390 ;
 wire \i43/n391 ;
 wire \i43/n392 ;
 wire \i43/n393 ;
 wire \i43/n394 ;
 wire \i43/n395 ;
 wire \i43/n396 ;
 wire \i43/n397 ;
 wire \i43/n398 ;
 wire \i43/n399 ;
 wire \i43/n4 ;
 wire \i43/n40 ;
 wire \i43/n400 ;
 wire \i43/n401 ;
 wire \i43/n402 ;
 wire \i43/n403 ;
 wire \i43/n404 ;
 wire \i43/n405 ;
 wire \i43/n406 ;
 wire \i43/n407 ;
 wire \i43/n408 ;
 wire \i43/n409 ;
 wire \i43/n41 ;
 wire \i43/n410 ;
 wire \i43/n411 ;
 wire \i43/n412 ;
 wire \i43/n413 ;
 wire \i43/n414 ;
 wire \i43/n415 ;
 wire \i43/n416 ;
 wire \i43/n417 ;
 wire \i43/n418 ;
 wire \i43/n419 ;
 wire \i43/n42 ;
 wire \i43/n420 ;
 wire \i43/n421 ;
 wire \i43/n422 ;
 wire \i43/n423 ;
 wire \i43/n424 ;
 wire \i43/n425 ;
 wire \i43/n426 ;
 wire \i43/n427 ;
 wire \i43/n428 ;
 wire \i43/n429 ;
 wire \i43/n43 ;
 wire \i43/n430 ;
 wire \i43/n431 ;
 wire \i43/n432 ;
 wire \i43/n433 ;
 wire \i43/n434 ;
 wire \i43/n435 ;
 wire \i43/n436 ;
 wire \i43/n437 ;
 wire \i43/n438 ;
 wire \i43/n439 ;
 wire \i43/n44 ;
 wire \i43/n440 ;
 wire \i43/n441 ;
 wire \i43/n442 ;
 wire \i43/n443 ;
 wire \i43/n444 ;
 wire \i43/n445 ;
 wire \i43/n446 ;
 wire \i43/n447 ;
 wire \i43/n448 ;
 wire \i43/n449 ;
 wire \i43/n45 ;
 wire \i43/n450 ;
 wire \i43/n451 ;
 wire \i43/n452 ;
 wire \i43/n453 ;
 wire \i43/n454 ;
 wire \i43/n455 ;
 wire \i43/n456 ;
 wire \i43/n457 ;
 wire \i43/n458 ;
 wire \i43/n459 ;
 wire \i43/n46 ;
 wire \i43/n460 ;
 wire \i43/n461 ;
 wire \i43/n462 ;
 wire \i43/n463 ;
 wire \i43/n464 ;
 wire \i43/n47 ;
 wire \i43/n48 ;
 wire \i43/n49 ;
 wire \i43/n5 ;
 wire \i43/n50 ;
 wire \i43/n51 ;
 wire \i43/n52 ;
 wire \i43/n53 ;
 wire \i43/n54 ;
 wire \i43/n55 ;
 wire \i43/n56 ;
 wire \i43/n57 ;
 wire \i43/n58 ;
 wire \i43/n59 ;
 wire \i43/n6 ;
 wire \i43/n60 ;
 wire \i43/n61 ;
 wire \i43/n62 ;
 wire \i43/n63 ;
 wire \i43/n64 ;
 wire \i43/n65 ;
 wire \i43/n66 ;
 wire \i43/n67 ;
 wire \i43/n68 ;
 wire \i43/n69 ;
 wire \i43/n7 ;
 wire \i43/n70 ;
 wire \i43/n71 ;
 wire \i43/n72 ;
 wire \i43/n73 ;
 wire \i43/n74 ;
 wire \i43/n75 ;
 wire \i43/n76 ;
 wire \i43/n77 ;
 wire \i43/n78 ;
 wire \i43/n79 ;
 wire \i43/n8 ;
 wire \i43/n80 ;
 wire \i43/n81 ;
 wire \i43/n82 ;
 wire \i43/n83 ;
 wire \i43/n84 ;
 wire \i43/n85 ;
 wire \i43/n86 ;
 wire \i43/n87 ;
 wire \i43/n88 ;
 wire \i43/n89 ;
 wire \i43/n9 ;
 wire \i43/n90 ;
 wire \i43/n91 ;
 wire \i43/n92 ;
 wire \i43/n93 ;
 wire \i43/n94 ;
 wire \i43/n95 ;
 wire \i43/n96 ;
 wire \i43/n97 ;
 wire \i43/n98 ;
 wire \i43/n99 ;
 wire \i43/i45/n10 ;
 wire \i43/i45/n11 ;
 wire \i43/i45/n12 ;
 wire \i43/i45/n13 ;
 wire \i43/i45/n14 ;
 wire \i43/i45/n15 ;
 wire \i43/i45/n16 ;
 wire \i43/i45/n17 ;
 wire \i43/i45/n18 ;
 wire \i43/i45/n19 ;
 wire \i43/i45/n2 ;
 wire \i43/i45/n20 ;
 wire \i43/i45/n21 ;
 wire \i43/i45/n22 ;
 wire \i43/i45/n23 ;
 wire \i43/i45/n24 ;
 wire \i43/i45/n25 ;
 wire \i43/i45/n26 ;
 wire \i43/i45/n27 ;
 wire \i43/i45/n3 ;
 wire \i43/i45/n4 ;
 wire \i43/i45/n5 ;
 wire \i43/i45/n6 ;
 wire \i43/i45/n7 ;
 wire \i43/i45/n8 ;
 wire \i43/i45/n9 ;
 wire \i43/i46/n0 ;
 wire \i43/i46/n1 ;
 wire \i43/i46/n10 ;
 wire \i43/i46/n100 ;
 wire \i43/i46/n101 ;
 wire \i43/i46/n102 ;
 wire \i43/i46/n103 ;
 wire \i43/i46/n104 ;
 wire \i43/i46/n105 ;
 wire \i43/i46/n106 ;
 wire \i43/i46/n107 ;
 wire \i43/i46/n108 ;
 wire \i43/i46/n109 ;
 wire \i43/i46/n11 ;
 wire \i43/i46/n110 ;
 wire \i43/i46/n111 ;
 wire \i43/i46/n112 ;
 wire \i43/i46/n113 ;
 wire \i43/i46/n114 ;
 wire \i43/i46/n115 ;
 wire \i43/i46/n116 ;
 wire \i43/i46/n117 ;
 wire \i43/i46/n118 ;
 wire \i43/i46/n119 ;
 wire \i43/i46/n12 ;
 wire \i43/i46/n120 ;
 wire \i43/i46/n121 ;
 wire \i43/i46/n122 ;
 wire \i43/i46/n123 ;
 wire \i43/i46/n124 ;
 wire \i43/i46/n125 ;
 wire \i43/i46/n126 ;
 wire \i43/i46/n127 ;
 wire \i43/i46/n128 ;
 wire \i43/i46/n129 ;
 wire \i43/i46/n13 ;
 wire \i43/i46/n130 ;
 wire \i43/i46/n131 ;
 wire \i43/i46/n132 ;
 wire \i43/i46/n133 ;
 wire \i43/i46/n134 ;
 wire \i43/i46/n135 ;
 wire \i43/i46/n136 ;
 wire \i43/i46/n137 ;
 wire \i43/i46/n138 ;
 wire \i43/i46/n139 ;
 wire \i43/i46/n14 ;
 wire \i43/i46/n140 ;
 wire \i43/i46/n141 ;
 wire \i43/i46/n142 ;
 wire \i43/i46/n143 ;
 wire \i43/i46/n144 ;
 wire \i43/i46/n145 ;
 wire \i43/i46/n146 ;
 wire \i43/i46/n147 ;
 wire \i43/i46/n148 ;
 wire \i43/i46/n149 ;
 wire \i43/i46/n15 ;
 wire \i43/i46/n150 ;
 wire \i43/i46/n151 ;
 wire \i43/i46/n152 ;
 wire \i43/i46/n153 ;
 wire \i43/i46/n154 ;
 wire \i43/i46/n155 ;
 wire \i43/i46/n156 ;
 wire \i43/i46/n157 ;
 wire \i43/i46/n158 ;
 wire \i43/i46/n159 ;
 wire \i43/i46/n16 ;
 wire \i43/i46/n160 ;
 wire \i43/i46/n161 ;
 wire \i43/i46/n162 ;
 wire \i43/i46/n163 ;
 wire \i43/i46/n164 ;
 wire \i43/i46/n165 ;
 wire \i43/i46/n166 ;
 wire \i43/i46/n167 ;
 wire \i43/i46/n168 ;
 wire \i43/i46/n169 ;
 wire \i43/i46/n17 ;
 wire \i43/i46/n170 ;
 wire \i43/i46/n171 ;
 wire \i43/i46/n172 ;
 wire \i43/i46/n173 ;
 wire \i43/i46/n174 ;
 wire \i43/i46/n175 ;
 wire \i43/i46/n176 ;
 wire \i43/i46/n177 ;
 wire \i43/i46/n178 ;
 wire \i43/i46/n179 ;
 wire \i43/i46/n18 ;
 wire \i43/i46/n180 ;
 wire \i43/i46/n181 ;
 wire \i43/i46/n182 ;
 wire \i43/i46/n183 ;
 wire \i43/i46/n184 ;
 wire \i43/i46/n185 ;
 wire \i43/i46/n186 ;
 wire \i43/i46/n187 ;
 wire \i43/i46/n188 ;
 wire \i43/i46/n189 ;
 wire \i43/i46/n19 ;
 wire \i43/i46/n190 ;
 wire \i43/i46/n191 ;
 wire \i43/i46/n192 ;
 wire \i43/i46/n193 ;
 wire \i43/i46/n194 ;
 wire \i43/i46/n195 ;
 wire \i43/i46/n196 ;
 wire \i43/i46/n197 ;
 wire \i43/i46/n198 ;
 wire \i43/i46/n199 ;
 wire \i43/i46/n2 ;
 wire \i43/i46/n20 ;
 wire \i43/i46/n200 ;
 wire \i43/i46/n201 ;
 wire \i43/i46/n202 ;
 wire \i43/i46/n203 ;
 wire \i43/i46/n204 ;
 wire \i43/i46/n205 ;
 wire \i43/i46/n206 ;
 wire \i43/i46/n207 ;
 wire \i43/i46/n208 ;
 wire \i43/i46/n209 ;
 wire \i43/i46/n21 ;
 wire \i43/i46/n210 ;
 wire \i43/i46/n211 ;
 wire \i43/i46/n212 ;
 wire \i43/i46/n213 ;
 wire \i43/i46/n214 ;
 wire \i43/i46/n215 ;
 wire \i43/i46/n216 ;
 wire \i43/i46/n217 ;
 wire \i43/i46/n218 ;
 wire \i43/i46/n219 ;
 wire \i43/i46/n22 ;
 wire \i43/i46/n220 ;
 wire \i43/i46/n221 ;
 wire \i43/i46/n222 ;
 wire \i43/i46/n223 ;
 wire \i43/i46/n224 ;
 wire \i43/i46/n225 ;
 wire \i43/i46/n226 ;
 wire \i43/i46/n227 ;
 wire \i43/i46/n228 ;
 wire \i43/i46/n229 ;
 wire \i43/i46/n23 ;
 wire \i43/i46/n230 ;
 wire \i43/i46/n231 ;
 wire \i43/i46/n232 ;
 wire \i43/i46/n233 ;
 wire \i43/i46/n234 ;
 wire \i43/i46/n235 ;
 wire \i43/i46/n236 ;
 wire \i43/i46/n237 ;
 wire \i43/i46/n238 ;
 wire \i43/i46/n239 ;
 wire \i43/i46/n24 ;
 wire \i43/i46/n240 ;
 wire \i43/i46/n241 ;
 wire \i43/i46/n242 ;
 wire \i43/i46/n243 ;
 wire \i43/i46/n244 ;
 wire \i43/i46/n245 ;
 wire \i43/i46/n246 ;
 wire \i43/i46/n247 ;
 wire \i43/i46/n248 ;
 wire \i43/i46/n249 ;
 wire \i43/i46/n25 ;
 wire \i43/i46/n250 ;
 wire \i43/i46/n251 ;
 wire \i43/i46/n252 ;
 wire \i43/i46/n253 ;
 wire \i43/i46/n254 ;
 wire \i43/i46/n255 ;
 wire \i43/i46/n256 ;
 wire \i43/i46/n257 ;
 wire \i43/i46/n258 ;
 wire \i43/i46/n259 ;
 wire \i43/i46/n26 ;
 wire \i43/i46/n260 ;
 wire \i43/i46/n261 ;
 wire \i43/i46/n262 ;
 wire \i43/i46/n263 ;
 wire \i43/i46/n264 ;
 wire \i43/i46/n265 ;
 wire \i43/i46/n266 ;
 wire \i43/i46/n267 ;
 wire \i43/i46/n268 ;
 wire \i43/i46/n269 ;
 wire \i43/i46/n27 ;
 wire \i43/i46/n270 ;
 wire \i43/i46/n271 ;
 wire \i43/i46/n272 ;
 wire \i43/i46/n273 ;
 wire \i43/i46/n274 ;
 wire \i43/i46/n275 ;
 wire \i43/i46/n276 ;
 wire \i43/i46/n277 ;
 wire \i43/i46/n278 ;
 wire \i43/i46/n279 ;
 wire \i43/i46/n28 ;
 wire \i43/i46/n280 ;
 wire \i43/i46/n281 ;
 wire \i43/i46/n282 ;
 wire \i43/i46/n283 ;
 wire \i43/i46/n284 ;
 wire \i43/i46/n285 ;
 wire \i43/i46/n286 ;
 wire \i43/i46/n287 ;
 wire \i43/i46/n288 ;
 wire \i43/i46/n289 ;
 wire \i43/i46/n29 ;
 wire \i43/i46/n290 ;
 wire \i43/i46/n291 ;
 wire \i43/i46/n292 ;
 wire \i43/i46/n293 ;
 wire \i43/i46/n294 ;
 wire \i43/i46/n295 ;
 wire \i43/i46/n296 ;
 wire \i43/i46/n297 ;
 wire \i43/i46/n298 ;
 wire \i43/i46/n299 ;
 wire \i43/i46/n3 ;
 wire \i43/i46/n30 ;
 wire \i43/i46/n300 ;
 wire \i43/i46/n301 ;
 wire \i43/i46/n302 ;
 wire \i43/i46/n303 ;
 wire \i43/i46/n304 ;
 wire \i43/i46/n305 ;
 wire \i43/i46/n306 ;
 wire \i43/i46/n307 ;
 wire \i43/i46/n308 ;
 wire \i43/i46/n309 ;
 wire \i43/i46/n31 ;
 wire \i43/i46/n310 ;
 wire \i43/i46/n311 ;
 wire \i43/i46/n312 ;
 wire \i43/i46/n313 ;
 wire \i43/i46/n314 ;
 wire \i43/i46/n315 ;
 wire \i43/i46/n316 ;
 wire \i43/i46/n317 ;
 wire \i43/i46/n318 ;
 wire \i43/i46/n319 ;
 wire \i43/i46/n32 ;
 wire \i43/i46/n320 ;
 wire \i43/i46/n321 ;
 wire \i43/i46/n322 ;
 wire \i43/i46/n323 ;
 wire \i43/i46/n324 ;
 wire \i43/i46/n325 ;
 wire \i43/i46/n326 ;
 wire \i43/i46/n327 ;
 wire \i43/i46/n328 ;
 wire \i43/i46/n329 ;
 wire \i43/i46/n33 ;
 wire \i43/i46/n330 ;
 wire \i43/i46/n331 ;
 wire \i43/i46/n332 ;
 wire \i43/i46/n333 ;
 wire \i43/i46/n334 ;
 wire \i43/i46/n335 ;
 wire \i43/i46/n336 ;
 wire \i43/i46/n337 ;
 wire \i43/i46/n338 ;
 wire \i43/i46/n339 ;
 wire \i43/i46/n34 ;
 wire \i43/i46/n340 ;
 wire \i43/i46/n341 ;
 wire \i43/i46/n342 ;
 wire \i43/i46/n343 ;
 wire \i43/i46/n344 ;
 wire \i43/i46/n345 ;
 wire \i43/i46/n346 ;
 wire \i43/i46/n347 ;
 wire \i43/i46/n348 ;
 wire \i43/i46/n349 ;
 wire \i43/i46/n35 ;
 wire \i43/i46/n350 ;
 wire \i43/i46/n351 ;
 wire \i43/i46/n352 ;
 wire \i43/i46/n353 ;
 wire \i43/i46/n354 ;
 wire \i43/i46/n355 ;
 wire \i43/i46/n356 ;
 wire \i43/i46/n357 ;
 wire \i43/i46/n358 ;
 wire \i43/i46/n359 ;
 wire \i43/i46/n36 ;
 wire \i43/i46/n360 ;
 wire \i43/i46/n361 ;
 wire \i43/i46/n362 ;
 wire \i43/i46/n363 ;
 wire \i43/i46/n364 ;
 wire \i43/i46/n365 ;
 wire \i43/i46/n366 ;
 wire \i43/i46/n367 ;
 wire \i43/i46/n368 ;
 wire \i43/i46/n369 ;
 wire \i43/i46/n37 ;
 wire \i43/i46/n370 ;
 wire \i43/i46/n371 ;
 wire \i43/i46/n372 ;
 wire \i43/i46/n373 ;
 wire \i43/i46/n374 ;
 wire \i43/i46/n375 ;
 wire \i43/i46/n376 ;
 wire \i43/i46/n377 ;
 wire \i43/i46/n378 ;
 wire \i43/i46/n379 ;
 wire \i43/i46/n38 ;
 wire \i43/i46/n380 ;
 wire \i43/i46/n381 ;
 wire \i43/i46/n382 ;
 wire \i43/i46/n383 ;
 wire \i43/i46/n384 ;
 wire \i43/i46/n385 ;
 wire \i43/i46/n386 ;
 wire \i43/i46/n387 ;
 wire \i43/i46/n388 ;
 wire \i43/i46/n389 ;
 wire \i43/i46/n39 ;
 wire \i43/i46/n390 ;
 wire \i43/i46/n391 ;
 wire \i43/i46/n392 ;
 wire \i43/i46/n393 ;
 wire \i43/i46/n394 ;
 wire \i43/i46/n395 ;
 wire \i43/i46/n396 ;
 wire \i43/i46/n397 ;
 wire \i43/i46/n398 ;
 wire \i43/i46/n399 ;
 wire \i43/i46/n4 ;
 wire \i43/i46/n40 ;
 wire \i43/i46/n400 ;
 wire \i43/i46/n401 ;
 wire \i43/i46/n402 ;
 wire \i43/i46/n403 ;
 wire \i43/i46/n404 ;
 wire \i43/i46/n405 ;
 wire \i43/i46/n406 ;
 wire \i43/i46/n407 ;
 wire \i43/i46/n408 ;
 wire \i43/i46/n409 ;
 wire \i43/i46/n41 ;
 wire \i43/i46/n410 ;
 wire \i43/i46/n411 ;
 wire \i43/i46/n412 ;
 wire \i43/i46/n413 ;
 wire \i43/i46/n414 ;
 wire \i43/i46/n415 ;
 wire \i43/i46/n416 ;
 wire \i43/i46/n417 ;
 wire \i43/i46/n418 ;
 wire \i43/i46/n419 ;
 wire \i43/i46/n42 ;
 wire \i43/i46/n420 ;
 wire \i43/i46/n421 ;
 wire \i43/i46/n422 ;
 wire \i43/i46/n423 ;
 wire \i43/i46/n424 ;
 wire \i43/i46/n425 ;
 wire \i43/i46/n426 ;
 wire \i43/i46/n427 ;
 wire \i43/i46/n428 ;
 wire \i43/i46/n429 ;
 wire \i43/i46/n43 ;
 wire \i43/i46/n430 ;
 wire \i43/i46/n431 ;
 wire \i43/i46/n432 ;
 wire \i43/i46/n433 ;
 wire \i43/i46/n434 ;
 wire \i43/i46/n435 ;
 wire \i43/i46/n436 ;
 wire \i43/i46/n437 ;
 wire \i43/i46/n438 ;
 wire \i43/i46/n439 ;
 wire \i43/i46/n44 ;
 wire \i43/i46/n440 ;
 wire \i43/i46/n441 ;
 wire \i43/i46/n442 ;
 wire \i43/i46/n443 ;
 wire \i43/i46/n444 ;
 wire \i43/i46/n445 ;
 wire \i43/i46/n446 ;
 wire \i43/i46/n447 ;
 wire \i43/i46/n448 ;
 wire \i43/i46/n449 ;
 wire \i43/i46/n45 ;
 wire \i43/i46/n450 ;
 wire \i43/i46/n451 ;
 wire \i43/i46/n452 ;
 wire \i43/i46/n453 ;
 wire \i43/i46/n454 ;
 wire \i43/i46/n455 ;
 wire \i43/i46/n456 ;
 wire \i43/i46/n457 ;
 wire \i43/i46/n458 ;
 wire \i43/i46/n459 ;
 wire \i43/i46/n46 ;
 wire \i43/i46/n460 ;
 wire \i43/i46/n461 ;
 wire \i43/i46/n462 ;
 wire \i43/i46/n463 ;
 wire \i43/i46/n464 ;
 wire \i43/i46/n465 ;
 wire \i43/i46/n466 ;
 wire \i43/i46/n467 ;
 wire \i43/i46/n468 ;
 wire \i43/i46/n469 ;
 wire \i43/i46/n47 ;
 wire \i43/i46/n470 ;
 wire \i43/i46/n471 ;
 wire \i43/i46/n472 ;
 wire \i43/i46/n473 ;
 wire \i43/i46/n474 ;
 wire \i43/i46/n475 ;
 wire \i43/i46/n476 ;
 wire \i43/i46/n477 ;
 wire \i43/i46/n478 ;
 wire \i43/i46/n479 ;
 wire \i43/i46/n48 ;
 wire \i43/i46/n480 ;
 wire \i43/i46/n481 ;
 wire \i43/i46/n482 ;
 wire \i43/i46/n483 ;
 wire \i43/i46/n484 ;
 wire \i43/i46/n485 ;
 wire \i43/i46/n486 ;
 wire \i43/i46/n487 ;
 wire \i43/i46/n488 ;
 wire \i43/i46/n489 ;
 wire \i43/i46/n49 ;
 wire \i43/i46/n490 ;
 wire \i43/i46/n491 ;
 wire \i43/i46/n492 ;
 wire \i43/i46/n493 ;
 wire \i43/i46/n494 ;
 wire \i43/i46/n495 ;
 wire \i43/i46/n496 ;
 wire \i43/i46/n497 ;
 wire \i43/i46/n498 ;
 wire \i43/i46/n499 ;
 wire \i43/i46/n5 ;
 wire \i43/i46/n50 ;
 wire \i43/i46/n500 ;
 wire \i43/i46/n501 ;
 wire \i43/i46/n502 ;
 wire \i43/i46/n503 ;
 wire \i43/i46/n504 ;
 wire \i43/i46/n505 ;
 wire \i43/i46/n506 ;
 wire \i43/i46/n507 ;
 wire \i43/i46/n508 ;
 wire \i43/i46/n509 ;
 wire \i43/i46/n51 ;
 wire \i43/i46/n510 ;
 wire \i43/i46/n511 ;
 wire \i43/i46/n512 ;
 wire \i43/i46/n513 ;
 wire \i43/i46/n514 ;
 wire \i43/i46/n515 ;
 wire \i43/i46/n516 ;
 wire \i43/i46/n517 ;
 wire \i43/i46/n518 ;
 wire \i43/i46/n519 ;
 wire \i43/i46/n52 ;
 wire \i43/i46/n53 ;
 wire \i43/i46/n54 ;
 wire \i43/i46/n55 ;
 wire \i43/i46/n56 ;
 wire \i43/i46/n57 ;
 wire \i43/i46/n58 ;
 wire \i43/i46/n59 ;
 wire \i43/i46/n6 ;
 wire \i43/i46/n60 ;
 wire \i43/i46/n61 ;
 wire \i43/i46/n62 ;
 wire \i43/i46/n63 ;
 wire \i43/i46/n64 ;
 wire \i43/i46/n65 ;
 wire \i43/i46/n66 ;
 wire \i43/i46/n67 ;
 wire \i43/i46/n68 ;
 wire \i43/i46/n69 ;
 wire \i43/i46/n7 ;
 wire \i43/i46/n70 ;
 wire \i43/i46/n71 ;
 wire \i43/i46/n72 ;
 wire \i43/i46/n73 ;
 wire \i43/i46/n74 ;
 wire \i43/i46/n75 ;
 wire \i43/i46/n76 ;
 wire \i43/i46/n77 ;
 wire \i43/i46/n78 ;
 wire \i43/i46/n79 ;
 wire \i43/i46/n8 ;
 wire \i43/i46/n80 ;
 wire \i43/i46/n81 ;
 wire \i43/i46/n82 ;
 wire \i43/i46/n83 ;
 wire \i43/i46/n84 ;
 wire \i43/i46/n85 ;
 wire \i43/i46/n86 ;
 wire \i43/i46/n87 ;
 wire \i43/i46/n88 ;
 wire \i43/i46/n89 ;
 wire \i43/i46/n9 ;
 wire \i43/i46/n90 ;
 wire \i43/i46/n91 ;
 wire \i43/i46/n92 ;
 wire \i43/i46/n93 ;
 wire \i43/i46/n94 ;
 wire \i43/i46/n95 ;
 wire \i43/i46/n96 ;
 wire \i43/i46/n97 ;
 wire \i43/i46/n98 ;
 wire \i43/i46/n99 ;
 wire \i43/i47/n0 ;
 wire \i43/i47/n1 ;
 wire \i43/i47/n10 ;
 wire \i43/i47/n100 ;
 wire \i43/i47/n101 ;
 wire \i43/i47/n102 ;
 wire \i43/i47/n103 ;
 wire \i43/i47/n104 ;
 wire \i43/i47/n105 ;
 wire \i43/i47/n106 ;
 wire \i43/i47/n107 ;
 wire \i43/i47/n108 ;
 wire \i43/i47/n109 ;
 wire \i43/i47/n11 ;
 wire \i43/i47/n110 ;
 wire \i43/i47/n111 ;
 wire \i43/i47/n112 ;
 wire \i43/i47/n113 ;
 wire \i43/i47/n114 ;
 wire \i43/i47/n115 ;
 wire \i43/i47/n116 ;
 wire \i43/i47/n117 ;
 wire \i43/i47/n118 ;
 wire \i43/i47/n119 ;
 wire \i43/i47/n12 ;
 wire \i43/i47/n120 ;
 wire \i43/i47/n121 ;
 wire \i43/i47/n122 ;
 wire \i43/i47/n123 ;
 wire \i43/i47/n124 ;
 wire \i43/i47/n125 ;
 wire \i43/i47/n126 ;
 wire \i43/i47/n127 ;
 wire \i43/i47/n128 ;
 wire \i43/i47/n129 ;
 wire \i43/i47/n13 ;
 wire \i43/i47/n130 ;
 wire \i43/i47/n131 ;
 wire \i43/i47/n132 ;
 wire \i43/i47/n133 ;
 wire \i43/i47/n134 ;
 wire \i43/i47/n135 ;
 wire \i43/i47/n136 ;
 wire \i43/i47/n137 ;
 wire \i43/i47/n138 ;
 wire \i43/i47/n139 ;
 wire \i43/i47/n14 ;
 wire \i43/i47/n140 ;
 wire \i43/i47/n141 ;
 wire \i43/i47/n142 ;
 wire \i43/i47/n143 ;
 wire \i43/i47/n144 ;
 wire \i43/i47/n145 ;
 wire \i43/i47/n146 ;
 wire \i43/i47/n147 ;
 wire \i43/i47/n148 ;
 wire \i43/i47/n149 ;
 wire \i43/i47/n15 ;
 wire \i43/i47/n150 ;
 wire \i43/i47/n151 ;
 wire \i43/i47/n152 ;
 wire \i43/i47/n153 ;
 wire \i43/i47/n154 ;
 wire \i43/i47/n155 ;
 wire \i43/i47/n156 ;
 wire \i43/i47/n157 ;
 wire \i43/i47/n158 ;
 wire \i43/i47/n159 ;
 wire \i43/i47/n16 ;
 wire \i43/i47/n160 ;
 wire \i43/i47/n161 ;
 wire \i43/i47/n162 ;
 wire \i43/i47/n163 ;
 wire \i43/i47/n164 ;
 wire \i43/i47/n165 ;
 wire \i43/i47/n166 ;
 wire \i43/i47/n167 ;
 wire \i43/i47/n168 ;
 wire \i43/i47/n169 ;
 wire \i43/i47/n17 ;
 wire \i43/i47/n170 ;
 wire \i43/i47/n171 ;
 wire \i43/i47/n172 ;
 wire \i43/i47/n173 ;
 wire \i43/i47/n174 ;
 wire \i43/i47/n175 ;
 wire \i43/i47/n176 ;
 wire \i43/i47/n177 ;
 wire \i43/i47/n178 ;
 wire \i43/i47/n179 ;
 wire \i43/i47/n18 ;
 wire \i43/i47/n180 ;
 wire \i43/i47/n181 ;
 wire \i43/i47/n182 ;
 wire \i43/i47/n183 ;
 wire \i43/i47/n184 ;
 wire \i43/i47/n185 ;
 wire \i43/i47/n186 ;
 wire \i43/i47/n187 ;
 wire \i43/i47/n188 ;
 wire \i43/i47/n189 ;
 wire \i43/i47/n19 ;
 wire \i43/i47/n190 ;
 wire \i43/i47/n191 ;
 wire \i43/i47/n192 ;
 wire \i43/i47/n193 ;
 wire \i43/i47/n194 ;
 wire \i43/i47/n195 ;
 wire \i43/i47/n196 ;
 wire \i43/i47/n197 ;
 wire \i43/i47/n198 ;
 wire \i43/i47/n199 ;
 wire \i43/i47/n2 ;
 wire \i43/i47/n20 ;
 wire \i43/i47/n200 ;
 wire \i43/i47/n201 ;
 wire \i43/i47/n202 ;
 wire \i43/i47/n203 ;
 wire \i43/i47/n204 ;
 wire \i43/i47/n205 ;
 wire \i43/i47/n206 ;
 wire \i43/i47/n207 ;
 wire \i43/i47/n208 ;
 wire \i43/i47/n209 ;
 wire \i43/i47/n21 ;
 wire \i43/i47/n210 ;
 wire \i43/i47/n211 ;
 wire \i43/i47/n212 ;
 wire \i43/i47/n213 ;
 wire \i43/i47/n214 ;
 wire \i43/i47/n215 ;
 wire \i43/i47/n216 ;
 wire \i43/i47/n217 ;
 wire \i43/i47/n218 ;
 wire \i43/i47/n219 ;
 wire \i43/i47/n22 ;
 wire \i43/i47/n220 ;
 wire \i43/i47/n221 ;
 wire \i43/i47/n222 ;
 wire \i43/i47/n223 ;
 wire \i43/i47/n224 ;
 wire \i43/i47/n225 ;
 wire \i43/i47/n226 ;
 wire \i43/i47/n227 ;
 wire \i43/i47/n228 ;
 wire \i43/i47/n229 ;
 wire \i43/i47/n23 ;
 wire \i43/i47/n230 ;
 wire \i43/i47/n231 ;
 wire \i43/i47/n232 ;
 wire \i43/i47/n233 ;
 wire \i43/i47/n234 ;
 wire \i43/i47/n235 ;
 wire \i43/i47/n236 ;
 wire \i43/i47/n237 ;
 wire \i43/i47/n238 ;
 wire \i43/i47/n239 ;
 wire \i43/i47/n24 ;
 wire \i43/i47/n240 ;
 wire \i43/i47/n241 ;
 wire \i43/i47/n242 ;
 wire \i43/i47/n243 ;
 wire \i43/i47/n244 ;
 wire \i43/i47/n245 ;
 wire \i43/i47/n246 ;
 wire \i43/i47/n247 ;
 wire \i43/i47/n248 ;
 wire \i43/i47/n249 ;
 wire \i43/i47/n25 ;
 wire \i43/i47/n250 ;
 wire \i43/i47/n251 ;
 wire \i43/i47/n252 ;
 wire \i43/i47/n253 ;
 wire \i43/i47/n254 ;
 wire \i43/i47/n255 ;
 wire \i43/i47/n256 ;
 wire \i43/i47/n257 ;
 wire \i43/i47/n258 ;
 wire \i43/i47/n259 ;
 wire \i43/i47/n26 ;
 wire \i43/i47/n260 ;
 wire \i43/i47/n261 ;
 wire \i43/i47/n262 ;
 wire \i43/i47/n263 ;
 wire \i43/i47/n264 ;
 wire \i43/i47/n265 ;
 wire \i43/i47/n266 ;
 wire \i43/i47/n267 ;
 wire \i43/i47/n268 ;
 wire \i43/i47/n269 ;
 wire \i43/i47/n27 ;
 wire \i43/i47/n270 ;
 wire \i43/i47/n271 ;
 wire \i43/i47/n272 ;
 wire \i43/i47/n273 ;
 wire \i43/i47/n274 ;
 wire \i43/i47/n275 ;
 wire \i43/i47/n276 ;
 wire \i43/i47/n277 ;
 wire \i43/i47/n278 ;
 wire \i43/i47/n279 ;
 wire \i43/i47/n28 ;
 wire \i43/i47/n280 ;
 wire \i43/i47/n281 ;
 wire \i43/i47/n282 ;
 wire \i43/i47/n283 ;
 wire \i43/i47/n284 ;
 wire \i43/i47/n285 ;
 wire \i43/i47/n286 ;
 wire \i43/i47/n287 ;
 wire \i43/i47/n288 ;
 wire \i43/i47/n289 ;
 wire \i43/i47/n29 ;
 wire \i43/i47/n290 ;
 wire \i43/i47/n291 ;
 wire \i43/i47/n292 ;
 wire \i43/i47/n293 ;
 wire \i43/i47/n294 ;
 wire \i43/i47/n295 ;
 wire \i43/i47/n296 ;
 wire \i43/i47/n297 ;
 wire \i43/i47/n298 ;
 wire \i43/i47/n299 ;
 wire \i43/i47/n3 ;
 wire \i43/i47/n30 ;
 wire \i43/i47/n300 ;
 wire \i43/i47/n301 ;
 wire \i43/i47/n302 ;
 wire \i43/i47/n303 ;
 wire \i43/i47/n304 ;
 wire \i43/i47/n305 ;
 wire \i43/i47/n306 ;
 wire \i43/i47/n307 ;
 wire \i43/i47/n308 ;
 wire \i43/i47/n309 ;
 wire \i43/i47/n31 ;
 wire \i43/i47/n310 ;
 wire \i43/i47/n311 ;
 wire \i43/i47/n312 ;
 wire \i43/i47/n313 ;
 wire \i43/i47/n314 ;
 wire \i43/i47/n315 ;
 wire \i43/i47/n316 ;
 wire \i43/i47/n317 ;
 wire \i43/i47/n318 ;
 wire \i43/i47/n319 ;
 wire \i43/i47/n32 ;
 wire \i43/i47/n320 ;
 wire \i43/i47/n321 ;
 wire \i43/i47/n322 ;
 wire \i43/i47/n323 ;
 wire \i43/i47/n324 ;
 wire \i43/i47/n325 ;
 wire \i43/i47/n326 ;
 wire \i43/i47/n327 ;
 wire \i43/i47/n328 ;
 wire \i43/i47/n329 ;
 wire \i43/i47/n33 ;
 wire \i43/i47/n330 ;
 wire \i43/i47/n331 ;
 wire \i43/i47/n332 ;
 wire \i43/i47/n333 ;
 wire \i43/i47/n334 ;
 wire \i43/i47/n335 ;
 wire \i43/i47/n336 ;
 wire \i43/i47/n337 ;
 wire \i43/i47/n338 ;
 wire \i43/i47/n339 ;
 wire \i43/i47/n34 ;
 wire \i43/i47/n340 ;
 wire \i43/i47/n341 ;
 wire \i43/i47/n342 ;
 wire \i43/i47/n343 ;
 wire \i43/i47/n344 ;
 wire \i43/i47/n345 ;
 wire \i43/i47/n346 ;
 wire \i43/i47/n347 ;
 wire \i43/i47/n348 ;
 wire \i43/i47/n349 ;
 wire \i43/i47/n35 ;
 wire \i43/i47/n350 ;
 wire \i43/i47/n351 ;
 wire \i43/i47/n352 ;
 wire \i43/i47/n353 ;
 wire \i43/i47/n354 ;
 wire \i43/i47/n355 ;
 wire \i43/i47/n356 ;
 wire \i43/i47/n357 ;
 wire \i43/i47/n358 ;
 wire \i43/i47/n359 ;
 wire \i43/i47/n36 ;
 wire \i43/i47/n360 ;
 wire \i43/i47/n361 ;
 wire \i43/i47/n362 ;
 wire \i43/i47/n363 ;
 wire \i43/i47/n364 ;
 wire \i43/i47/n365 ;
 wire \i43/i47/n366 ;
 wire \i43/i47/n367 ;
 wire \i43/i47/n368 ;
 wire \i43/i47/n369 ;
 wire \i43/i47/n37 ;
 wire \i43/i47/n370 ;
 wire \i43/i47/n371 ;
 wire \i43/i47/n372 ;
 wire \i43/i47/n373 ;
 wire \i43/i47/n374 ;
 wire \i43/i47/n375 ;
 wire \i43/i47/n376 ;
 wire \i43/i47/n377 ;
 wire \i43/i47/n378 ;
 wire \i43/i47/n379 ;
 wire \i43/i47/n38 ;
 wire \i43/i47/n380 ;
 wire \i43/i47/n381 ;
 wire \i43/i47/n382 ;
 wire \i43/i47/n383 ;
 wire \i43/i47/n384 ;
 wire \i43/i47/n385 ;
 wire \i43/i47/n386 ;
 wire \i43/i47/n387 ;
 wire \i43/i47/n388 ;
 wire \i43/i47/n389 ;
 wire \i43/i47/n39 ;
 wire \i43/i47/n390 ;
 wire \i43/i47/n391 ;
 wire \i43/i47/n392 ;
 wire \i43/i47/n393 ;
 wire \i43/i47/n394 ;
 wire \i43/i47/n395 ;
 wire \i43/i47/n396 ;
 wire \i43/i47/n397 ;
 wire \i43/i47/n398 ;
 wire \i43/i47/n399 ;
 wire \i43/i47/n4 ;
 wire \i43/i47/n40 ;
 wire \i43/i47/n400 ;
 wire \i43/i47/n401 ;
 wire \i43/i47/n402 ;
 wire \i43/i47/n403 ;
 wire \i43/i47/n404 ;
 wire \i43/i47/n405 ;
 wire \i43/i47/n406 ;
 wire \i43/i47/n407 ;
 wire \i43/i47/n408 ;
 wire \i43/i47/n409 ;
 wire \i43/i47/n41 ;
 wire \i43/i47/n410 ;
 wire \i43/i47/n411 ;
 wire \i43/i47/n412 ;
 wire \i43/i47/n413 ;
 wire \i43/i47/n414 ;
 wire \i43/i47/n415 ;
 wire \i43/i47/n416 ;
 wire \i43/i47/n417 ;
 wire \i43/i47/n418 ;
 wire \i43/i47/n419 ;
 wire \i43/i47/n42 ;
 wire \i43/i47/n420 ;
 wire \i43/i47/n421 ;
 wire \i43/i47/n422 ;
 wire \i43/i47/n423 ;
 wire \i43/i47/n424 ;
 wire \i43/i47/n425 ;
 wire \i43/i47/n426 ;
 wire \i43/i47/n427 ;
 wire \i43/i47/n428 ;
 wire \i43/i47/n429 ;
 wire \i43/i47/n43 ;
 wire \i43/i47/n430 ;
 wire \i43/i47/n431 ;
 wire \i43/i47/n432 ;
 wire \i43/i47/n433 ;
 wire \i43/i47/n434 ;
 wire \i43/i47/n435 ;
 wire \i43/i47/n436 ;
 wire \i43/i47/n437 ;
 wire \i43/i47/n438 ;
 wire \i43/i47/n439 ;
 wire \i43/i47/n44 ;
 wire \i43/i47/n440 ;
 wire \i43/i47/n441 ;
 wire \i43/i47/n442 ;
 wire \i43/i47/n443 ;
 wire \i43/i47/n444 ;
 wire \i43/i47/n445 ;
 wire \i43/i47/n446 ;
 wire \i43/i47/n447 ;
 wire \i43/i47/n448 ;
 wire \i43/i47/n449 ;
 wire \i43/i47/n45 ;
 wire \i43/i47/n450 ;
 wire \i43/i47/n451 ;
 wire \i43/i47/n452 ;
 wire \i43/i47/n453 ;
 wire \i43/i47/n454 ;
 wire \i43/i47/n455 ;
 wire \i43/i47/n456 ;
 wire \i43/i47/n457 ;
 wire \i43/i47/n458 ;
 wire \i43/i47/n459 ;
 wire \i43/i47/n46 ;
 wire \i43/i47/n460 ;
 wire \i43/i47/n461 ;
 wire \i43/i47/n462 ;
 wire \i43/i47/n463 ;
 wire \i43/i47/n464 ;
 wire \i43/i47/n465 ;
 wire \i43/i47/n466 ;
 wire \i43/i47/n467 ;
 wire \i43/i47/n468 ;
 wire \i43/i47/n469 ;
 wire \i43/i47/n47 ;
 wire \i43/i47/n470 ;
 wire \i43/i47/n471 ;
 wire \i43/i47/n472 ;
 wire \i43/i47/n473 ;
 wire \i43/i47/n474 ;
 wire \i43/i47/n475 ;
 wire \i43/i47/n476 ;
 wire \i43/i47/n477 ;
 wire \i43/i47/n478 ;
 wire \i43/i47/n479 ;
 wire \i43/i47/n48 ;
 wire \i43/i47/n480 ;
 wire \i43/i47/n481 ;
 wire \i43/i47/n482 ;
 wire \i43/i47/n483 ;
 wire \i43/i47/n484 ;
 wire \i43/i47/n485 ;
 wire \i43/i47/n486 ;
 wire \i43/i47/n487 ;
 wire \i43/i47/n488 ;
 wire \i43/i47/n489 ;
 wire \i43/i47/n49 ;
 wire \i43/i47/n490 ;
 wire \i43/i47/n491 ;
 wire \i43/i47/n492 ;
 wire \i43/i47/n493 ;
 wire \i43/i47/n494 ;
 wire \i43/i47/n495 ;
 wire \i43/i47/n496 ;
 wire \i43/i47/n497 ;
 wire \i43/i47/n498 ;
 wire \i43/i47/n499 ;
 wire \i43/i47/n5 ;
 wire \i43/i47/n50 ;
 wire \i43/i47/n500 ;
 wire \i43/i47/n501 ;
 wire \i43/i47/n502 ;
 wire \i43/i47/n503 ;
 wire \i43/i47/n504 ;
 wire \i43/i47/n505 ;
 wire \i43/i47/n506 ;
 wire \i43/i47/n507 ;
 wire \i43/i47/n508 ;
 wire \i43/i47/n509 ;
 wire \i43/i47/n51 ;
 wire \i43/i47/n510 ;
 wire \i43/i47/n511 ;
 wire \i43/i47/n512 ;
 wire \i43/i47/n513 ;
 wire \i43/i47/n514 ;
 wire \i43/i47/n52 ;
 wire \i43/i47/n53 ;
 wire \i43/i47/n54 ;
 wire \i43/i47/n55 ;
 wire \i43/i47/n56 ;
 wire \i43/i47/n57 ;
 wire \i43/i47/n58 ;
 wire \i43/i47/n59 ;
 wire \i43/i47/n6 ;
 wire \i43/i47/n60 ;
 wire \i43/i47/n61 ;
 wire \i43/i47/n62 ;
 wire \i43/i47/n63 ;
 wire \i43/i47/n64 ;
 wire \i43/i47/n65 ;
 wire \i43/i47/n66 ;
 wire \i43/i47/n67 ;
 wire \i43/i47/n68 ;
 wire \i43/i47/n69 ;
 wire \i43/i47/n7 ;
 wire \i43/i47/n70 ;
 wire \i43/i47/n71 ;
 wire \i43/i47/n72 ;
 wire \i43/i47/n73 ;
 wire \i43/i47/n74 ;
 wire \i43/i47/n75 ;
 wire \i43/i47/n76 ;
 wire \i43/i47/n77 ;
 wire \i43/i47/n78 ;
 wire \i43/i47/n79 ;
 wire \i43/i47/n8 ;
 wire \i43/i47/n80 ;
 wire \i43/i47/n81 ;
 wire \i43/i47/n82 ;
 wire \i43/i47/n83 ;
 wire \i43/i47/n84 ;
 wire \i43/i47/n85 ;
 wire \i43/i47/n86 ;
 wire \i43/i47/n87 ;
 wire \i43/i47/n88 ;
 wire \i43/i47/n89 ;
 wire \i43/i47/n9 ;
 wire \i43/i47/n90 ;
 wire \i43/i47/n91 ;
 wire \i43/i47/n92 ;
 wire \i43/i47/n93 ;
 wire \i43/i47/n94 ;
 wire \i43/i47/n95 ;
 wire \i43/i47/n96 ;
 wire \i43/i47/n97 ;
 wire \i43/i47/n98 ;
 wire \i43/i47/n99 ;
 wire \i43/i48/n0 ;
 wire \i43/i48/n1 ;
 wire \i43/i48/n10 ;
 wire \i43/i48/n100 ;
 wire \i43/i48/n101 ;
 wire \i43/i48/n102 ;
 wire \i43/i48/n103 ;
 wire \i43/i48/n104 ;
 wire \i43/i48/n105 ;
 wire \i43/i48/n106 ;
 wire \i43/i48/n107 ;
 wire \i43/i48/n108 ;
 wire \i43/i48/n109 ;
 wire \i43/i48/n11 ;
 wire \i43/i48/n110 ;
 wire \i43/i48/n111 ;
 wire \i43/i48/n112 ;
 wire \i43/i48/n113 ;
 wire \i43/i48/n114 ;
 wire \i43/i48/n115 ;
 wire \i43/i48/n116 ;
 wire \i43/i48/n117 ;
 wire \i43/i48/n118 ;
 wire \i43/i48/n119 ;
 wire \i43/i48/n12 ;
 wire \i43/i48/n120 ;
 wire \i43/i48/n121 ;
 wire \i43/i48/n122 ;
 wire \i43/i48/n123 ;
 wire \i43/i48/n124 ;
 wire \i43/i48/n125 ;
 wire \i43/i48/n126 ;
 wire \i43/i48/n127 ;
 wire \i43/i48/n128 ;
 wire \i43/i48/n129 ;
 wire \i43/i48/n13 ;
 wire \i43/i48/n130 ;
 wire \i43/i48/n131 ;
 wire \i43/i48/n132 ;
 wire \i43/i48/n133 ;
 wire \i43/i48/n134 ;
 wire \i43/i48/n135 ;
 wire \i43/i48/n136 ;
 wire \i43/i48/n137 ;
 wire \i43/i48/n138 ;
 wire \i43/i48/n139 ;
 wire \i43/i48/n14 ;
 wire \i43/i48/n140 ;
 wire \i43/i48/n141 ;
 wire \i43/i48/n142 ;
 wire \i43/i48/n143 ;
 wire \i43/i48/n144 ;
 wire \i43/i48/n145 ;
 wire \i43/i48/n146 ;
 wire \i43/i48/n147 ;
 wire \i43/i48/n148 ;
 wire \i43/i48/n149 ;
 wire \i43/i48/n15 ;
 wire \i43/i48/n150 ;
 wire \i43/i48/n151 ;
 wire \i43/i48/n152 ;
 wire \i43/i48/n153 ;
 wire \i43/i48/n154 ;
 wire \i43/i48/n155 ;
 wire \i43/i48/n156 ;
 wire \i43/i48/n157 ;
 wire \i43/i48/n158 ;
 wire \i43/i48/n159 ;
 wire \i43/i48/n16 ;
 wire \i43/i48/n160 ;
 wire \i43/i48/n161 ;
 wire \i43/i48/n162 ;
 wire \i43/i48/n163 ;
 wire \i43/i48/n164 ;
 wire \i43/i48/n165 ;
 wire \i43/i48/n166 ;
 wire \i43/i48/n167 ;
 wire \i43/i48/n168 ;
 wire \i43/i48/n169 ;
 wire \i43/i48/n17 ;
 wire \i43/i48/n170 ;
 wire \i43/i48/n171 ;
 wire \i43/i48/n172 ;
 wire \i43/i48/n173 ;
 wire \i43/i48/n174 ;
 wire \i43/i48/n175 ;
 wire \i43/i48/n176 ;
 wire \i43/i48/n177 ;
 wire \i43/i48/n178 ;
 wire \i43/i48/n179 ;
 wire \i43/i48/n18 ;
 wire \i43/i48/n180 ;
 wire \i43/i48/n181 ;
 wire \i43/i48/n182 ;
 wire \i43/i48/n183 ;
 wire \i43/i48/n184 ;
 wire \i43/i48/n185 ;
 wire \i43/i48/n186 ;
 wire \i43/i48/n187 ;
 wire \i43/i48/n188 ;
 wire \i43/i48/n189 ;
 wire \i43/i48/n19 ;
 wire \i43/i48/n190 ;
 wire \i43/i48/n191 ;
 wire \i43/i48/n192 ;
 wire \i43/i48/n193 ;
 wire \i43/i48/n194 ;
 wire \i43/i48/n195 ;
 wire \i43/i48/n196 ;
 wire \i43/i48/n197 ;
 wire \i43/i48/n198 ;
 wire \i43/i48/n199 ;
 wire \i43/i48/n2 ;
 wire \i43/i48/n20 ;
 wire \i43/i48/n200 ;
 wire \i43/i48/n201 ;
 wire \i43/i48/n202 ;
 wire \i43/i48/n203 ;
 wire \i43/i48/n204 ;
 wire \i43/i48/n205 ;
 wire \i43/i48/n206 ;
 wire \i43/i48/n207 ;
 wire \i43/i48/n208 ;
 wire \i43/i48/n209 ;
 wire \i43/i48/n21 ;
 wire \i43/i48/n210 ;
 wire \i43/i48/n211 ;
 wire \i43/i48/n212 ;
 wire \i43/i48/n213 ;
 wire \i43/i48/n214 ;
 wire \i43/i48/n215 ;
 wire \i43/i48/n216 ;
 wire \i43/i48/n217 ;
 wire \i43/i48/n218 ;
 wire \i43/i48/n219 ;
 wire \i43/i48/n22 ;
 wire \i43/i48/n220 ;
 wire \i43/i48/n221 ;
 wire \i43/i48/n222 ;
 wire \i43/i48/n223 ;
 wire \i43/i48/n224 ;
 wire \i43/i48/n225 ;
 wire \i43/i48/n226 ;
 wire \i43/i48/n227 ;
 wire \i43/i48/n228 ;
 wire \i43/i48/n229 ;
 wire \i43/i48/n23 ;
 wire \i43/i48/n230 ;
 wire \i43/i48/n231 ;
 wire \i43/i48/n232 ;
 wire \i43/i48/n233 ;
 wire \i43/i48/n234 ;
 wire \i43/i48/n235 ;
 wire \i43/i48/n236 ;
 wire \i43/i48/n237 ;
 wire \i43/i48/n238 ;
 wire \i43/i48/n239 ;
 wire \i43/i48/n24 ;
 wire \i43/i48/n240 ;
 wire \i43/i48/n241 ;
 wire \i43/i48/n242 ;
 wire \i43/i48/n243 ;
 wire \i43/i48/n244 ;
 wire \i43/i48/n245 ;
 wire \i43/i48/n246 ;
 wire \i43/i48/n247 ;
 wire \i43/i48/n248 ;
 wire \i43/i48/n249 ;
 wire \i43/i48/n25 ;
 wire \i43/i48/n250 ;
 wire \i43/i48/n251 ;
 wire \i43/i48/n252 ;
 wire \i43/i48/n253 ;
 wire \i43/i48/n254 ;
 wire \i43/i48/n255 ;
 wire \i43/i48/n256 ;
 wire \i43/i48/n257 ;
 wire \i43/i48/n258 ;
 wire \i43/i48/n259 ;
 wire \i43/i48/n26 ;
 wire \i43/i48/n260 ;
 wire \i43/i48/n261 ;
 wire \i43/i48/n262 ;
 wire \i43/i48/n263 ;
 wire \i43/i48/n264 ;
 wire \i43/i48/n265 ;
 wire \i43/i48/n266 ;
 wire \i43/i48/n267 ;
 wire \i43/i48/n268 ;
 wire \i43/i48/n269 ;
 wire \i43/i48/n27 ;
 wire \i43/i48/n270 ;
 wire \i43/i48/n271 ;
 wire \i43/i48/n272 ;
 wire \i43/i48/n273 ;
 wire \i43/i48/n274 ;
 wire \i43/i48/n275 ;
 wire \i43/i48/n276 ;
 wire \i43/i48/n277 ;
 wire \i43/i48/n278 ;
 wire \i43/i48/n279 ;
 wire \i43/i48/n28 ;
 wire \i43/i48/n280 ;
 wire \i43/i48/n281 ;
 wire \i43/i48/n282 ;
 wire \i43/i48/n283 ;
 wire \i43/i48/n284 ;
 wire \i43/i48/n285 ;
 wire \i43/i48/n286 ;
 wire \i43/i48/n287 ;
 wire \i43/i48/n288 ;
 wire \i43/i48/n289 ;
 wire \i43/i48/n29 ;
 wire \i43/i48/n290 ;
 wire \i43/i48/n291 ;
 wire \i43/i48/n292 ;
 wire \i43/i48/n293 ;
 wire \i43/i48/n294 ;
 wire \i43/i48/n295 ;
 wire \i43/i48/n296 ;
 wire \i43/i48/n297 ;
 wire \i43/i48/n298 ;
 wire \i43/i48/n299 ;
 wire \i43/i48/n3 ;
 wire \i43/i48/n30 ;
 wire \i43/i48/n300 ;
 wire \i43/i48/n301 ;
 wire \i43/i48/n302 ;
 wire \i43/i48/n303 ;
 wire \i43/i48/n304 ;
 wire \i43/i48/n305 ;
 wire \i43/i48/n306 ;
 wire \i43/i48/n307 ;
 wire \i43/i48/n308 ;
 wire \i43/i48/n309 ;
 wire \i43/i48/n31 ;
 wire \i43/i48/n310 ;
 wire \i43/i48/n311 ;
 wire \i43/i48/n312 ;
 wire \i43/i48/n313 ;
 wire \i43/i48/n314 ;
 wire \i43/i48/n315 ;
 wire \i43/i48/n316 ;
 wire \i43/i48/n317 ;
 wire \i43/i48/n318 ;
 wire \i43/i48/n319 ;
 wire \i43/i48/n32 ;
 wire \i43/i48/n320 ;
 wire \i43/i48/n321 ;
 wire \i43/i48/n322 ;
 wire \i43/i48/n323 ;
 wire \i43/i48/n324 ;
 wire \i43/i48/n325 ;
 wire \i43/i48/n326 ;
 wire \i43/i48/n327 ;
 wire \i43/i48/n328 ;
 wire \i43/i48/n329 ;
 wire \i43/i48/n33 ;
 wire \i43/i48/n330 ;
 wire \i43/i48/n331 ;
 wire \i43/i48/n332 ;
 wire \i43/i48/n333 ;
 wire \i43/i48/n334 ;
 wire \i43/i48/n335 ;
 wire \i43/i48/n336 ;
 wire \i43/i48/n337 ;
 wire \i43/i48/n338 ;
 wire \i43/i48/n339 ;
 wire \i43/i48/n34 ;
 wire \i43/i48/n340 ;
 wire \i43/i48/n341 ;
 wire \i43/i48/n342 ;
 wire \i43/i48/n343 ;
 wire \i43/i48/n344 ;
 wire \i43/i48/n345 ;
 wire \i43/i48/n346 ;
 wire \i43/i48/n347 ;
 wire \i43/i48/n348 ;
 wire \i43/i48/n349 ;
 wire \i43/i48/n35 ;
 wire \i43/i48/n350 ;
 wire \i43/i48/n351 ;
 wire \i43/i48/n352 ;
 wire \i43/i48/n353 ;
 wire \i43/i48/n354 ;
 wire \i43/i48/n355 ;
 wire \i43/i48/n356 ;
 wire \i43/i48/n357 ;
 wire \i43/i48/n358 ;
 wire \i43/i48/n359 ;
 wire \i43/i48/n36 ;
 wire \i43/i48/n360 ;
 wire \i43/i48/n361 ;
 wire \i43/i48/n362 ;
 wire \i43/i48/n363 ;
 wire \i43/i48/n364 ;
 wire \i43/i48/n365 ;
 wire \i43/i48/n366 ;
 wire \i43/i48/n367 ;
 wire \i43/i48/n368 ;
 wire \i43/i48/n369 ;
 wire \i43/i48/n37 ;
 wire \i43/i48/n370 ;
 wire \i43/i48/n371 ;
 wire \i43/i48/n372 ;
 wire \i43/i48/n373 ;
 wire \i43/i48/n374 ;
 wire \i43/i48/n375 ;
 wire \i43/i48/n376 ;
 wire \i43/i48/n377 ;
 wire \i43/i48/n378 ;
 wire \i43/i48/n379 ;
 wire \i43/i48/n38 ;
 wire \i43/i48/n380 ;
 wire \i43/i48/n381 ;
 wire \i43/i48/n382 ;
 wire \i43/i48/n383 ;
 wire \i43/i48/n384 ;
 wire \i43/i48/n385 ;
 wire \i43/i48/n386 ;
 wire \i43/i48/n387 ;
 wire \i43/i48/n388 ;
 wire \i43/i48/n389 ;
 wire \i43/i48/n39 ;
 wire \i43/i48/n390 ;
 wire \i43/i48/n391 ;
 wire \i43/i48/n392 ;
 wire \i43/i48/n393 ;
 wire \i43/i48/n394 ;
 wire \i43/i48/n395 ;
 wire \i43/i48/n396 ;
 wire \i43/i48/n397 ;
 wire \i43/i48/n398 ;
 wire \i43/i48/n399 ;
 wire \i43/i48/n4 ;
 wire \i43/i48/n40 ;
 wire \i43/i48/n400 ;
 wire \i43/i48/n401 ;
 wire \i43/i48/n402 ;
 wire \i43/i48/n403 ;
 wire \i43/i48/n404 ;
 wire \i43/i48/n405 ;
 wire \i43/i48/n406 ;
 wire \i43/i48/n407 ;
 wire \i43/i48/n408 ;
 wire \i43/i48/n409 ;
 wire \i43/i48/n41 ;
 wire \i43/i48/n410 ;
 wire \i43/i48/n411 ;
 wire \i43/i48/n412 ;
 wire \i43/i48/n413 ;
 wire \i43/i48/n414 ;
 wire \i43/i48/n415 ;
 wire \i43/i48/n416 ;
 wire \i43/i48/n417 ;
 wire \i43/i48/n418 ;
 wire \i43/i48/n419 ;
 wire \i43/i48/n42 ;
 wire \i43/i48/n420 ;
 wire \i43/i48/n421 ;
 wire \i43/i48/n422 ;
 wire \i43/i48/n423 ;
 wire \i43/i48/n424 ;
 wire \i43/i48/n425 ;
 wire \i43/i48/n426 ;
 wire \i43/i48/n427 ;
 wire \i43/i48/n428 ;
 wire \i43/i48/n429 ;
 wire \i43/i48/n43 ;
 wire \i43/i48/n430 ;
 wire \i43/i48/n431 ;
 wire \i43/i48/n432 ;
 wire \i43/i48/n433 ;
 wire \i43/i48/n434 ;
 wire \i43/i48/n435 ;
 wire \i43/i48/n436 ;
 wire \i43/i48/n437 ;
 wire \i43/i48/n438 ;
 wire \i43/i48/n439 ;
 wire \i43/i48/n44 ;
 wire \i43/i48/n440 ;
 wire \i43/i48/n441 ;
 wire \i43/i48/n442 ;
 wire \i43/i48/n443 ;
 wire \i43/i48/n444 ;
 wire \i43/i48/n445 ;
 wire \i43/i48/n446 ;
 wire \i43/i48/n447 ;
 wire \i43/i48/n448 ;
 wire \i43/i48/n449 ;
 wire \i43/i48/n45 ;
 wire \i43/i48/n450 ;
 wire \i43/i48/n451 ;
 wire \i43/i48/n452 ;
 wire \i43/i48/n453 ;
 wire \i43/i48/n454 ;
 wire \i43/i48/n455 ;
 wire \i43/i48/n456 ;
 wire \i43/i48/n457 ;
 wire \i43/i48/n458 ;
 wire \i43/i48/n459 ;
 wire \i43/i48/n46 ;
 wire \i43/i48/n460 ;
 wire \i43/i48/n461 ;
 wire \i43/i48/n462 ;
 wire \i43/i48/n463 ;
 wire \i43/i48/n464 ;
 wire \i43/i48/n465 ;
 wire \i43/i48/n466 ;
 wire \i43/i48/n467 ;
 wire \i43/i48/n468 ;
 wire \i43/i48/n469 ;
 wire \i43/i48/n47 ;
 wire \i43/i48/n470 ;
 wire \i43/i48/n471 ;
 wire \i43/i48/n472 ;
 wire \i43/i48/n473 ;
 wire \i43/i48/n474 ;
 wire \i43/i48/n475 ;
 wire \i43/i48/n476 ;
 wire \i43/i48/n477 ;
 wire \i43/i48/n478 ;
 wire \i43/i48/n479 ;
 wire \i43/i48/n48 ;
 wire \i43/i48/n480 ;
 wire \i43/i48/n481 ;
 wire \i43/i48/n482 ;
 wire \i43/i48/n483 ;
 wire \i43/i48/n484 ;
 wire \i43/i48/n485 ;
 wire \i43/i48/n486 ;
 wire \i43/i48/n487 ;
 wire \i43/i48/n488 ;
 wire \i43/i48/n489 ;
 wire \i43/i48/n49 ;
 wire \i43/i48/n490 ;
 wire \i43/i48/n491 ;
 wire \i43/i48/n492 ;
 wire \i43/i48/n493 ;
 wire \i43/i48/n494 ;
 wire \i43/i48/n495 ;
 wire \i43/i48/n496 ;
 wire \i43/i48/n497 ;
 wire \i43/i48/n498 ;
 wire \i43/i48/n499 ;
 wire \i43/i48/n5 ;
 wire \i43/i48/n50 ;
 wire \i43/i48/n500 ;
 wire \i43/i48/n501 ;
 wire \i43/i48/n502 ;
 wire \i43/i48/n503 ;
 wire \i43/i48/n504 ;
 wire \i43/i48/n505 ;
 wire \i43/i48/n506 ;
 wire \i43/i48/n507 ;
 wire \i43/i48/n508 ;
 wire \i43/i48/n509 ;
 wire \i43/i48/n51 ;
 wire \i43/i48/n510 ;
 wire \i43/i48/n511 ;
 wire \i43/i48/n512 ;
 wire \i43/i48/n513 ;
 wire \i43/i48/n514 ;
 wire \i43/i48/n52 ;
 wire \i43/i48/n53 ;
 wire \i43/i48/n54 ;
 wire \i43/i48/n55 ;
 wire \i43/i48/n56 ;
 wire \i43/i48/n57 ;
 wire \i43/i48/n58 ;
 wire \i43/i48/n59 ;
 wire \i43/i48/n6 ;
 wire \i43/i48/n60 ;
 wire \i43/i48/n61 ;
 wire \i43/i48/n62 ;
 wire \i43/i48/n63 ;
 wire \i43/i48/n64 ;
 wire \i43/i48/n65 ;
 wire \i43/i48/n66 ;
 wire \i43/i48/n67 ;
 wire \i43/i48/n68 ;
 wire \i43/i48/n69 ;
 wire \i43/i48/n7 ;
 wire \i43/i48/n70 ;
 wire \i43/i48/n71 ;
 wire \i43/i48/n72 ;
 wire \i43/i48/n73 ;
 wire \i43/i48/n74 ;
 wire \i43/i48/n75 ;
 wire \i43/i48/n76 ;
 wire \i43/i48/n77 ;
 wire \i43/i48/n78 ;
 wire \i43/i48/n79 ;
 wire \i43/i48/n8 ;
 wire \i43/i48/n80 ;
 wire \i43/i48/n81 ;
 wire \i43/i48/n82 ;
 wire \i43/i48/n83 ;
 wire \i43/i48/n84 ;
 wire \i43/i48/n85 ;
 wire \i43/i48/n86 ;
 wire \i43/i48/n87 ;
 wire \i43/i48/n88 ;
 wire \i43/i48/n89 ;
 wire \i43/i48/n9 ;
 wire \i43/i48/n90 ;
 wire \i43/i48/n91 ;
 wire \i43/i48/n92 ;
 wire \i43/i48/n93 ;
 wire \i43/i48/n94 ;
 wire \i43/i48/n95 ;
 wire \i43/i48/n96 ;
 wire \i43/i48/n97 ;
 wire \i43/i48/n98 ;
 wire \i43/i48/n99 ;
 wire \i43/i49/n0 ;
 wire \i43/i49/n1 ;
 wire \i43/i49/n10 ;
 wire \i43/i49/n100 ;
 wire \i43/i49/n101 ;
 wire \i43/i49/n102 ;
 wire \i43/i49/n103 ;
 wire \i43/i49/n104 ;
 wire \i43/i49/n105 ;
 wire \i43/i49/n106 ;
 wire \i43/i49/n107 ;
 wire \i43/i49/n108 ;
 wire \i43/i49/n109 ;
 wire \i43/i49/n11 ;
 wire \i43/i49/n110 ;
 wire \i43/i49/n111 ;
 wire \i43/i49/n112 ;
 wire \i43/i49/n113 ;
 wire \i43/i49/n114 ;
 wire \i43/i49/n115 ;
 wire \i43/i49/n116 ;
 wire \i43/i49/n117 ;
 wire \i43/i49/n118 ;
 wire \i43/i49/n119 ;
 wire \i43/i49/n12 ;
 wire \i43/i49/n120 ;
 wire \i43/i49/n121 ;
 wire \i43/i49/n122 ;
 wire \i43/i49/n123 ;
 wire \i43/i49/n124 ;
 wire \i43/i49/n125 ;
 wire \i43/i49/n126 ;
 wire \i43/i49/n127 ;
 wire \i43/i49/n128 ;
 wire \i43/i49/n129 ;
 wire \i43/i49/n13 ;
 wire \i43/i49/n130 ;
 wire \i43/i49/n131 ;
 wire \i43/i49/n132 ;
 wire \i43/i49/n133 ;
 wire \i43/i49/n134 ;
 wire \i43/i49/n135 ;
 wire \i43/i49/n136 ;
 wire \i43/i49/n137 ;
 wire \i43/i49/n138 ;
 wire \i43/i49/n139 ;
 wire \i43/i49/n14 ;
 wire \i43/i49/n140 ;
 wire \i43/i49/n141 ;
 wire \i43/i49/n142 ;
 wire \i43/i49/n143 ;
 wire \i43/i49/n144 ;
 wire \i43/i49/n145 ;
 wire \i43/i49/n146 ;
 wire \i43/i49/n147 ;
 wire \i43/i49/n148 ;
 wire \i43/i49/n149 ;
 wire \i43/i49/n15 ;
 wire \i43/i49/n150 ;
 wire \i43/i49/n151 ;
 wire \i43/i49/n152 ;
 wire \i43/i49/n153 ;
 wire \i43/i49/n154 ;
 wire \i43/i49/n155 ;
 wire \i43/i49/n156 ;
 wire \i43/i49/n157 ;
 wire \i43/i49/n158 ;
 wire \i43/i49/n159 ;
 wire \i43/i49/n16 ;
 wire \i43/i49/n160 ;
 wire \i43/i49/n161 ;
 wire \i43/i49/n162 ;
 wire \i43/i49/n163 ;
 wire \i43/i49/n164 ;
 wire \i43/i49/n165 ;
 wire \i43/i49/n166 ;
 wire \i43/i49/n167 ;
 wire \i43/i49/n168 ;
 wire \i43/i49/n169 ;
 wire \i43/i49/n17 ;
 wire \i43/i49/n170 ;
 wire \i43/i49/n171 ;
 wire \i43/i49/n172 ;
 wire \i43/i49/n173 ;
 wire \i43/i49/n174 ;
 wire \i43/i49/n175 ;
 wire \i43/i49/n176 ;
 wire \i43/i49/n177 ;
 wire \i43/i49/n178 ;
 wire \i43/i49/n179 ;
 wire \i43/i49/n18 ;
 wire \i43/i49/n180 ;
 wire \i43/i49/n181 ;
 wire \i43/i49/n182 ;
 wire \i43/i49/n183 ;
 wire \i43/i49/n184 ;
 wire \i43/i49/n185 ;
 wire \i43/i49/n186 ;
 wire \i43/i49/n187 ;
 wire \i43/i49/n188 ;
 wire \i43/i49/n189 ;
 wire \i43/i49/n19 ;
 wire \i43/i49/n190 ;
 wire \i43/i49/n191 ;
 wire \i43/i49/n192 ;
 wire \i43/i49/n193 ;
 wire \i43/i49/n194 ;
 wire \i43/i49/n195 ;
 wire \i43/i49/n196 ;
 wire \i43/i49/n197 ;
 wire \i43/i49/n198 ;
 wire \i43/i49/n199 ;
 wire \i43/i49/n2 ;
 wire \i43/i49/n20 ;
 wire \i43/i49/n200 ;
 wire \i43/i49/n201 ;
 wire \i43/i49/n202 ;
 wire \i43/i49/n203 ;
 wire \i43/i49/n204 ;
 wire \i43/i49/n205 ;
 wire \i43/i49/n206 ;
 wire \i43/i49/n207 ;
 wire \i43/i49/n208 ;
 wire \i43/i49/n209 ;
 wire \i43/i49/n21 ;
 wire \i43/i49/n210 ;
 wire \i43/i49/n211 ;
 wire \i43/i49/n212 ;
 wire \i43/i49/n213 ;
 wire \i43/i49/n214 ;
 wire \i43/i49/n215 ;
 wire \i43/i49/n216 ;
 wire \i43/i49/n217 ;
 wire \i43/i49/n218 ;
 wire \i43/i49/n219 ;
 wire \i43/i49/n22 ;
 wire \i43/i49/n220 ;
 wire \i43/i49/n221 ;
 wire \i43/i49/n222 ;
 wire \i43/i49/n223 ;
 wire \i43/i49/n224 ;
 wire \i43/i49/n225 ;
 wire \i43/i49/n226 ;
 wire \i43/i49/n227 ;
 wire \i43/i49/n228 ;
 wire \i43/i49/n229 ;
 wire \i43/i49/n23 ;
 wire \i43/i49/n230 ;
 wire \i43/i49/n231 ;
 wire \i43/i49/n232 ;
 wire \i43/i49/n233 ;
 wire \i43/i49/n234 ;
 wire \i43/i49/n235 ;
 wire \i43/i49/n236 ;
 wire \i43/i49/n237 ;
 wire \i43/i49/n238 ;
 wire \i43/i49/n239 ;
 wire \i43/i49/n24 ;
 wire \i43/i49/n240 ;
 wire \i43/i49/n241 ;
 wire \i43/i49/n242 ;
 wire \i43/i49/n243 ;
 wire \i43/i49/n244 ;
 wire \i43/i49/n245 ;
 wire \i43/i49/n246 ;
 wire \i43/i49/n247 ;
 wire \i43/i49/n248 ;
 wire \i43/i49/n249 ;
 wire \i43/i49/n25 ;
 wire \i43/i49/n250 ;
 wire \i43/i49/n251 ;
 wire \i43/i49/n252 ;
 wire \i43/i49/n253 ;
 wire \i43/i49/n254 ;
 wire \i43/i49/n255 ;
 wire \i43/i49/n256 ;
 wire \i43/i49/n257 ;
 wire \i43/i49/n258 ;
 wire \i43/i49/n259 ;
 wire \i43/i49/n26 ;
 wire \i43/i49/n260 ;
 wire \i43/i49/n261 ;
 wire \i43/i49/n262 ;
 wire \i43/i49/n263 ;
 wire \i43/i49/n264 ;
 wire \i43/i49/n265 ;
 wire \i43/i49/n266 ;
 wire \i43/i49/n267 ;
 wire \i43/i49/n268 ;
 wire \i43/i49/n269 ;
 wire \i43/i49/n27 ;
 wire \i43/i49/n270 ;
 wire \i43/i49/n271 ;
 wire \i43/i49/n272 ;
 wire \i43/i49/n273 ;
 wire \i43/i49/n274 ;
 wire \i43/i49/n275 ;
 wire \i43/i49/n276 ;
 wire \i43/i49/n277 ;
 wire \i43/i49/n278 ;
 wire \i43/i49/n279 ;
 wire \i43/i49/n28 ;
 wire \i43/i49/n280 ;
 wire \i43/i49/n281 ;
 wire \i43/i49/n282 ;
 wire \i43/i49/n283 ;
 wire \i43/i49/n284 ;
 wire \i43/i49/n285 ;
 wire \i43/i49/n286 ;
 wire \i43/i49/n287 ;
 wire \i43/i49/n288 ;
 wire \i43/i49/n289 ;
 wire \i43/i49/n29 ;
 wire \i43/i49/n290 ;
 wire \i43/i49/n291 ;
 wire \i43/i49/n292 ;
 wire \i43/i49/n293 ;
 wire \i43/i49/n294 ;
 wire \i43/i49/n295 ;
 wire \i43/i49/n296 ;
 wire \i43/i49/n297 ;
 wire \i43/i49/n298 ;
 wire \i43/i49/n299 ;
 wire \i43/i49/n3 ;
 wire \i43/i49/n30 ;
 wire \i43/i49/n300 ;
 wire \i43/i49/n301 ;
 wire \i43/i49/n302 ;
 wire \i43/i49/n303 ;
 wire \i43/i49/n304 ;
 wire \i43/i49/n305 ;
 wire \i43/i49/n306 ;
 wire \i43/i49/n307 ;
 wire \i43/i49/n308 ;
 wire \i43/i49/n309 ;
 wire \i43/i49/n31 ;
 wire \i43/i49/n310 ;
 wire \i43/i49/n311 ;
 wire \i43/i49/n312 ;
 wire \i43/i49/n313 ;
 wire \i43/i49/n314 ;
 wire \i43/i49/n315 ;
 wire \i43/i49/n316 ;
 wire \i43/i49/n317 ;
 wire \i43/i49/n318 ;
 wire \i43/i49/n319 ;
 wire \i43/i49/n32 ;
 wire \i43/i49/n320 ;
 wire \i43/i49/n321 ;
 wire \i43/i49/n322 ;
 wire \i43/i49/n323 ;
 wire \i43/i49/n324 ;
 wire \i43/i49/n325 ;
 wire \i43/i49/n326 ;
 wire \i43/i49/n327 ;
 wire \i43/i49/n328 ;
 wire \i43/i49/n329 ;
 wire \i43/i49/n33 ;
 wire \i43/i49/n330 ;
 wire \i43/i49/n331 ;
 wire \i43/i49/n332 ;
 wire \i43/i49/n333 ;
 wire \i43/i49/n334 ;
 wire \i43/i49/n335 ;
 wire \i43/i49/n336 ;
 wire \i43/i49/n337 ;
 wire \i43/i49/n338 ;
 wire \i43/i49/n339 ;
 wire \i43/i49/n34 ;
 wire \i43/i49/n340 ;
 wire \i43/i49/n341 ;
 wire \i43/i49/n342 ;
 wire \i43/i49/n343 ;
 wire \i43/i49/n344 ;
 wire \i43/i49/n345 ;
 wire \i43/i49/n346 ;
 wire \i43/i49/n347 ;
 wire \i43/i49/n348 ;
 wire \i43/i49/n349 ;
 wire \i43/i49/n35 ;
 wire \i43/i49/n350 ;
 wire \i43/i49/n351 ;
 wire \i43/i49/n352 ;
 wire \i43/i49/n353 ;
 wire \i43/i49/n354 ;
 wire \i43/i49/n355 ;
 wire \i43/i49/n356 ;
 wire \i43/i49/n357 ;
 wire \i43/i49/n358 ;
 wire \i43/i49/n359 ;
 wire \i43/i49/n36 ;
 wire \i43/i49/n360 ;
 wire \i43/i49/n361 ;
 wire \i43/i49/n362 ;
 wire \i43/i49/n363 ;
 wire \i43/i49/n364 ;
 wire \i43/i49/n365 ;
 wire \i43/i49/n366 ;
 wire \i43/i49/n367 ;
 wire \i43/i49/n368 ;
 wire \i43/i49/n369 ;
 wire \i43/i49/n37 ;
 wire \i43/i49/n370 ;
 wire \i43/i49/n371 ;
 wire \i43/i49/n372 ;
 wire \i43/i49/n373 ;
 wire \i43/i49/n374 ;
 wire \i43/i49/n375 ;
 wire \i43/i49/n376 ;
 wire \i43/i49/n377 ;
 wire \i43/i49/n378 ;
 wire \i43/i49/n379 ;
 wire \i43/i49/n38 ;
 wire \i43/i49/n380 ;
 wire \i43/i49/n381 ;
 wire \i43/i49/n382 ;
 wire \i43/i49/n383 ;
 wire \i43/i49/n384 ;
 wire \i43/i49/n385 ;
 wire \i43/i49/n386 ;
 wire \i43/i49/n387 ;
 wire \i43/i49/n388 ;
 wire \i43/i49/n389 ;
 wire \i43/i49/n39 ;
 wire \i43/i49/n390 ;
 wire \i43/i49/n391 ;
 wire \i43/i49/n392 ;
 wire \i43/i49/n393 ;
 wire \i43/i49/n394 ;
 wire \i43/i49/n395 ;
 wire \i43/i49/n396 ;
 wire \i43/i49/n397 ;
 wire \i43/i49/n398 ;
 wire \i43/i49/n399 ;
 wire \i43/i49/n4 ;
 wire \i43/i49/n40 ;
 wire \i43/i49/n400 ;
 wire \i43/i49/n401 ;
 wire \i43/i49/n402 ;
 wire \i43/i49/n403 ;
 wire \i43/i49/n404 ;
 wire \i43/i49/n405 ;
 wire \i43/i49/n406 ;
 wire \i43/i49/n407 ;
 wire \i43/i49/n408 ;
 wire \i43/i49/n409 ;
 wire \i43/i49/n41 ;
 wire \i43/i49/n410 ;
 wire \i43/i49/n411 ;
 wire \i43/i49/n412 ;
 wire \i43/i49/n413 ;
 wire \i43/i49/n414 ;
 wire \i43/i49/n415 ;
 wire \i43/i49/n416 ;
 wire \i43/i49/n417 ;
 wire \i43/i49/n418 ;
 wire \i43/i49/n419 ;
 wire \i43/i49/n42 ;
 wire \i43/i49/n420 ;
 wire \i43/i49/n421 ;
 wire \i43/i49/n422 ;
 wire \i43/i49/n423 ;
 wire \i43/i49/n424 ;
 wire \i43/i49/n425 ;
 wire \i43/i49/n426 ;
 wire \i43/i49/n427 ;
 wire \i43/i49/n428 ;
 wire \i43/i49/n429 ;
 wire \i43/i49/n43 ;
 wire \i43/i49/n430 ;
 wire \i43/i49/n431 ;
 wire \i43/i49/n432 ;
 wire \i43/i49/n433 ;
 wire \i43/i49/n434 ;
 wire \i43/i49/n435 ;
 wire \i43/i49/n436 ;
 wire \i43/i49/n437 ;
 wire \i43/i49/n438 ;
 wire \i43/i49/n439 ;
 wire \i43/i49/n44 ;
 wire \i43/i49/n440 ;
 wire \i43/i49/n441 ;
 wire \i43/i49/n442 ;
 wire \i43/i49/n443 ;
 wire \i43/i49/n444 ;
 wire \i43/i49/n445 ;
 wire \i43/i49/n446 ;
 wire \i43/i49/n447 ;
 wire \i43/i49/n448 ;
 wire \i43/i49/n449 ;
 wire \i43/i49/n45 ;
 wire \i43/i49/n450 ;
 wire \i43/i49/n451 ;
 wire \i43/i49/n452 ;
 wire \i43/i49/n453 ;
 wire \i43/i49/n454 ;
 wire \i43/i49/n455 ;
 wire \i43/i49/n456 ;
 wire \i43/i49/n457 ;
 wire \i43/i49/n458 ;
 wire \i43/i49/n459 ;
 wire \i43/i49/n46 ;
 wire \i43/i49/n460 ;
 wire \i43/i49/n461 ;
 wire \i43/i49/n462 ;
 wire \i43/i49/n463 ;
 wire \i43/i49/n464 ;
 wire \i43/i49/n465 ;
 wire \i43/i49/n466 ;
 wire \i43/i49/n467 ;
 wire \i43/i49/n468 ;
 wire \i43/i49/n469 ;
 wire \i43/i49/n47 ;
 wire \i43/i49/n470 ;
 wire \i43/i49/n471 ;
 wire \i43/i49/n472 ;
 wire \i43/i49/n473 ;
 wire \i43/i49/n474 ;
 wire \i43/i49/n475 ;
 wire \i43/i49/n476 ;
 wire \i43/i49/n477 ;
 wire \i43/i49/n478 ;
 wire \i43/i49/n479 ;
 wire \i43/i49/n48 ;
 wire \i43/i49/n480 ;
 wire \i43/i49/n481 ;
 wire \i43/i49/n482 ;
 wire \i43/i49/n483 ;
 wire \i43/i49/n484 ;
 wire \i43/i49/n485 ;
 wire \i43/i49/n486 ;
 wire \i43/i49/n487 ;
 wire \i43/i49/n488 ;
 wire \i43/i49/n489 ;
 wire \i43/i49/n49 ;
 wire \i43/i49/n490 ;
 wire \i43/i49/n491 ;
 wire \i43/i49/n492 ;
 wire \i43/i49/n493 ;
 wire \i43/i49/n494 ;
 wire \i43/i49/n495 ;
 wire \i43/i49/n496 ;
 wire \i43/i49/n497 ;
 wire \i43/i49/n498 ;
 wire \i43/i49/n499 ;
 wire \i43/i49/n5 ;
 wire \i43/i49/n50 ;
 wire \i43/i49/n500 ;
 wire \i43/i49/n501 ;
 wire \i43/i49/n502 ;
 wire \i43/i49/n503 ;
 wire \i43/i49/n504 ;
 wire \i43/i49/n505 ;
 wire \i43/i49/n506 ;
 wire \i43/i49/n507 ;
 wire \i43/i49/n508 ;
 wire \i43/i49/n509 ;
 wire \i43/i49/n51 ;
 wire \i43/i49/n510 ;
 wire \i43/i49/n511 ;
 wire \i43/i49/n512 ;
 wire \i43/i49/n513 ;
 wire \i43/i49/n514 ;
 wire \i43/i49/n52 ;
 wire \i43/i49/n53 ;
 wire \i43/i49/n54 ;
 wire \i43/i49/n55 ;
 wire \i43/i49/n56 ;
 wire \i43/i49/n57 ;
 wire \i43/i49/n58 ;
 wire \i43/i49/n59 ;
 wire \i43/i49/n6 ;
 wire \i43/i49/n60 ;
 wire \i43/i49/n61 ;
 wire \i43/i49/n62 ;
 wire \i43/i49/n63 ;
 wire \i43/i49/n64 ;
 wire \i43/i49/n65 ;
 wire \i43/i49/n66 ;
 wire \i43/i49/n67 ;
 wire \i43/i49/n68 ;
 wire \i43/i49/n69 ;
 wire \i43/i49/n7 ;
 wire \i43/i49/n70 ;
 wire \i43/i49/n71 ;
 wire \i43/i49/n72 ;
 wire \i43/i49/n73 ;
 wire \i43/i49/n74 ;
 wire \i43/i49/n75 ;
 wire \i43/i49/n76 ;
 wire \i43/i49/n77 ;
 wire \i43/i49/n78 ;
 wire \i43/i49/n79 ;
 wire \i43/i49/n8 ;
 wire \i43/i49/n80 ;
 wire \i43/i49/n81 ;
 wire \i43/i49/n82 ;
 wire \i43/i49/n83 ;
 wire \i43/i49/n84 ;
 wire \i43/i49/n85 ;
 wire \i43/i49/n86 ;
 wire \i43/i49/n87 ;
 wire \i43/i49/n88 ;
 wire \i43/i49/n89 ;
 wire \i43/i49/n9 ;
 wire \i43/i49/n90 ;
 wire \i43/i49/n91 ;
 wire \i43/i49/n92 ;
 wire \i43/i49/n93 ;
 wire \i43/i49/n94 ;
 wire \i43/i49/n95 ;
 wire \i43/i49/n96 ;
 wire \i43/i49/n97 ;
 wire \i43/i49/n98 ;
 wire \i43/i49/n99 ;
 wire \i44/n0 ;
 wire \i44/n1 ;
 wire \i44/n10 ;
 wire \i44/n100 ;
 wire \i44/n101 ;
 wire \i44/n102 ;
 wire \i44/n103 ;
 wire \i44/n104 ;
 wire \i44/n105 ;
 wire \i44/n106 ;
 wire \i44/n107 ;
 wire \i44/n108 ;
 wire \i44/n109 ;
 wire \i44/n11 ;
 wire \i44/n110 ;
 wire \i44/n111 ;
 wire \i44/n112 ;
 wire \i44/n113 ;
 wire \i44/n114 ;
 wire \i44/n115 ;
 wire \i44/n116 ;
 wire \i44/n117 ;
 wire \i44/n118 ;
 wire \i44/n119 ;
 wire \i44/n12 ;
 wire \i44/n120 ;
 wire \i44/n121 ;
 wire \i44/n122 ;
 wire \i44/n123 ;
 wire \i44/n124 ;
 wire \i44/n125 ;
 wire \i44/n126 ;
 wire \i44/n127 ;
 wire \i44/n128 ;
 wire \i44/n129 ;
 wire \i44/n13 ;
 wire \i44/n130 ;
 wire \i44/n131 ;
 wire \i44/n132 ;
 wire \i44/n133 ;
 wire \i44/n134 ;
 wire \i44/n135 ;
 wire \i44/n136 ;
 wire \i44/n137 ;
 wire \i44/n138 ;
 wire \i44/n139 ;
 wire \i44/n14 ;
 wire \i44/n140 ;
 wire \i44/n141 ;
 wire \i44/n142 ;
 wire \i44/n143 ;
 wire \i44/n144 ;
 wire \i44/n145 ;
 wire \i44/n146 ;
 wire \i44/n147 ;
 wire \i44/n148 ;
 wire \i44/n149 ;
 wire \i44/n15 ;
 wire \i44/n150 ;
 wire \i44/n151 ;
 wire \i44/n152 ;
 wire \i44/n153 ;
 wire \i44/n154 ;
 wire \i44/n155 ;
 wire \i44/n156 ;
 wire \i44/n157 ;
 wire \i44/n158 ;
 wire \i44/n159 ;
 wire \i44/n16 ;
 wire \i44/n160 ;
 wire \i44/n161 ;
 wire \i44/n162 ;
 wire \i44/n163 ;
 wire \i44/n164 ;
 wire \i44/n165 ;
 wire \i44/n166 ;
 wire \i44/n167 ;
 wire \i44/n168 ;
 wire \i44/n169 ;
 wire \i44/n17 ;
 wire \i44/n170 ;
 wire \i44/n171 ;
 wire \i44/n172 ;
 wire \i44/n173 ;
 wire \i44/n174 ;
 wire \i44/n175 ;
 wire \i44/n176 ;
 wire \i44/n177 ;
 wire \i44/n178 ;
 wire \i44/n179 ;
 wire \i44/n18 ;
 wire \i44/n180 ;
 wire \i44/n181 ;
 wire \i44/n182 ;
 wire \i44/n183 ;
 wire \i44/n184 ;
 wire \i44/n185 ;
 wire \i44/n186 ;
 wire \i44/n187 ;
 wire \i44/n188 ;
 wire \i44/n189 ;
 wire \i44/n19 ;
 wire \i44/n190 ;
 wire \i44/n191 ;
 wire \i44/n192 ;
 wire \i44/n193 ;
 wire \i44/n194 ;
 wire \i44/n195 ;
 wire \i44/n196 ;
 wire \i44/n197 ;
 wire \i44/n198 ;
 wire \i44/n199 ;
 wire \i44/n2 ;
 wire \i44/n20 ;
 wire \i44/n200 ;
 wire \i44/n201 ;
 wire \i44/n202 ;
 wire \i44/n203 ;
 wire \i44/n204 ;
 wire \i44/n205 ;
 wire \i44/n206 ;
 wire \i44/n207 ;
 wire \i44/n208 ;
 wire \i44/n209 ;
 wire \i44/n21 ;
 wire \i44/n210 ;
 wire \i44/n211 ;
 wire \i44/n212 ;
 wire \i44/n213 ;
 wire \i44/n214 ;
 wire \i44/n215 ;
 wire \i44/n216 ;
 wire \i44/n217 ;
 wire \i44/n218 ;
 wire \i44/n219 ;
 wire \i44/n22 ;
 wire \i44/n220 ;
 wire \i44/n221 ;
 wire \i44/n222 ;
 wire \i44/n223 ;
 wire \i44/n224 ;
 wire \i44/n225 ;
 wire \i44/n226 ;
 wire \i44/n227 ;
 wire \i44/n228 ;
 wire \i44/n229 ;
 wire \i44/n23 ;
 wire \i44/n230 ;
 wire \i44/n231 ;
 wire \i44/n232 ;
 wire \i44/n233 ;
 wire \i44/n234 ;
 wire \i44/n235 ;
 wire \i44/n236 ;
 wire \i44/n237 ;
 wire \i44/n238 ;
 wire \i44/n239 ;
 wire \i44/n24 ;
 wire \i44/n240 ;
 wire \i44/n241 ;
 wire \i44/n242 ;
 wire \i44/n243 ;
 wire \i44/n244 ;
 wire \i44/n245 ;
 wire \i44/n246 ;
 wire \i44/n247 ;
 wire \i44/n248 ;
 wire \i44/n249 ;
 wire \i44/n25 ;
 wire \i44/n250 ;
 wire \i44/n251 ;
 wire \i44/n252 ;
 wire \i44/n253 ;
 wire \i44/n254 ;
 wire \i44/n255 ;
 wire \i44/n256 ;
 wire \i44/n257 ;
 wire \i44/n258 ;
 wire \i44/n259 ;
 wire \i44/n26 ;
 wire \i44/n260 ;
 wire \i44/n261 ;
 wire \i44/n262 ;
 wire \i44/n263 ;
 wire \i44/n264 ;
 wire \i44/n265 ;
 wire \i44/n266 ;
 wire \i44/n267 ;
 wire \i44/n268 ;
 wire \i44/n269 ;
 wire \i44/n27 ;
 wire \i44/n270 ;
 wire \i44/n271 ;
 wire \i44/n272 ;
 wire \i44/n273 ;
 wire \i44/n274 ;
 wire \i44/n275 ;
 wire \i44/n276 ;
 wire \i44/n277 ;
 wire \i44/n278 ;
 wire \i44/n279 ;
 wire \i44/n28 ;
 wire \i44/n280 ;
 wire \i44/n281 ;
 wire \i44/n282 ;
 wire \i44/n283 ;
 wire \i44/n284 ;
 wire \i44/n285 ;
 wire \i44/n286 ;
 wire \i44/n287 ;
 wire \i44/n288 ;
 wire \i44/n289 ;
 wire \i44/n29 ;
 wire \i44/n290 ;
 wire \i44/n291 ;
 wire \i44/n292 ;
 wire \i44/n293 ;
 wire \i44/n294 ;
 wire \i44/n295 ;
 wire \i44/n296 ;
 wire \i44/n297 ;
 wire \i44/n298 ;
 wire \i44/n299 ;
 wire \i44/n3 ;
 wire \i44/n30 ;
 wire \i44/n300 ;
 wire \i44/n301 ;
 wire \i44/n302 ;
 wire \i44/n303 ;
 wire \i44/n304 ;
 wire \i44/n305 ;
 wire \i44/n306 ;
 wire \i44/n307 ;
 wire \i44/n308 ;
 wire \i44/n309 ;
 wire \i44/n31 ;
 wire \i44/n310 ;
 wire \i44/n311 ;
 wire \i44/n312 ;
 wire \i44/n313 ;
 wire \i44/n314 ;
 wire \i44/n315 ;
 wire \i44/n316 ;
 wire \i44/n317 ;
 wire \i44/n318 ;
 wire \i44/n319 ;
 wire \i44/n32 ;
 wire \i44/n320 ;
 wire \i44/n321 ;
 wire \i44/n322 ;
 wire \i44/n323 ;
 wire \i44/n324 ;
 wire \i44/n325 ;
 wire \i44/n326 ;
 wire \i44/n327 ;
 wire \i44/n328 ;
 wire \i44/n329 ;
 wire \i44/n33 ;
 wire \i44/n330 ;
 wire \i44/n331 ;
 wire \i44/n332 ;
 wire \i44/n333 ;
 wire \i44/n334 ;
 wire \i44/n335 ;
 wire \i44/n336 ;
 wire \i44/n337 ;
 wire \i44/n338 ;
 wire \i44/n339 ;
 wire \i44/n34 ;
 wire \i44/n340 ;
 wire \i44/n341 ;
 wire \i44/n342 ;
 wire \i44/n343 ;
 wire \i44/n344 ;
 wire \i44/n345 ;
 wire \i44/n346 ;
 wire \i44/n347 ;
 wire \i44/n348 ;
 wire \i44/n349 ;
 wire \i44/n35 ;
 wire \i44/n350 ;
 wire \i44/n351 ;
 wire \i44/n352 ;
 wire \i44/n353 ;
 wire \i44/n354 ;
 wire \i44/n355 ;
 wire \i44/n356 ;
 wire \i44/n357 ;
 wire \i44/n358 ;
 wire \i44/n359 ;
 wire \i44/n36 ;
 wire \i44/n360 ;
 wire \i44/n361 ;
 wire \i44/n362 ;
 wire \i44/n363 ;
 wire \i44/n364 ;
 wire \i44/n365 ;
 wire \i44/n366 ;
 wire \i44/n367 ;
 wire \i44/n368 ;
 wire \i44/n369 ;
 wire \i44/n37 ;
 wire \i44/n370 ;
 wire \i44/n371 ;
 wire \i44/n372 ;
 wire \i44/n373 ;
 wire \i44/n374 ;
 wire \i44/n375 ;
 wire \i44/n376 ;
 wire \i44/n377 ;
 wire \i44/n378 ;
 wire \i44/n379 ;
 wire \i44/n38 ;
 wire \i44/n380 ;
 wire \i44/n381 ;
 wire \i44/n382 ;
 wire \i44/n383 ;
 wire \i44/n384 ;
 wire \i44/n385 ;
 wire \i44/n386 ;
 wire \i44/n387 ;
 wire \i44/n388 ;
 wire \i44/n389 ;
 wire \i44/n39 ;
 wire \i44/n390 ;
 wire \i44/n391 ;
 wire \i44/n392 ;
 wire \i44/n393 ;
 wire \i44/n394 ;
 wire \i44/n395 ;
 wire \i44/n396 ;
 wire \i44/n397 ;
 wire \i44/n398 ;
 wire \i44/n399 ;
 wire \i44/n4 ;
 wire \i44/n40 ;
 wire \i44/n400 ;
 wire \i44/n401 ;
 wire \i44/n402 ;
 wire \i44/n403 ;
 wire \i44/n404 ;
 wire \i44/n405 ;
 wire \i44/n406 ;
 wire \i44/n407 ;
 wire \i44/n408 ;
 wire \i44/n409 ;
 wire \i44/n41 ;
 wire \i44/n410 ;
 wire \i44/n411 ;
 wire \i44/n412 ;
 wire \i44/n413 ;
 wire \i44/n414 ;
 wire \i44/n415 ;
 wire \i44/n416 ;
 wire \i44/n417 ;
 wire \i44/n418 ;
 wire \i44/n419 ;
 wire \i44/n42 ;
 wire \i44/n420 ;
 wire \i44/n421 ;
 wire \i44/n422 ;
 wire \i44/n423 ;
 wire \i44/n424 ;
 wire \i44/n425 ;
 wire \i44/n426 ;
 wire \i44/n427 ;
 wire \i44/n428 ;
 wire \i44/n429 ;
 wire \i44/n43 ;
 wire \i44/n430 ;
 wire \i44/n431 ;
 wire \i44/n432 ;
 wire \i44/n433 ;
 wire \i44/n434 ;
 wire \i44/n435 ;
 wire \i44/n436 ;
 wire \i44/n437 ;
 wire \i44/n438 ;
 wire \i44/n439 ;
 wire \i44/n44 ;
 wire \i44/n440 ;
 wire \i44/n441 ;
 wire \i44/n442 ;
 wire \i44/n443 ;
 wire \i44/n444 ;
 wire \i44/n445 ;
 wire \i44/n446 ;
 wire \i44/n447 ;
 wire \i44/n448 ;
 wire \i44/n449 ;
 wire \i44/n45 ;
 wire \i44/n450 ;
 wire \i44/n451 ;
 wire \i44/n452 ;
 wire \i44/n453 ;
 wire \i44/n454 ;
 wire \i44/n455 ;
 wire \i44/n456 ;
 wire \i44/n457 ;
 wire \i44/n458 ;
 wire \i44/n459 ;
 wire \i44/n46 ;
 wire \i44/n460 ;
 wire \i44/n461 ;
 wire \i44/n462 ;
 wire \i44/n463 ;
 wire \i44/n464 ;
 wire \i44/n465 ;
 wire \i44/n466 ;
 wire \i44/n467 ;
 wire \i44/n468 ;
 wire \i44/n469 ;
 wire \i44/n47 ;
 wire \i44/n470 ;
 wire \i44/n471 ;
 wire \i44/n472 ;
 wire \i44/n473 ;
 wire \i44/n474 ;
 wire \i44/n475 ;
 wire \i44/n476 ;
 wire \i44/n477 ;
 wire \i44/n478 ;
 wire \i44/n479 ;
 wire \i44/n48 ;
 wire \i44/n480 ;
 wire \i44/n481 ;
 wire \i44/n482 ;
 wire \i44/n483 ;
 wire \i44/n484 ;
 wire \i44/n485 ;
 wire \i44/n486 ;
 wire \i44/n487 ;
 wire \i44/n488 ;
 wire \i44/n489 ;
 wire \i44/n49 ;
 wire \i44/n490 ;
 wire \i44/n491 ;
 wire \i44/n492 ;
 wire \i44/n493 ;
 wire \i44/n494 ;
 wire \i44/n495 ;
 wire \i44/n496 ;
 wire \i44/n497 ;
 wire \i44/n498 ;
 wire \i44/n499 ;
 wire \i44/n5 ;
 wire \i44/n50 ;
 wire \i44/n500 ;
 wire \i44/n501 ;
 wire \i44/n502 ;
 wire \i44/n503 ;
 wire \i44/n504 ;
 wire \i44/n505 ;
 wire \i44/n506 ;
 wire \i44/n507 ;
 wire \i44/n508 ;
 wire \i44/n509 ;
 wire \i44/n51 ;
 wire \i44/n510 ;
 wire \i44/n511 ;
 wire \i44/n512 ;
 wire \i44/n513 ;
 wire \i44/n514 ;
 wire \i44/n515 ;
 wire \i44/n516 ;
 wire \i44/n517 ;
 wire \i44/n518 ;
 wire \i44/n519 ;
 wire \i44/n52 ;
 wire \i44/n520 ;
 wire \i44/n521 ;
 wire \i44/n522 ;
 wire \i44/n523 ;
 wire \i44/n524 ;
 wire \i44/n525 ;
 wire \i44/n526 ;
 wire \i44/n527 ;
 wire \i44/n528 ;
 wire \i44/n529 ;
 wire \i44/n53 ;
 wire \i44/n530 ;
 wire \i44/n531 ;
 wire \i44/n532 ;
 wire \i44/n533 ;
 wire \i44/n534 ;
 wire \i44/n535 ;
 wire \i44/n536 ;
 wire \i44/n537 ;
 wire \i44/n538 ;
 wire \i44/n539 ;
 wire \i44/n54 ;
 wire \i44/n540 ;
 wire \i44/n541 ;
 wire \i44/n542 ;
 wire \i44/n543 ;
 wire \i44/n544 ;
 wire \i44/n545 ;
 wire \i44/n546 ;
 wire \i44/n547 ;
 wire \i44/n548 ;
 wire \i44/n549 ;
 wire \i44/n55 ;
 wire \i44/n550 ;
 wire \i44/n551 ;
 wire \i44/n552 ;
 wire \i44/n553 ;
 wire \i44/n554 ;
 wire \i44/n555 ;
 wire \i44/n556 ;
 wire \i44/n557 ;
 wire \i44/n558 ;
 wire \i44/n559 ;
 wire \i44/n56 ;
 wire \i44/n560 ;
 wire \i44/n561 ;
 wire \i44/n562 ;
 wire \i44/n563 ;
 wire \i44/n564 ;
 wire \i44/n565 ;
 wire \i44/n566 ;
 wire \i44/n567 ;
 wire \i44/n568 ;
 wire \i44/n569 ;
 wire \i44/n57 ;
 wire \i44/n570 ;
 wire \i44/n571 ;
 wire \i44/n572 ;
 wire \i44/n573 ;
 wire \i44/n574 ;
 wire \i44/n575 ;
 wire \i44/n576 ;
 wire \i44/n577 ;
 wire \i44/n578 ;
 wire \i44/n579 ;
 wire \i44/n58 ;
 wire \i44/n580 ;
 wire \i44/n581 ;
 wire \i44/n582 ;
 wire \i44/n59 ;
 wire \i44/n6 ;
 wire \i44/n60 ;
 wire \i44/n61 ;
 wire \i44/n62 ;
 wire \i44/n63 ;
 wire \i44/n64 ;
 wire \i44/n65 ;
 wire \i44/n66 ;
 wire \i44/n67 ;
 wire \i44/n68 ;
 wire \i44/n69 ;
 wire \i44/n7 ;
 wire \i44/n70 ;
 wire \i44/n71 ;
 wire \i44/n72 ;
 wire \i44/n73 ;
 wire \i44/n74 ;
 wire \i44/n75 ;
 wire \i44/n76 ;
 wire \i44/n77 ;
 wire \i44/n78 ;
 wire \i44/n79 ;
 wire \i44/n8 ;
 wire \i44/n80 ;
 wire \i44/n81 ;
 wire \i44/n82 ;
 wire \i44/n83 ;
 wire \i44/n84 ;
 wire \i44/n85 ;
 wire \i44/n86 ;
 wire \i44/n87 ;
 wire \i44/n88 ;
 wire \i44/n89 ;
 wire \i44/n9 ;
 wire \i44/n90 ;
 wire \i44/n91 ;
 wire \i44/n92 ;
 wire \i44/n93 ;
 wire \i44/n94 ;
 wire \i44/n95 ;
 wire \i44/n96 ;
 wire \i44/n97 ;
 wire \i44/n98 ;
 wire \i44/n99 ;
 wire \i45/n0 ;
 wire \i45/n1 ;
 wire \i45/n10 ;
 wire \i45/n100 ;
 wire \i45/n101 ;
 wire \i45/n102 ;
 wire \i45/n103 ;
 wire \i45/n104 ;
 wire \i45/n105 ;
 wire \i45/n106 ;
 wire \i45/n107 ;
 wire \i45/n108 ;
 wire \i45/n109 ;
 wire \i45/n11 ;
 wire \i45/n110 ;
 wire \i45/n111 ;
 wire \i45/n112 ;
 wire \i45/n113 ;
 wire \i45/n114 ;
 wire \i45/n115 ;
 wire \i45/n116 ;
 wire \i45/n117 ;
 wire \i45/n118 ;
 wire \i45/n119 ;
 wire \i45/n12 ;
 wire \i45/n120 ;
 wire \i45/n121 ;
 wire \i45/n122 ;
 wire \i45/n123 ;
 wire \i45/n124 ;
 wire \i45/n125 ;
 wire \i45/n126 ;
 wire \i45/n127 ;
 wire \i45/n128 ;
 wire \i45/n129 ;
 wire \i45/n13 ;
 wire \i45/n130 ;
 wire \i45/n131 ;
 wire \i45/n132 ;
 wire \i45/n133 ;
 wire \i45/n134 ;
 wire \i45/n135 ;
 wire \i45/n136 ;
 wire \i45/n137 ;
 wire \i45/n138 ;
 wire \i45/n139 ;
 wire \i45/n14 ;
 wire \i45/n140 ;
 wire \i45/n141 ;
 wire \i45/n142 ;
 wire \i45/n143 ;
 wire \i45/n144 ;
 wire \i45/n145 ;
 wire \i45/n146 ;
 wire \i45/n147 ;
 wire \i45/n148 ;
 wire \i45/n149 ;
 wire \i45/n15 ;
 wire \i45/n150 ;
 wire \i45/n151 ;
 wire \i45/n152 ;
 wire \i45/n153 ;
 wire \i45/n154 ;
 wire \i45/n155 ;
 wire \i45/n156 ;
 wire \i45/n157 ;
 wire \i45/n158 ;
 wire \i45/n159 ;
 wire \i45/n16 ;
 wire \i45/n160 ;
 wire \i45/n161 ;
 wire \i45/n162 ;
 wire \i45/n163 ;
 wire \i45/n164 ;
 wire \i45/n165 ;
 wire \i45/n166 ;
 wire \i45/n167 ;
 wire \i45/n168 ;
 wire \i45/n169 ;
 wire \i45/n17 ;
 wire \i45/n170 ;
 wire \i45/n171 ;
 wire \i45/n172 ;
 wire \i45/n173 ;
 wire \i45/n174 ;
 wire \i45/n175 ;
 wire \i45/n176 ;
 wire \i45/n177 ;
 wire \i45/n178 ;
 wire \i45/n179 ;
 wire \i45/n18 ;
 wire \i45/n180 ;
 wire \i45/n181 ;
 wire \i45/n182 ;
 wire \i45/n183 ;
 wire \i45/n184 ;
 wire \i45/n185 ;
 wire \i45/n186 ;
 wire \i45/n187 ;
 wire \i45/n188 ;
 wire \i45/n189 ;
 wire \i45/n19 ;
 wire \i45/n190 ;
 wire \i45/n191 ;
 wire \i45/n192 ;
 wire \i45/n193 ;
 wire \i45/n194 ;
 wire \i45/n195 ;
 wire \i45/n196 ;
 wire \i45/n197 ;
 wire \i45/n198 ;
 wire \i45/n199 ;
 wire \i45/n2 ;
 wire \i45/n20 ;
 wire \i45/n200 ;
 wire \i45/n201 ;
 wire \i45/n202 ;
 wire \i45/n203 ;
 wire \i45/n204 ;
 wire \i45/n205 ;
 wire \i45/n206 ;
 wire \i45/n207 ;
 wire \i45/n208 ;
 wire \i45/n209 ;
 wire \i45/n21 ;
 wire \i45/n210 ;
 wire \i45/n211 ;
 wire \i45/n212 ;
 wire \i45/n213 ;
 wire \i45/n214 ;
 wire \i45/n215 ;
 wire \i45/n216 ;
 wire \i45/n217 ;
 wire \i45/n218 ;
 wire \i45/n219 ;
 wire \i45/n22 ;
 wire \i45/n220 ;
 wire \i45/n221 ;
 wire \i45/n222 ;
 wire \i45/n223 ;
 wire \i45/n224 ;
 wire \i45/n225 ;
 wire \i45/n226 ;
 wire \i45/n227 ;
 wire \i45/n228 ;
 wire \i45/n229 ;
 wire \i45/n23 ;
 wire \i45/n230 ;
 wire \i45/n231 ;
 wire \i45/n232 ;
 wire \i45/n233 ;
 wire \i45/n234 ;
 wire \i45/n235 ;
 wire \i45/n236 ;
 wire \i45/n237 ;
 wire \i45/n238 ;
 wire \i45/n239 ;
 wire \i45/n24 ;
 wire \i45/n240 ;
 wire \i45/n241 ;
 wire \i45/n242 ;
 wire \i45/n243 ;
 wire \i45/n244 ;
 wire \i45/n245 ;
 wire \i45/n246 ;
 wire \i45/n247 ;
 wire \i45/n248 ;
 wire \i45/n249 ;
 wire \i45/n25 ;
 wire \i45/n250 ;
 wire \i45/n251 ;
 wire \i45/n252 ;
 wire \i45/n253 ;
 wire \i45/n254 ;
 wire \i45/n255 ;
 wire \i45/n256 ;
 wire \i45/n257 ;
 wire \i45/n258 ;
 wire \i45/n259 ;
 wire \i45/n26 ;
 wire \i45/n260 ;
 wire \i45/n261 ;
 wire \i45/n262 ;
 wire \i45/n263 ;
 wire \i45/n264 ;
 wire \i45/n265 ;
 wire \i45/n266 ;
 wire \i45/n267 ;
 wire \i45/n268 ;
 wire \i45/n269 ;
 wire \i45/n27 ;
 wire \i45/n270 ;
 wire \i45/n271 ;
 wire \i45/n272 ;
 wire \i45/n273 ;
 wire \i45/n274 ;
 wire \i45/n275 ;
 wire \i45/n276 ;
 wire \i45/n277 ;
 wire \i45/n278 ;
 wire \i45/n279 ;
 wire \i45/n28 ;
 wire \i45/n280 ;
 wire \i45/n281 ;
 wire \i45/n282 ;
 wire \i45/n283 ;
 wire \i45/n284 ;
 wire \i45/n285 ;
 wire \i45/n286 ;
 wire \i45/n287 ;
 wire \i45/n288 ;
 wire \i45/n289 ;
 wire \i45/n29 ;
 wire \i45/n290 ;
 wire \i45/n291 ;
 wire \i45/n292 ;
 wire \i45/n293 ;
 wire \i45/n294 ;
 wire \i45/n295 ;
 wire \i45/n296 ;
 wire \i45/n297 ;
 wire \i45/n298 ;
 wire \i45/n299 ;
 wire \i45/n3 ;
 wire \i45/n30 ;
 wire \i45/n300 ;
 wire \i45/n301 ;
 wire \i45/n302 ;
 wire \i45/n303 ;
 wire \i45/n304 ;
 wire \i45/n305 ;
 wire \i45/n306 ;
 wire \i45/n307 ;
 wire \i45/n308 ;
 wire \i45/n309 ;
 wire \i45/n31 ;
 wire \i45/n310 ;
 wire \i45/n311 ;
 wire \i45/n312 ;
 wire \i45/n313 ;
 wire \i45/n314 ;
 wire \i45/n315 ;
 wire \i45/n316 ;
 wire \i45/n317 ;
 wire \i45/n318 ;
 wire \i45/n319 ;
 wire \i45/n32 ;
 wire \i45/n320 ;
 wire \i45/n321 ;
 wire \i45/n322 ;
 wire \i45/n323 ;
 wire \i45/n324 ;
 wire \i45/n325 ;
 wire \i45/n326 ;
 wire \i45/n327 ;
 wire \i45/n328 ;
 wire \i45/n329 ;
 wire \i45/n33 ;
 wire \i45/n330 ;
 wire \i45/n331 ;
 wire \i45/n332 ;
 wire \i45/n333 ;
 wire \i45/n334 ;
 wire \i45/n335 ;
 wire \i45/n336 ;
 wire \i45/n337 ;
 wire \i45/n338 ;
 wire \i45/n339 ;
 wire \i45/n34 ;
 wire \i45/n340 ;
 wire \i45/n341 ;
 wire \i45/n342 ;
 wire \i45/n343 ;
 wire \i45/n344 ;
 wire \i45/n345 ;
 wire \i45/n346 ;
 wire \i45/n347 ;
 wire \i45/n348 ;
 wire \i45/n349 ;
 wire \i45/n35 ;
 wire \i45/n350 ;
 wire \i45/n351 ;
 wire \i45/n352 ;
 wire \i45/n353 ;
 wire \i45/n354 ;
 wire \i45/n355 ;
 wire \i45/n356 ;
 wire \i45/n357 ;
 wire \i45/n358 ;
 wire \i45/n359 ;
 wire \i45/n36 ;
 wire \i45/n360 ;
 wire \i45/n361 ;
 wire \i45/n362 ;
 wire \i45/n363 ;
 wire \i45/n364 ;
 wire \i45/n365 ;
 wire \i45/n366 ;
 wire \i45/n367 ;
 wire \i45/n368 ;
 wire \i45/n369 ;
 wire \i45/n37 ;
 wire \i45/n370 ;
 wire \i45/n371 ;
 wire \i45/n372 ;
 wire \i45/n373 ;
 wire \i45/n374 ;
 wire \i45/n375 ;
 wire \i45/n376 ;
 wire \i45/n377 ;
 wire \i45/n378 ;
 wire \i45/n379 ;
 wire \i45/n38 ;
 wire \i45/n380 ;
 wire \i45/n381 ;
 wire \i45/n382 ;
 wire \i45/n383 ;
 wire \i45/n384 ;
 wire \i45/n385 ;
 wire \i45/n386 ;
 wire \i45/n387 ;
 wire \i45/n388 ;
 wire \i45/n389 ;
 wire \i45/n39 ;
 wire \i45/n390 ;
 wire \i45/n391 ;
 wire \i45/n392 ;
 wire \i45/n393 ;
 wire \i45/n394 ;
 wire \i45/n395 ;
 wire \i45/n396 ;
 wire \i45/n397 ;
 wire \i45/n398 ;
 wire \i45/n399 ;
 wire \i45/n4 ;
 wire \i45/n40 ;
 wire \i45/n400 ;
 wire \i45/n401 ;
 wire \i45/n402 ;
 wire \i45/n403 ;
 wire \i45/n404 ;
 wire \i45/n405 ;
 wire \i45/n406 ;
 wire \i45/n407 ;
 wire \i45/n408 ;
 wire \i45/n409 ;
 wire \i45/n41 ;
 wire \i45/n410 ;
 wire \i45/n411 ;
 wire \i45/n412 ;
 wire \i45/n413 ;
 wire \i45/n414 ;
 wire \i45/n415 ;
 wire \i45/n416 ;
 wire \i45/n417 ;
 wire \i45/n418 ;
 wire \i45/n419 ;
 wire \i45/n42 ;
 wire \i45/n420 ;
 wire \i45/n421 ;
 wire \i45/n422 ;
 wire \i45/n423 ;
 wire \i45/n424 ;
 wire \i45/n425 ;
 wire \i45/n426 ;
 wire \i45/n427 ;
 wire \i45/n428 ;
 wire \i45/n429 ;
 wire \i45/n43 ;
 wire \i45/n430 ;
 wire \i45/n431 ;
 wire \i45/n432 ;
 wire \i45/n433 ;
 wire \i45/n434 ;
 wire \i45/n435 ;
 wire \i45/n436 ;
 wire \i45/n437 ;
 wire \i45/n438 ;
 wire \i45/n439 ;
 wire \i45/n44 ;
 wire \i45/n440 ;
 wire \i45/n441 ;
 wire \i45/n442 ;
 wire \i45/n443 ;
 wire \i45/n444 ;
 wire \i45/n445 ;
 wire \i45/n446 ;
 wire \i45/n447 ;
 wire \i45/n448 ;
 wire \i45/n449 ;
 wire \i45/n45 ;
 wire \i45/n450 ;
 wire \i45/n451 ;
 wire \i45/n452 ;
 wire \i45/n453 ;
 wire \i45/n454 ;
 wire \i45/n455 ;
 wire \i45/n456 ;
 wire \i45/n457 ;
 wire \i45/n458 ;
 wire \i45/n459 ;
 wire \i45/n46 ;
 wire \i45/n460 ;
 wire \i45/n461 ;
 wire \i45/n462 ;
 wire \i45/n463 ;
 wire \i45/n464 ;
 wire \i45/n465 ;
 wire \i45/n466 ;
 wire \i45/n467 ;
 wire \i45/n468 ;
 wire \i45/n469 ;
 wire \i45/n47 ;
 wire \i45/n470 ;
 wire \i45/n471 ;
 wire \i45/n472 ;
 wire \i45/n473 ;
 wire \i45/n474 ;
 wire \i45/n475 ;
 wire \i45/n476 ;
 wire \i45/n477 ;
 wire \i45/n478 ;
 wire \i45/n479 ;
 wire \i45/n48 ;
 wire \i45/n480 ;
 wire \i45/n481 ;
 wire \i45/n482 ;
 wire \i45/n483 ;
 wire \i45/n484 ;
 wire \i45/n485 ;
 wire \i45/n486 ;
 wire \i45/n487 ;
 wire \i45/n488 ;
 wire \i45/n489 ;
 wire \i45/n49 ;
 wire \i45/n490 ;
 wire \i45/n491 ;
 wire \i45/n492 ;
 wire \i45/n493 ;
 wire \i45/n494 ;
 wire \i45/n495 ;
 wire \i45/n496 ;
 wire \i45/n497 ;
 wire \i45/n498 ;
 wire \i45/n499 ;
 wire \i45/n5 ;
 wire \i45/n50 ;
 wire \i45/n500 ;
 wire \i45/n501 ;
 wire \i45/n502 ;
 wire \i45/n503 ;
 wire \i45/n504 ;
 wire \i45/n505 ;
 wire \i45/n506 ;
 wire \i45/n507 ;
 wire \i45/n508 ;
 wire \i45/n509 ;
 wire \i45/n51 ;
 wire \i45/n510 ;
 wire \i45/n511 ;
 wire \i45/n512 ;
 wire \i45/n513 ;
 wire \i45/n514 ;
 wire \i45/n515 ;
 wire \i45/n516 ;
 wire \i45/n517 ;
 wire \i45/n518 ;
 wire \i45/n519 ;
 wire \i45/n52 ;
 wire \i45/n520 ;
 wire \i45/n521 ;
 wire \i45/n522 ;
 wire \i45/n523 ;
 wire \i45/n524 ;
 wire \i45/n525 ;
 wire \i45/n526 ;
 wire \i45/n527 ;
 wire \i45/n528 ;
 wire \i45/n529 ;
 wire \i45/n53 ;
 wire \i45/n530 ;
 wire \i45/n531 ;
 wire \i45/n532 ;
 wire \i45/n533 ;
 wire \i45/n534 ;
 wire \i45/n535 ;
 wire \i45/n536 ;
 wire \i45/n537 ;
 wire \i45/n538 ;
 wire \i45/n539 ;
 wire \i45/n54 ;
 wire \i45/n540 ;
 wire \i45/n541 ;
 wire \i45/n542 ;
 wire \i45/n543 ;
 wire \i45/n544 ;
 wire \i45/n545 ;
 wire \i45/n546 ;
 wire \i45/n547 ;
 wire \i45/n548 ;
 wire \i45/n549 ;
 wire \i45/n55 ;
 wire \i45/n550 ;
 wire \i45/n551 ;
 wire \i45/n552 ;
 wire \i45/n553 ;
 wire \i45/n554 ;
 wire \i45/n555 ;
 wire \i45/n556 ;
 wire \i45/n557 ;
 wire \i45/n558 ;
 wire \i45/n559 ;
 wire \i45/n56 ;
 wire \i45/n560 ;
 wire \i45/n561 ;
 wire \i45/n562 ;
 wire \i45/n563 ;
 wire \i45/n564 ;
 wire \i45/n565 ;
 wire \i45/n566 ;
 wire \i45/n567 ;
 wire \i45/n568 ;
 wire \i45/n569 ;
 wire \i45/n57 ;
 wire \i45/n570 ;
 wire \i45/n571 ;
 wire \i45/n572 ;
 wire \i45/n573 ;
 wire \i45/n574 ;
 wire \i45/n575 ;
 wire \i45/n576 ;
 wire \i45/n577 ;
 wire \i45/n578 ;
 wire \i45/n579 ;
 wire \i45/n58 ;
 wire \i45/n580 ;
 wire \i45/n581 ;
 wire \i45/n582 ;
 wire \i45/n59 ;
 wire \i45/n6 ;
 wire \i45/n60 ;
 wire \i45/n61 ;
 wire \i45/n62 ;
 wire \i45/n63 ;
 wire \i45/n64 ;
 wire \i45/n65 ;
 wire \i45/n66 ;
 wire \i45/n67 ;
 wire \i45/n68 ;
 wire \i45/n69 ;
 wire \i45/n7 ;
 wire \i45/n70 ;
 wire \i45/n71 ;
 wire \i45/n72 ;
 wire \i45/n73 ;
 wire \i45/n74 ;
 wire \i45/n75 ;
 wire \i45/n76 ;
 wire \i45/n77 ;
 wire \i45/n78 ;
 wire \i45/n79 ;
 wire \i45/n8 ;
 wire \i45/n80 ;
 wire \i45/n81 ;
 wire \i45/n82 ;
 wire \i45/n83 ;
 wire \i45/n84 ;
 wire \i45/n85 ;
 wire \i45/n86 ;
 wire \i45/n87 ;
 wire \i45/n88 ;
 wire \i45/n89 ;
 wire \i45/n9 ;
 wire \i45/n90 ;
 wire \i45/n91 ;
 wire \i45/n92 ;
 wire \i45/n93 ;
 wire \i45/n94 ;
 wire \i45/n95 ;
 wire \i45/n96 ;
 wire \i45/n97 ;
 wire \i45/n98 ;
 wire \i45/n99 ;
 wire \i46/n0 ;
 wire \i46/n1 ;
 wire \i46/n10 ;
 wire \i46/n100 ;
 wire \i46/n101 ;
 wire \i46/n102 ;
 wire \i46/n103 ;
 wire \i46/n104 ;
 wire \i46/n105 ;
 wire \i46/n106 ;
 wire \i46/n107 ;
 wire \i46/n108 ;
 wire \i46/n109 ;
 wire \i46/n11 ;
 wire \i46/n110 ;
 wire \i46/n111 ;
 wire \i46/n112 ;
 wire \i46/n113 ;
 wire \i46/n114 ;
 wire \i46/n115 ;
 wire \i46/n116 ;
 wire \i46/n117 ;
 wire \i46/n118 ;
 wire \i46/n119 ;
 wire \i46/n12 ;
 wire \i46/n120 ;
 wire \i46/n121 ;
 wire \i46/n122 ;
 wire \i46/n123 ;
 wire \i46/n124 ;
 wire \i46/n125 ;
 wire \i46/n126 ;
 wire \i46/n127 ;
 wire \i46/n128 ;
 wire \i46/n129 ;
 wire \i46/n13 ;
 wire \i46/n130 ;
 wire \i46/n131 ;
 wire \i46/n132 ;
 wire \i46/n133 ;
 wire \i46/n134 ;
 wire \i46/n135 ;
 wire \i46/n136 ;
 wire \i46/n137 ;
 wire \i46/n138 ;
 wire \i46/n139 ;
 wire \i46/n14 ;
 wire \i46/n140 ;
 wire \i46/n141 ;
 wire \i46/n142 ;
 wire \i46/n143 ;
 wire \i46/n144 ;
 wire \i46/n145 ;
 wire \i46/n146 ;
 wire \i46/n147 ;
 wire \i46/n148 ;
 wire \i46/n149 ;
 wire \i46/n15 ;
 wire \i46/n150 ;
 wire \i46/n151 ;
 wire \i46/n152 ;
 wire \i46/n153 ;
 wire \i46/n154 ;
 wire \i46/n155 ;
 wire \i46/n156 ;
 wire \i46/n157 ;
 wire \i46/n158 ;
 wire \i46/n159 ;
 wire \i46/n16 ;
 wire \i46/n160 ;
 wire \i46/n161 ;
 wire \i46/n162 ;
 wire \i46/n163 ;
 wire \i46/n164 ;
 wire \i46/n165 ;
 wire \i46/n166 ;
 wire \i46/n167 ;
 wire \i46/n168 ;
 wire \i46/n169 ;
 wire \i46/n17 ;
 wire \i46/n170 ;
 wire \i46/n171 ;
 wire \i46/n172 ;
 wire \i46/n173 ;
 wire \i46/n174 ;
 wire \i46/n175 ;
 wire \i46/n176 ;
 wire \i46/n177 ;
 wire \i46/n178 ;
 wire \i46/n179 ;
 wire \i46/n18 ;
 wire \i46/n180 ;
 wire \i46/n181 ;
 wire \i46/n182 ;
 wire \i46/n183 ;
 wire \i46/n184 ;
 wire \i46/n185 ;
 wire \i46/n186 ;
 wire \i46/n187 ;
 wire \i46/n188 ;
 wire \i46/n189 ;
 wire \i46/n19 ;
 wire \i46/n190 ;
 wire \i46/n191 ;
 wire \i46/n192 ;
 wire \i46/n193 ;
 wire \i46/n194 ;
 wire \i46/n195 ;
 wire \i46/n196 ;
 wire \i46/n197 ;
 wire \i46/n198 ;
 wire \i46/n199 ;
 wire \i46/n2 ;
 wire \i46/n20 ;
 wire \i46/n200 ;
 wire \i46/n201 ;
 wire \i46/n202 ;
 wire \i46/n203 ;
 wire \i46/n204 ;
 wire \i46/n205 ;
 wire \i46/n206 ;
 wire \i46/n207 ;
 wire \i46/n208 ;
 wire \i46/n209 ;
 wire \i46/n21 ;
 wire \i46/n210 ;
 wire \i46/n211 ;
 wire \i46/n212 ;
 wire \i46/n213 ;
 wire \i46/n214 ;
 wire \i46/n215 ;
 wire \i46/n216 ;
 wire \i46/n217 ;
 wire \i46/n218 ;
 wire \i46/n219 ;
 wire \i46/n22 ;
 wire \i46/n220 ;
 wire \i46/n221 ;
 wire \i46/n222 ;
 wire \i46/n223 ;
 wire \i46/n224 ;
 wire \i46/n225 ;
 wire \i46/n226 ;
 wire \i46/n227 ;
 wire \i46/n228 ;
 wire \i46/n229 ;
 wire \i46/n23 ;
 wire \i46/n230 ;
 wire \i46/n231 ;
 wire \i46/n232 ;
 wire \i46/n233 ;
 wire \i46/n234 ;
 wire \i46/n235 ;
 wire \i46/n236 ;
 wire \i46/n237 ;
 wire \i46/n238 ;
 wire \i46/n239 ;
 wire \i46/n24 ;
 wire \i46/n240 ;
 wire \i46/n241 ;
 wire \i46/n242 ;
 wire \i46/n243 ;
 wire \i46/n244 ;
 wire \i46/n245 ;
 wire \i46/n246 ;
 wire \i46/n247 ;
 wire \i46/n248 ;
 wire \i46/n249 ;
 wire \i46/n25 ;
 wire \i46/n250 ;
 wire \i46/n251 ;
 wire \i46/n252 ;
 wire \i46/n253 ;
 wire \i46/n254 ;
 wire \i46/n255 ;
 wire \i46/n256 ;
 wire \i46/n257 ;
 wire \i46/n258 ;
 wire \i46/n259 ;
 wire \i46/n26 ;
 wire \i46/n260 ;
 wire \i46/n261 ;
 wire \i46/n262 ;
 wire \i46/n263 ;
 wire \i46/n264 ;
 wire \i46/n265 ;
 wire \i46/n266 ;
 wire \i46/n267 ;
 wire \i46/n268 ;
 wire \i46/n269 ;
 wire \i46/n27 ;
 wire \i46/n270 ;
 wire \i46/n271 ;
 wire \i46/n272 ;
 wire \i46/n273 ;
 wire \i46/n274 ;
 wire \i46/n275 ;
 wire \i46/n276 ;
 wire \i46/n277 ;
 wire \i46/n278 ;
 wire \i46/n279 ;
 wire \i46/n28 ;
 wire \i46/n280 ;
 wire \i46/n281 ;
 wire \i46/n282 ;
 wire \i46/n283 ;
 wire \i46/n284 ;
 wire \i46/n285 ;
 wire \i46/n286 ;
 wire \i46/n287 ;
 wire \i46/n288 ;
 wire \i46/n289 ;
 wire \i46/n29 ;
 wire \i46/n290 ;
 wire \i46/n291 ;
 wire \i46/n292 ;
 wire \i46/n293 ;
 wire \i46/n294 ;
 wire \i46/n295 ;
 wire \i46/n296 ;
 wire \i46/n297 ;
 wire \i46/n298 ;
 wire \i46/n299 ;
 wire \i46/n3 ;
 wire \i46/n30 ;
 wire \i46/n300 ;
 wire \i46/n301 ;
 wire \i46/n302 ;
 wire \i46/n303 ;
 wire \i46/n304 ;
 wire \i46/n305 ;
 wire \i46/n306 ;
 wire \i46/n307 ;
 wire \i46/n308 ;
 wire \i46/n309 ;
 wire \i46/n31 ;
 wire \i46/n310 ;
 wire \i46/n311 ;
 wire \i46/n312 ;
 wire \i46/n313 ;
 wire \i46/n314 ;
 wire \i46/n315 ;
 wire \i46/n316 ;
 wire \i46/n317 ;
 wire \i46/n318 ;
 wire \i46/n319 ;
 wire \i46/n32 ;
 wire \i46/n320 ;
 wire \i46/n321 ;
 wire \i46/n322 ;
 wire \i46/n323 ;
 wire \i46/n324 ;
 wire \i46/n325 ;
 wire \i46/n326 ;
 wire \i46/n327 ;
 wire \i46/n328 ;
 wire \i46/n329 ;
 wire \i46/n33 ;
 wire \i46/n330 ;
 wire \i46/n331 ;
 wire \i46/n332 ;
 wire \i46/n333 ;
 wire \i46/n334 ;
 wire \i46/n335 ;
 wire \i46/n336 ;
 wire \i46/n337 ;
 wire \i46/n338 ;
 wire \i46/n339 ;
 wire \i46/n34 ;
 wire \i46/n340 ;
 wire \i46/n341 ;
 wire \i46/n342 ;
 wire \i46/n343 ;
 wire \i46/n344 ;
 wire \i46/n345 ;
 wire \i46/n346 ;
 wire \i46/n347 ;
 wire \i46/n348 ;
 wire \i46/n349 ;
 wire \i46/n35 ;
 wire \i46/n350 ;
 wire \i46/n351 ;
 wire \i46/n352 ;
 wire \i46/n353 ;
 wire \i46/n354 ;
 wire \i46/n355 ;
 wire \i46/n356 ;
 wire \i46/n357 ;
 wire \i46/n358 ;
 wire \i46/n359 ;
 wire \i46/n36 ;
 wire \i46/n360 ;
 wire \i46/n361 ;
 wire \i46/n362 ;
 wire \i46/n363 ;
 wire \i46/n364 ;
 wire \i46/n365 ;
 wire \i46/n366 ;
 wire \i46/n367 ;
 wire \i46/n368 ;
 wire \i46/n369 ;
 wire \i46/n37 ;
 wire \i46/n370 ;
 wire \i46/n371 ;
 wire \i46/n372 ;
 wire \i46/n373 ;
 wire \i46/n374 ;
 wire \i46/n375 ;
 wire \i46/n376 ;
 wire \i46/n377 ;
 wire \i46/n378 ;
 wire \i46/n379 ;
 wire \i46/n38 ;
 wire \i46/n380 ;
 wire \i46/n381 ;
 wire \i46/n382 ;
 wire \i46/n383 ;
 wire \i46/n384 ;
 wire \i46/n385 ;
 wire \i46/n386 ;
 wire \i46/n387 ;
 wire \i46/n388 ;
 wire \i46/n389 ;
 wire \i46/n39 ;
 wire \i46/n390 ;
 wire \i46/n391 ;
 wire \i46/n392 ;
 wire \i46/n393 ;
 wire \i46/n394 ;
 wire \i46/n395 ;
 wire \i46/n396 ;
 wire \i46/n397 ;
 wire \i46/n398 ;
 wire \i46/n399 ;
 wire \i46/n4 ;
 wire \i46/n40 ;
 wire \i46/n400 ;
 wire \i46/n401 ;
 wire \i46/n402 ;
 wire \i46/n403 ;
 wire \i46/n404 ;
 wire \i46/n405 ;
 wire \i46/n406 ;
 wire \i46/n407 ;
 wire \i46/n408 ;
 wire \i46/n409 ;
 wire \i46/n41 ;
 wire \i46/n410 ;
 wire \i46/n411 ;
 wire \i46/n412 ;
 wire \i46/n413 ;
 wire \i46/n414 ;
 wire \i46/n415 ;
 wire \i46/n416 ;
 wire \i46/n417 ;
 wire \i46/n418 ;
 wire \i46/n419 ;
 wire \i46/n42 ;
 wire \i46/n420 ;
 wire \i46/n421 ;
 wire \i46/n422 ;
 wire \i46/n423 ;
 wire \i46/n424 ;
 wire \i46/n425 ;
 wire \i46/n426 ;
 wire \i46/n427 ;
 wire \i46/n428 ;
 wire \i46/n429 ;
 wire \i46/n43 ;
 wire \i46/n430 ;
 wire \i46/n431 ;
 wire \i46/n432 ;
 wire \i46/n433 ;
 wire \i46/n434 ;
 wire \i46/n435 ;
 wire \i46/n436 ;
 wire \i46/n437 ;
 wire \i46/n438 ;
 wire \i46/n439 ;
 wire \i46/n44 ;
 wire \i46/n440 ;
 wire \i46/n441 ;
 wire \i46/n442 ;
 wire \i46/n443 ;
 wire \i46/n444 ;
 wire \i46/n445 ;
 wire \i46/n446 ;
 wire \i46/n447 ;
 wire \i46/n448 ;
 wire \i46/n449 ;
 wire \i46/n45 ;
 wire \i46/n450 ;
 wire \i46/n451 ;
 wire \i46/n452 ;
 wire \i46/n453 ;
 wire \i46/n454 ;
 wire \i46/n455 ;
 wire \i46/n456 ;
 wire \i46/n457 ;
 wire \i46/n458 ;
 wire \i46/n459 ;
 wire \i46/n46 ;
 wire \i46/n460 ;
 wire \i46/n461 ;
 wire \i46/n462 ;
 wire \i46/n463 ;
 wire \i46/n464 ;
 wire \i46/n465 ;
 wire \i46/n466 ;
 wire \i46/n467 ;
 wire \i46/n468 ;
 wire \i46/n469 ;
 wire \i46/n47 ;
 wire \i46/n470 ;
 wire \i46/n471 ;
 wire \i46/n472 ;
 wire \i46/n473 ;
 wire \i46/n474 ;
 wire \i46/n475 ;
 wire \i46/n476 ;
 wire \i46/n477 ;
 wire \i46/n478 ;
 wire \i46/n479 ;
 wire \i46/n48 ;
 wire \i46/n480 ;
 wire \i46/n481 ;
 wire \i46/n482 ;
 wire \i46/n483 ;
 wire \i46/n484 ;
 wire \i46/n485 ;
 wire \i46/n486 ;
 wire \i46/n487 ;
 wire \i46/n488 ;
 wire \i46/n489 ;
 wire \i46/n49 ;
 wire \i46/n490 ;
 wire \i46/n491 ;
 wire \i46/n492 ;
 wire \i46/n493 ;
 wire \i46/n494 ;
 wire \i46/n495 ;
 wire \i46/n496 ;
 wire \i46/n497 ;
 wire \i46/n498 ;
 wire \i46/n499 ;
 wire \i46/n5 ;
 wire \i46/n50 ;
 wire \i46/n500 ;
 wire \i46/n501 ;
 wire \i46/n502 ;
 wire \i46/n503 ;
 wire \i46/n504 ;
 wire \i46/n505 ;
 wire \i46/n506 ;
 wire \i46/n507 ;
 wire \i46/n508 ;
 wire \i46/n509 ;
 wire \i46/n51 ;
 wire \i46/n510 ;
 wire \i46/n511 ;
 wire \i46/n512 ;
 wire \i46/n513 ;
 wire \i46/n514 ;
 wire \i46/n515 ;
 wire \i46/n516 ;
 wire \i46/n517 ;
 wire \i46/n518 ;
 wire \i46/n519 ;
 wire \i46/n52 ;
 wire \i46/n520 ;
 wire \i46/n521 ;
 wire \i46/n522 ;
 wire \i46/n523 ;
 wire \i46/n524 ;
 wire \i46/n525 ;
 wire \i46/n526 ;
 wire \i46/n527 ;
 wire \i46/n528 ;
 wire \i46/n529 ;
 wire \i46/n53 ;
 wire \i46/n530 ;
 wire \i46/n531 ;
 wire \i46/n532 ;
 wire \i46/n533 ;
 wire \i46/n534 ;
 wire \i46/n535 ;
 wire \i46/n536 ;
 wire \i46/n537 ;
 wire \i46/n538 ;
 wire \i46/n539 ;
 wire \i46/n54 ;
 wire \i46/n540 ;
 wire \i46/n541 ;
 wire \i46/n542 ;
 wire \i46/n543 ;
 wire \i46/n544 ;
 wire \i46/n545 ;
 wire \i46/n546 ;
 wire \i46/n547 ;
 wire \i46/n548 ;
 wire \i46/n549 ;
 wire \i46/n55 ;
 wire \i46/n550 ;
 wire \i46/n551 ;
 wire \i46/n552 ;
 wire \i46/n553 ;
 wire \i46/n554 ;
 wire \i46/n555 ;
 wire \i46/n556 ;
 wire \i46/n557 ;
 wire \i46/n558 ;
 wire \i46/n559 ;
 wire \i46/n56 ;
 wire \i46/n560 ;
 wire \i46/n561 ;
 wire \i46/n562 ;
 wire \i46/n563 ;
 wire \i46/n564 ;
 wire \i46/n565 ;
 wire \i46/n566 ;
 wire \i46/n567 ;
 wire \i46/n568 ;
 wire \i46/n569 ;
 wire \i46/n57 ;
 wire \i46/n570 ;
 wire \i46/n571 ;
 wire \i46/n572 ;
 wire \i46/n573 ;
 wire \i46/n574 ;
 wire \i46/n575 ;
 wire \i46/n576 ;
 wire \i46/n577 ;
 wire \i46/n578 ;
 wire \i46/n579 ;
 wire \i46/n58 ;
 wire \i46/n580 ;
 wire \i46/n581 ;
 wire \i46/n59 ;
 wire \i46/n6 ;
 wire \i46/n60 ;
 wire \i46/n61 ;
 wire \i46/n62 ;
 wire \i46/n63 ;
 wire \i46/n64 ;
 wire \i46/n65 ;
 wire \i46/n66 ;
 wire \i46/n67 ;
 wire \i46/n68 ;
 wire \i46/n69 ;
 wire \i46/n7 ;
 wire \i46/n70 ;
 wire \i46/n71 ;
 wire \i46/n72 ;
 wire \i46/n73 ;
 wire \i46/n74 ;
 wire \i46/n75 ;
 wire \i46/n76 ;
 wire \i46/n77 ;
 wire \i46/n78 ;
 wire \i46/n79 ;
 wire \i46/n8 ;
 wire \i46/n80 ;
 wire \i46/n81 ;
 wire \i46/n82 ;
 wire \i46/n83 ;
 wire \i46/n84 ;
 wire \i46/n85 ;
 wire \i46/n86 ;
 wire \i46/n87 ;
 wire \i46/n88 ;
 wire \i46/n89 ;
 wire \i46/n9 ;
 wire \i46/n90 ;
 wire \i46/n91 ;
 wire \i46/n92 ;
 wire \i46/n93 ;
 wire \i46/n94 ;
 wire \i46/n95 ;
 wire \i46/n96 ;
 wire \i46/n97 ;
 wire \i46/n98 ;
 wire \i46/n99 ;
 wire \i47/n0 ;
 wire \i47/n1 ;
 wire \i47/n10 ;
 wire \i47/n100 ;
 wire \i47/n101 ;
 wire \i47/n102 ;
 wire \i47/n103 ;
 wire \i47/n104 ;
 wire \i47/n105 ;
 wire \i47/n106 ;
 wire \i47/n107 ;
 wire \i47/n108 ;
 wire \i47/n109 ;
 wire \i47/n11 ;
 wire \i47/n110 ;
 wire \i47/n111 ;
 wire \i47/n112 ;
 wire \i47/n113 ;
 wire \i47/n114 ;
 wire \i47/n115 ;
 wire \i47/n116 ;
 wire \i47/n117 ;
 wire \i47/n118 ;
 wire \i47/n119 ;
 wire \i47/n12 ;
 wire \i47/n120 ;
 wire \i47/n121 ;
 wire \i47/n122 ;
 wire \i47/n123 ;
 wire \i47/n124 ;
 wire \i47/n125 ;
 wire \i47/n126 ;
 wire \i47/n127 ;
 wire \i47/n128 ;
 wire \i47/n129 ;
 wire \i47/n13 ;
 wire \i47/n130 ;
 wire \i47/n131 ;
 wire \i47/n132 ;
 wire \i47/n133 ;
 wire \i47/n134 ;
 wire \i47/n135 ;
 wire \i47/n136 ;
 wire \i47/n137 ;
 wire \i47/n138 ;
 wire \i47/n139 ;
 wire \i47/n14 ;
 wire \i47/n140 ;
 wire \i47/n141 ;
 wire \i47/n142 ;
 wire \i47/n143 ;
 wire \i47/n144 ;
 wire \i47/n145 ;
 wire \i47/n146 ;
 wire \i47/n147 ;
 wire \i47/n148 ;
 wire \i47/n149 ;
 wire \i47/n15 ;
 wire \i47/n150 ;
 wire \i47/n151 ;
 wire \i47/n152 ;
 wire \i47/n153 ;
 wire \i47/n154 ;
 wire \i47/n155 ;
 wire \i47/n156 ;
 wire \i47/n157 ;
 wire \i47/n158 ;
 wire \i47/n159 ;
 wire \i47/n16 ;
 wire \i47/n160 ;
 wire \i47/n161 ;
 wire \i47/n162 ;
 wire \i47/n163 ;
 wire \i47/n164 ;
 wire \i47/n165 ;
 wire \i47/n166 ;
 wire \i47/n167 ;
 wire \i47/n168 ;
 wire \i47/n169 ;
 wire \i47/n17 ;
 wire \i47/n170 ;
 wire \i47/n171 ;
 wire \i47/n172 ;
 wire \i47/n173 ;
 wire \i47/n174 ;
 wire \i47/n175 ;
 wire \i47/n176 ;
 wire \i47/n177 ;
 wire \i47/n178 ;
 wire \i47/n179 ;
 wire \i47/n18 ;
 wire \i47/n180 ;
 wire \i47/n181 ;
 wire \i47/n182 ;
 wire \i47/n183 ;
 wire \i47/n184 ;
 wire \i47/n185 ;
 wire \i47/n186 ;
 wire \i47/n187 ;
 wire \i47/n188 ;
 wire \i47/n189 ;
 wire \i47/n19 ;
 wire \i47/n190 ;
 wire \i47/n191 ;
 wire \i47/n192 ;
 wire \i47/n193 ;
 wire \i47/n194 ;
 wire \i47/n195 ;
 wire \i47/n196 ;
 wire \i47/n197 ;
 wire \i47/n198 ;
 wire \i47/n199 ;
 wire \i47/n2 ;
 wire \i47/n20 ;
 wire \i47/n200 ;
 wire \i47/n201 ;
 wire \i47/n202 ;
 wire \i47/n203 ;
 wire \i47/n204 ;
 wire \i47/n205 ;
 wire \i47/n206 ;
 wire \i47/n207 ;
 wire \i47/n208 ;
 wire \i47/n209 ;
 wire \i47/n21 ;
 wire \i47/n210 ;
 wire \i47/n211 ;
 wire \i47/n212 ;
 wire \i47/n213 ;
 wire \i47/n214 ;
 wire \i47/n215 ;
 wire \i47/n216 ;
 wire \i47/n217 ;
 wire \i47/n218 ;
 wire \i47/n219 ;
 wire \i47/n22 ;
 wire \i47/n220 ;
 wire \i47/n221 ;
 wire \i47/n222 ;
 wire \i47/n223 ;
 wire \i47/n224 ;
 wire \i47/n225 ;
 wire \i47/n226 ;
 wire \i47/n227 ;
 wire \i47/n228 ;
 wire \i47/n229 ;
 wire \i47/n23 ;
 wire \i47/n230 ;
 wire \i47/n231 ;
 wire \i47/n232 ;
 wire \i47/n233 ;
 wire \i47/n234 ;
 wire \i47/n235 ;
 wire \i47/n236 ;
 wire \i47/n237 ;
 wire \i47/n238 ;
 wire \i47/n239 ;
 wire \i47/n24 ;
 wire \i47/n240 ;
 wire \i47/n241 ;
 wire \i47/n242 ;
 wire \i47/n243 ;
 wire \i47/n244 ;
 wire \i47/n245 ;
 wire \i47/n246 ;
 wire \i47/n247 ;
 wire \i47/n248 ;
 wire \i47/n249 ;
 wire \i47/n25 ;
 wire \i47/n250 ;
 wire \i47/n251 ;
 wire \i47/n252 ;
 wire \i47/n253 ;
 wire \i47/n254 ;
 wire \i47/n255 ;
 wire \i47/n256 ;
 wire \i47/n257 ;
 wire \i47/n258 ;
 wire \i47/n259 ;
 wire \i47/n26 ;
 wire \i47/n260 ;
 wire \i47/n261 ;
 wire \i47/n262 ;
 wire \i47/n263 ;
 wire \i47/n264 ;
 wire \i47/n265 ;
 wire \i47/n266 ;
 wire \i47/n267 ;
 wire \i47/n268 ;
 wire \i47/n269 ;
 wire \i47/n27 ;
 wire \i47/n270 ;
 wire \i47/n271 ;
 wire \i47/n272 ;
 wire \i47/n273 ;
 wire \i47/n274 ;
 wire \i47/n275 ;
 wire \i47/n276 ;
 wire \i47/n277 ;
 wire \i47/n278 ;
 wire \i47/n279 ;
 wire \i47/n28 ;
 wire \i47/n280 ;
 wire \i47/n281 ;
 wire \i47/n282 ;
 wire \i47/n283 ;
 wire \i47/n284 ;
 wire \i47/n285 ;
 wire \i47/n286 ;
 wire \i47/n287 ;
 wire \i47/n288 ;
 wire \i47/n289 ;
 wire \i47/n29 ;
 wire \i47/n290 ;
 wire \i47/n291 ;
 wire \i47/n292 ;
 wire \i47/n293 ;
 wire \i47/n294 ;
 wire \i47/n295 ;
 wire \i47/n296 ;
 wire \i47/n297 ;
 wire \i47/n298 ;
 wire \i47/n299 ;
 wire \i47/n3 ;
 wire \i47/n30 ;
 wire \i47/n300 ;
 wire \i47/n301 ;
 wire \i47/n302 ;
 wire \i47/n303 ;
 wire \i47/n304 ;
 wire \i47/n305 ;
 wire \i47/n306 ;
 wire \i47/n307 ;
 wire \i47/n308 ;
 wire \i47/n309 ;
 wire \i47/n31 ;
 wire \i47/n310 ;
 wire \i47/n311 ;
 wire \i47/n312 ;
 wire \i47/n313 ;
 wire \i47/n314 ;
 wire \i47/n315 ;
 wire \i47/n316 ;
 wire \i47/n317 ;
 wire \i47/n318 ;
 wire \i47/n319 ;
 wire \i47/n32 ;
 wire \i47/n320 ;
 wire \i47/n321 ;
 wire \i47/n322 ;
 wire \i47/n323 ;
 wire \i47/n324 ;
 wire \i47/n325 ;
 wire \i47/n326 ;
 wire \i47/n327 ;
 wire \i47/n328 ;
 wire \i47/n329 ;
 wire \i47/n33 ;
 wire \i47/n330 ;
 wire \i47/n331 ;
 wire \i47/n332 ;
 wire \i47/n333 ;
 wire \i47/n334 ;
 wire \i47/n335 ;
 wire \i47/n336 ;
 wire \i47/n337 ;
 wire \i47/n338 ;
 wire \i47/n339 ;
 wire \i47/n34 ;
 wire \i47/n340 ;
 wire \i47/n341 ;
 wire \i47/n342 ;
 wire \i47/n343 ;
 wire \i47/n344 ;
 wire \i47/n345 ;
 wire \i47/n346 ;
 wire \i47/n347 ;
 wire \i47/n348 ;
 wire \i47/n349 ;
 wire \i47/n35 ;
 wire \i47/n350 ;
 wire \i47/n351 ;
 wire \i47/n352 ;
 wire \i47/n353 ;
 wire \i47/n354 ;
 wire \i47/n355 ;
 wire \i47/n356 ;
 wire \i47/n357 ;
 wire \i47/n358 ;
 wire \i47/n359 ;
 wire \i47/n36 ;
 wire \i47/n360 ;
 wire \i47/n361 ;
 wire \i47/n362 ;
 wire \i47/n363 ;
 wire \i47/n364 ;
 wire \i47/n365 ;
 wire \i47/n366 ;
 wire \i47/n367 ;
 wire \i47/n368 ;
 wire \i47/n369 ;
 wire \i47/n37 ;
 wire \i47/n370 ;
 wire \i47/n371 ;
 wire \i47/n372 ;
 wire \i47/n373 ;
 wire \i47/n374 ;
 wire \i47/n375 ;
 wire \i47/n376 ;
 wire \i47/n377 ;
 wire \i47/n378 ;
 wire \i47/n379 ;
 wire \i47/n38 ;
 wire \i47/n380 ;
 wire \i47/n381 ;
 wire \i47/n382 ;
 wire \i47/n383 ;
 wire \i47/n384 ;
 wire \i47/n385 ;
 wire \i47/n386 ;
 wire \i47/n387 ;
 wire \i47/n388 ;
 wire \i47/n389 ;
 wire \i47/n39 ;
 wire \i47/n390 ;
 wire \i47/n391 ;
 wire \i47/n392 ;
 wire \i47/n393 ;
 wire \i47/n394 ;
 wire \i47/n395 ;
 wire \i47/n396 ;
 wire \i47/n397 ;
 wire \i47/n398 ;
 wire \i47/n399 ;
 wire \i47/n4 ;
 wire \i47/n40 ;
 wire \i47/n400 ;
 wire \i47/n401 ;
 wire \i47/n402 ;
 wire \i47/n403 ;
 wire \i47/n404 ;
 wire \i47/n405 ;
 wire \i47/n406 ;
 wire \i47/n407 ;
 wire \i47/n408 ;
 wire \i47/n409 ;
 wire \i47/n41 ;
 wire \i47/n410 ;
 wire \i47/n411 ;
 wire \i47/n412 ;
 wire \i47/n413 ;
 wire \i47/n414 ;
 wire \i47/n415 ;
 wire \i47/n416 ;
 wire \i47/n417 ;
 wire \i47/n418 ;
 wire \i47/n419 ;
 wire \i47/n42 ;
 wire \i47/n420 ;
 wire \i47/n421 ;
 wire \i47/n422 ;
 wire \i47/n423 ;
 wire \i47/n424 ;
 wire \i47/n425 ;
 wire \i47/n426 ;
 wire \i47/n427 ;
 wire \i47/n428 ;
 wire \i47/n429 ;
 wire \i47/n43 ;
 wire \i47/n430 ;
 wire \i47/n431 ;
 wire \i47/n432 ;
 wire \i47/n433 ;
 wire \i47/n434 ;
 wire \i47/n435 ;
 wire \i47/n436 ;
 wire \i47/n437 ;
 wire \i47/n438 ;
 wire \i47/n439 ;
 wire \i47/n44 ;
 wire \i47/n440 ;
 wire \i47/n441 ;
 wire \i47/n442 ;
 wire \i47/n443 ;
 wire \i47/n444 ;
 wire \i47/n445 ;
 wire \i47/n446 ;
 wire \i47/n447 ;
 wire \i47/n448 ;
 wire \i47/n449 ;
 wire \i47/n45 ;
 wire \i47/n450 ;
 wire \i47/n451 ;
 wire \i47/n452 ;
 wire \i47/n453 ;
 wire \i47/n454 ;
 wire \i47/n455 ;
 wire \i47/n456 ;
 wire \i47/n457 ;
 wire \i47/n458 ;
 wire \i47/n459 ;
 wire \i47/n46 ;
 wire \i47/n460 ;
 wire \i47/n461 ;
 wire \i47/n462 ;
 wire \i47/n463 ;
 wire \i47/n464 ;
 wire \i47/n465 ;
 wire \i47/n466 ;
 wire \i47/n467 ;
 wire \i47/n468 ;
 wire \i47/n469 ;
 wire \i47/n47 ;
 wire \i47/n470 ;
 wire \i47/n471 ;
 wire \i47/n472 ;
 wire \i47/n473 ;
 wire \i47/n474 ;
 wire \i47/n475 ;
 wire \i47/n476 ;
 wire \i47/n477 ;
 wire \i47/n478 ;
 wire \i47/n479 ;
 wire \i47/n48 ;
 wire \i47/n480 ;
 wire \i47/n481 ;
 wire \i47/n482 ;
 wire \i47/n483 ;
 wire \i47/n484 ;
 wire \i47/n485 ;
 wire \i47/n486 ;
 wire \i47/n487 ;
 wire \i47/n488 ;
 wire \i47/n489 ;
 wire \i47/n49 ;
 wire \i47/n490 ;
 wire \i47/n491 ;
 wire \i47/n492 ;
 wire \i47/n493 ;
 wire \i47/n494 ;
 wire \i47/n495 ;
 wire \i47/n496 ;
 wire \i47/n497 ;
 wire \i47/n498 ;
 wire \i47/n499 ;
 wire \i47/n5 ;
 wire \i47/n50 ;
 wire \i47/n500 ;
 wire \i47/n501 ;
 wire \i47/n502 ;
 wire \i47/n503 ;
 wire \i47/n504 ;
 wire \i47/n505 ;
 wire \i47/n506 ;
 wire \i47/n507 ;
 wire \i47/n508 ;
 wire \i47/n509 ;
 wire \i47/n51 ;
 wire \i47/n510 ;
 wire \i47/n511 ;
 wire \i47/n512 ;
 wire \i47/n513 ;
 wire \i47/n514 ;
 wire \i47/n515 ;
 wire \i47/n516 ;
 wire \i47/n517 ;
 wire \i47/n518 ;
 wire \i47/n519 ;
 wire \i47/n52 ;
 wire \i47/n520 ;
 wire \i47/n521 ;
 wire \i47/n522 ;
 wire \i47/n523 ;
 wire \i47/n524 ;
 wire \i47/n525 ;
 wire \i47/n526 ;
 wire \i47/n527 ;
 wire \i47/n528 ;
 wire \i47/n529 ;
 wire \i47/n53 ;
 wire \i47/n530 ;
 wire \i47/n531 ;
 wire \i47/n532 ;
 wire \i47/n533 ;
 wire \i47/n534 ;
 wire \i47/n535 ;
 wire \i47/n536 ;
 wire \i47/n537 ;
 wire \i47/n538 ;
 wire \i47/n539 ;
 wire \i47/n54 ;
 wire \i47/n540 ;
 wire \i47/n541 ;
 wire \i47/n542 ;
 wire \i47/n543 ;
 wire \i47/n544 ;
 wire \i47/n545 ;
 wire \i47/n546 ;
 wire \i47/n547 ;
 wire \i47/n548 ;
 wire \i47/n549 ;
 wire \i47/n55 ;
 wire \i47/n550 ;
 wire \i47/n551 ;
 wire \i47/n552 ;
 wire \i47/n553 ;
 wire \i47/n554 ;
 wire \i47/n555 ;
 wire \i47/n556 ;
 wire \i47/n557 ;
 wire \i47/n558 ;
 wire \i47/n559 ;
 wire \i47/n56 ;
 wire \i47/n560 ;
 wire \i47/n561 ;
 wire \i47/n562 ;
 wire \i47/n563 ;
 wire \i47/n564 ;
 wire \i47/n565 ;
 wire \i47/n566 ;
 wire \i47/n567 ;
 wire \i47/n568 ;
 wire \i47/n569 ;
 wire \i47/n57 ;
 wire \i47/n570 ;
 wire \i47/n571 ;
 wire \i47/n572 ;
 wire \i47/n573 ;
 wire \i47/n574 ;
 wire \i47/n575 ;
 wire \i47/n576 ;
 wire \i47/n577 ;
 wire \i47/n578 ;
 wire \i47/n579 ;
 wire \i47/n58 ;
 wire \i47/n59 ;
 wire \i47/n6 ;
 wire \i47/n60 ;
 wire \i47/n61 ;
 wire \i47/n62 ;
 wire \i47/n63 ;
 wire \i47/n64 ;
 wire \i47/n65 ;
 wire \i47/n66 ;
 wire \i47/n67 ;
 wire \i47/n68 ;
 wire \i47/n69 ;
 wire \i47/n7 ;
 wire \i47/n70 ;
 wire \i47/n71 ;
 wire \i47/n72 ;
 wire \i47/n73 ;
 wire \i47/n74 ;
 wire \i47/n75 ;
 wire \i47/n76 ;
 wire \i47/n77 ;
 wire \i47/n78 ;
 wire \i47/n79 ;
 wire \i47/n8 ;
 wire \i47/n80 ;
 wire \i47/n81 ;
 wire \i47/n82 ;
 wire \i47/n83 ;
 wire \i47/n84 ;
 wire \i47/n85 ;
 wire \i47/n86 ;
 wire \i47/n87 ;
 wire \i47/n88 ;
 wire \i47/n89 ;
 wire \i47/n9 ;
 wire \i47/n90 ;
 wire \i47/n91 ;
 wire \i47/n92 ;
 wire \i47/n93 ;
 wire \i47/n94 ;
 wire \i47/n95 ;
 wire \i47/n96 ;
 wire \i47/n97 ;
 wire \i47/n98 ;
 wire \i47/n99 ;
 wire \i48/n0 ;
 wire \i48/n1 ;
 wire \i48/n10 ;
 wire \i48/n100 ;
 wire \i48/n101 ;
 wire \i48/n102 ;
 wire \i48/n103 ;
 wire \i48/n104 ;
 wire \i48/n105 ;
 wire \i48/n106 ;
 wire \i48/n107 ;
 wire \i48/n108 ;
 wire \i48/n109 ;
 wire \i48/n11 ;
 wire \i48/n110 ;
 wire \i48/n111 ;
 wire \i48/n112 ;
 wire \i48/n113 ;
 wire \i48/n114 ;
 wire \i48/n115 ;
 wire \i48/n116 ;
 wire \i48/n117 ;
 wire \i48/n118 ;
 wire \i48/n119 ;
 wire \i48/n12 ;
 wire \i48/n120 ;
 wire \i48/n121 ;
 wire \i48/n122 ;
 wire \i48/n123 ;
 wire \i48/n124 ;
 wire \i48/n125 ;
 wire \i48/n126 ;
 wire \i48/n127 ;
 wire \i48/n128 ;
 wire \i48/n129 ;
 wire \i48/n13 ;
 wire \i48/n130 ;
 wire \i48/n131 ;
 wire \i48/n132 ;
 wire \i48/n133 ;
 wire \i48/n134 ;
 wire \i48/n135 ;
 wire \i48/n136 ;
 wire \i48/n137 ;
 wire \i48/n138 ;
 wire \i48/n139 ;
 wire \i48/n14 ;
 wire \i48/n140 ;
 wire \i48/n141 ;
 wire \i48/n142 ;
 wire \i48/n143 ;
 wire \i48/n144 ;
 wire \i48/n145 ;
 wire \i48/n146 ;
 wire \i48/n147 ;
 wire \i48/n148 ;
 wire \i48/n149 ;
 wire \i48/n15 ;
 wire \i48/n150 ;
 wire \i48/n151 ;
 wire \i48/n152 ;
 wire \i48/n153 ;
 wire \i48/n154 ;
 wire \i48/n155 ;
 wire \i48/n156 ;
 wire \i48/n157 ;
 wire \i48/n158 ;
 wire \i48/n159 ;
 wire \i48/n16 ;
 wire \i48/n160 ;
 wire \i48/n161 ;
 wire \i48/n162 ;
 wire \i48/n163 ;
 wire \i48/n164 ;
 wire \i48/n165 ;
 wire \i48/n166 ;
 wire \i48/n167 ;
 wire \i48/n168 ;
 wire \i48/n169 ;
 wire \i48/n17 ;
 wire \i48/n170 ;
 wire \i48/n171 ;
 wire \i48/n172 ;
 wire \i48/n173 ;
 wire \i48/n174 ;
 wire \i48/n175 ;
 wire \i48/n176 ;
 wire \i48/n177 ;
 wire \i48/n178 ;
 wire \i48/n179 ;
 wire \i48/n18 ;
 wire \i48/n180 ;
 wire \i48/n181 ;
 wire \i48/n182 ;
 wire \i48/n183 ;
 wire \i48/n184 ;
 wire \i48/n185 ;
 wire \i48/n186 ;
 wire \i48/n187 ;
 wire \i48/n188 ;
 wire \i48/n189 ;
 wire \i48/n19 ;
 wire \i48/n190 ;
 wire \i48/n191 ;
 wire \i48/n192 ;
 wire \i48/n193 ;
 wire \i48/n194 ;
 wire \i48/n195 ;
 wire \i48/n196 ;
 wire \i48/n197 ;
 wire \i48/n198 ;
 wire \i48/n199 ;
 wire \i48/n2 ;
 wire \i48/n20 ;
 wire \i48/n200 ;
 wire \i48/n201 ;
 wire \i48/n202 ;
 wire \i48/n203 ;
 wire \i48/n204 ;
 wire \i48/n205 ;
 wire \i48/n206 ;
 wire \i48/n207 ;
 wire \i48/n208 ;
 wire \i48/n209 ;
 wire \i48/n21 ;
 wire \i48/n210 ;
 wire \i48/n211 ;
 wire \i48/n212 ;
 wire \i48/n213 ;
 wire \i48/n214 ;
 wire \i48/n215 ;
 wire \i48/n216 ;
 wire \i48/n217 ;
 wire \i48/n218 ;
 wire \i48/n219 ;
 wire \i48/n22 ;
 wire \i48/n220 ;
 wire \i48/n221 ;
 wire \i48/n222 ;
 wire \i48/n223 ;
 wire \i48/n224 ;
 wire \i48/n225 ;
 wire \i48/n226 ;
 wire \i48/n227 ;
 wire \i48/n228 ;
 wire \i48/n229 ;
 wire \i48/n23 ;
 wire \i48/n230 ;
 wire \i48/n231 ;
 wire \i48/n232 ;
 wire \i48/n233 ;
 wire \i48/n234 ;
 wire \i48/n235 ;
 wire \i48/n236 ;
 wire \i48/n237 ;
 wire \i48/n238 ;
 wire \i48/n239 ;
 wire \i48/n24 ;
 wire \i48/n240 ;
 wire \i48/n241 ;
 wire \i48/n242 ;
 wire \i48/n243 ;
 wire \i48/n244 ;
 wire \i48/n245 ;
 wire \i48/n246 ;
 wire \i48/n247 ;
 wire \i48/n248 ;
 wire \i48/n249 ;
 wire \i48/n25 ;
 wire \i48/n250 ;
 wire \i48/n251 ;
 wire \i48/n252 ;
 wire \i48/n253 ;
 wire \i48/n254 ;
 wire \i48/n255 ;
 wire \i48/n256 ;
 wire \i48/n257 ;
 wire \i48/n258 ;
 wire \i48/n259 ;
 wire \i48/n26 ;
 wire \i48/n260 ;
 wire \i48/n261 ;
 wire \i48/n262 ;
 wire \i48/n263 ;
 wire \i48/n264 ;
 wire \i48/n265 ;
 wire \i48/n266 ;
 wire \i48/n267 ;
 wire \i48/n268 ;
 wire \i48/n269 ;
 wire \i48/n27 ;
 wire \i48/n270 ;
 wire \i48/n271 ;
 wire \i48/n272 ;
 wire \i48/n273 ;
 wire \i48/n274 ;
 wire \i48/n275 ;
 wire \i48/n276 ;
 wire \i48/n277 ;
 wire \i48/n278 ;
 wire \i48/n279 ;
 wire \i48/n28 ;
 wire \i48/n280 ;
 wire \i48/n281 ;
 wire \i48/n282 ;
 wire \i48/n283 ;
 wire \i48/n284 ;
 wire \i48/n285 ;
 wire \i48/n286 ;
 wire \i48/n287 ;
 wire \i48/n288 ;
 wire \i48/n289 ;
 wire \i48/n29 ;
 wire \i48/n290 ;
 wire \i48/n291 ;
 wire \i48/n292 ;
 wire \i48/n293 ;
 wire \i48/n294 ;
 wire \i48/n295 ;
 wire \i48/n296 ;
 wire \i48/n297 ;
 wire \i48/n298 ;
 wire \i48/n299 ;
 wire \i48/n3 ;
 wire \i48/n30 ;
 wire \i48/n300 ;
 wire \i48/n301 ;
 wire \i48/n302 ;
 wire \i48/n303 ;
 wire \i48/n304 ;
 wire \i48/n305 ;
 wire \i48/n306 ;
 wire \i48/n307 ;
 wire \i48/n308 ;
 wire \i48/n309 ;
 wire \i48/n31 ;
 wire \i48/n310 ;
 wire \i48/n311 ;
 wire \i48/n312 ;
 wire \i48/n313 ;
 wire \i48/n314 ;
 wire \i48/n315 ;
 wire \i48/n316 ;
 wire \i48/n317 ;
 wire \i48/n318 ;
 wire \i48/n319 ;
 wire \i48/n32 ;
 wire \i48/n320 ;
 wire \i48/n321 ;
 wire \i48/n322 ;
 wire \i48/n323 ;
 wire \i48/n324 ;
 wire \i48/n325 ;
 wire \i48/n326 ;
 wire \i48/n327 ;
 wire \i48/n328 ;
 wire \i48/n329 ;
 wire \i48/n33 ;
 wire \i48/n330 ;
 wire \i48/n331 ;
 wire \i48/n332 ;
 wire \i48/n333 ;
 wire \i48/n334 ;
 wire \i48/n335 ;
 wire \i48/n336 ;
 wire \i48/n337 ;
 wire \i48/n338 ;
 wire \i48/n339 ;
 wire \i48/n34 ;
 wire \i48/n340 ;
 wire \i48/n341 ;
 wire \i48/n342 ;
 wire \i48/n343 ;
 wire \i48/n344 ;
 wire \i48/n345 ;
 wire \i48/n346 ;
 wire \i48/n347 ;
 wire \i48/n348 ;
 wire \i48/n349 ;
 wire \i48/n35 ;
 wire \i48/n350 ;
 wire \i48/n351 ;
 wire \i48/n352 ;
 wire \i48/n353 ;
 wire \i48/n354 ;
 wire \i48/n355 ;
 wire \i48/n356 ;
 wire \i48/n357 ;
 wire \i48/n358 ;
 wire \i48/n359 ;
 wire \i48/n36 ;
 wire \i48/n360 ;
 wire \i48/n361 ;
 wire \i48/n362 ;
 wire \i48/n363 ;
 wire \i48/n364 ;
 wire \i48/n365 ;
 wire \i48/n366 ;
 wire \i48/n367 ;
 wire \i48/n368 ;
 wire \i48/n369 ;
 wire \i48/n37 ;
 wire \i48/n370 ;
 wire \i48/n371 ;
 wire \i48/n372 ;
 wire \i48/n373 ;
 wire \i48/n374 ;
 wire \i48/n375 ;
 wire \i48/n376 ;
 wire \i48/n377 ;
 wire \i48/n378 ;
 wire \i48/n379 ;
 wire \i48/n38 ;
 wire \i48/n380 ;
 wire \i48/n381 ;
 wire \i48/n382 ;
 wire \i48/n383 ;
 wire \i48/n384 ;
 wire \i48/n385 ;
 wire \i48/n386 ;
 wire \i48/n387 ;
 wire \i48/n388 ;
 wire \i48/n389 ;
 wire \i48/n39 ;
 wire \i48/n390 ;
 wire \i48/n391 ;
 wire \i48/n392 ;
 wire \i48/n393 ;
 wire \i48/n394 ;
 wire \i48/n395 ;
 wire \i48/n396 ;
 wire \i48/n397 ;
 wire \i48/n398 ;
 wire \i48/n399 ;
 wire \i48/n4 ;
 wire \i48/n40 ;
 wire \i48/n400 ;
 wire \i48/n401 ;
 wire \i48/n402 ;
 wire \i48/n403 ;
 wire \i48/n404 ;
 wire \i48/n405 ;
 wire \i48/n406 ;
 wire \i48/n407 ;
 wire \i48/n408 ;
 wire \i48/n409 ;
 wire \i48/n41 ;
 wire \i48/n410 ;
 wire \i48/n411 ;
 wire \i48/n412 ;
 wire \i48/n413 ;
 wire \i48/n414 ;
 wire \i48/n415 ;
 wire \i48/n416 ;
 wire \i48/n417 ;
 wire \i48/n418 ;
 wire \i48/n419 ;
 wire \i48/n42 ;
 wire \i48/n420 ;
 wire \i48/n421 ;
 wire \i48/n422 ;
 wire \i48/n423 ;
 wire \i48/n424 ;
 wire \i48/n425 ;
 wire \i48/n426 ;
 wire \i48/n427 ;
 wire \i48/n428 ;
 wire \i48/n429 ;
 wire \i48/n43 ;
 wire \i48/n430 ;
 wire \i48/n431 ;
 wire \i48/n432 ;
 wire \i48/n433 ;
 wire \i48/n434 ;
 wire \i48/n435 ;
 wire \i48/n436 ;
 wire \i48/n437 ;
 wire \i48/n438 ;
 wire \i48/n439 ;
 wire \i48/n44 ;
 wire \i48/n440 ;
 wire \i48/n441 ;
 wire \i48/n442 ;
 wire \i48/n443 ;
 wire \i48/n444 ;
 wire \i48/n445 ;
 wire \i48/n446 ;
 wire \i48/n447 ;
 wire \i48/n448 ;
 wire \i48/n449 ;
 wire \i48/n45 ;
 wire \i48/n450 ;
 wire \i48/n451 ;
 wire \i48/n452 ;
 wire \i48/n453 ;
 wire \i48/n454 ;
 wire \i48/n455 ;
 wire \i48/n456 ;
 wire \i48/n457 ;
 wire \i48/n458 ;
 wire \i48/n459 ;
 wire \i48/n46 ;
 wire \i48/n460 ;
 wire \i48/n461 ;
 wire \i48/n462 ;
 wire \i48/n463 ;
 wire \i48/n464 ;
 wire \i48/n465 ;
 wire \i48/n466 ;
 wire \i48/n467 ;
 wire \i48/n468 ;
 wire \i48/n469 ;
 wire \i48/n47 ;
 wire \i48/n470 ;
 wire \i48/n471 ;
 wire \i48/n472 ;
 wire \i48/n473 ;
 wire \i48/n474 ;
 wire \i48/n475 ;
 wire \i48/n476 ;
 wire \i48/n477 ;
 wire \i48/n478 ;
 wire \i48/n479 ;
 wire \i48/n48 ;
 wire \i48/n480 ;
 wire \i48/n481 ;
 wire \i48/n482 ;
 wire \i48/n483 ;
 wire \i48/n484 ;
 wire \i48/n485 ;
 wire \i48/n486 ;
 wire \i48/n487 ;
 wire \i48/n488 ;
 wire \i48/n489 ;
 wire \i48/n49 ;
 wire \i48/n490 ;
 wire \i48/n491 ;
 wire \i48/n492 ;
 wire \i48/n493 ;
 wire \i48/n494 ;
 wire \i48/n495 ;
 wire \i48/n496 ;
 wire \i48/n497 ;
 wire \i48/n498 ;
 wire \i48/n499 ;
 wire \i48/n5 ;
 wire \i48/n50 ;
 wire \i48/n500 ;
 wire \i48/n501 ;
 wire \i48/n502 ;
 wire \i48/n503 ;
 wire \i48/n504 ;
 wire \i48/n505 ;
 wire \i48/n506 ;
 wire \i48/n507 ;
 wire \i48/n508 ;
 wire \i48/n509 ;
 wire \i48/n51 ;
 wire \i48/n510 ;
 wire \i48/n511 ;
 wire \i48/n512 ;
 wire \i48/n513 ;
 wire \i48/n514 ;
 wire \i48/n515 ;
 wire \i48/n516 ;
 wire \i48/n517 ;
 wire \i48/n518 ;
 wire \i48/n519 ;
 wire \i48/n52 ;
 wire \i48/n520 ;
 wire \i48/n521 ;
 wire \i48/n522 ;
 wire \i48/n523 ;
 wire \i48/n524 ;
 wire \i48/n525 ;
 wire \i48/n526 ;
 wire \i48/n527 ;
 wire \i48/n528 ;
 wire \i48/n529 ;
 wire \i48/n53 ;
 wire \i48/n530 ;
 wire \i48/n531 ;
 wire \i48/n532 ;
 wire \i48/n533 ;
 wire \i48/n534 ;
 wire \i48/n535 ;
 wire \i48/n536 ;
 wire \i48/n537 ;
 wire \i48/n538 ;
 wire \i48/n539 ;
 wire \i48/n54 ;
 wire \i48/n540 ;
 wire \i48/n541 ;
 wire \i48/n542 ;
 wire \i48/n543 ;
 wire \i48/n544 ;
 wire \i48/n545 ;
 wire \i48/n546 ;
 wire \i48/n547 ;
 wire \i48/n548 ;
 wire \i48/n549 ;
 wire \i48/n55 ;
 wire \i48/n550 ;
 wire \i48/n551 ;
 wire \i48/n552 ;
 wire \i48/n553 ;
 wire \i48/n554 ;
 wire \i48/n555 ;
 wire \i48/n556 ;
 wire \i48/n557 ;
 wire \i48/n558 ;
 wire \i48/n559 ;
 wire \i48/n56 ;
 wire \i48/n560 ;
 wire \i48/n561 ;
 wire \i48/n562 ;
 wire \i48/n563 ;
 wire \i48/n564 ;
 wire \i48/n565 ;
 wire \i48/n566 ;
 wire \i48/n567 ;
 wire \i48/n568 ;
 wire \i48/n569 ;
 wire \i48/n57 ;
 wire \i48/n570 ;
 wire \i48/n571 ;
 wire \i48/n572 ;
 wire \i48/n573 ;
 wire \i48/n574 ;
 wire \i48/n575 ;
 wire \i48/n576 ;
 wire \i48/n577 ;
 wire \i48/n578 ;
 wire \i48/n579 ;
 wire \i48/n58 ;
 wire \i48/n580 ;
 wire \i48/n581 ;
 wire \i48/n59 ;
 wire \i48/n6 ;
 wire \i48/n60 ;
 wire \i48/n61 ;
 wire \i48/n62 ;
 wire \i48/n63 ;
 wire \i48/n64 ;
 wire \i48/n65 ;
 wire \i48/n66 ;
 wire \i48/n67 ;
 wire \i48/n68 ;
 wire \i48/n69 ;
 wire \i48/n7 ;
 wire \i48/n70 ;
 wire \i48/n71 ;
 wire \i48/n72 ;
 wire \i48/n73 ;
 wire \i48/n74 ;
 wire \i48/n75 ;
 wire \i48/n76 ;
 wire \i48/n77 ;
 wire \i48/n78 ;
 wire \i48/n79 ;
 wire \i48/n8 ;
 wire \i48/n80 ;
 wire \i48/n81 ;
 wire \i48/n82 ;
 wire \i48/n83 ;
 wire \i48/n84 ;
 wire \i48/n85 ;
 wire \i48/n86 ;
 wire \i48/n87 ;
 wire \i48/n88 ;
 wire \i48/n89 ;
 wire \i48/n9 ;
 wire \i48/n90 ;
 wire \i48/n91 ;
 wire \i48/n92 ;
 wire \i48/n93 ;
 wire \i48/n94 ;
 wire \i48/n95 ;
 wire \i48/n96 ;
 wire \i48/n97 ;
 wire \i48/n98 ;
 wire \i48/n99 ;
 wire \i49/n0 ;
 wire \i49/n1 ;
 wire \i49/n10 ;
 wire \i49/n100 ;
 wire \i49/n101 ;
 wire \i49/n102 ;
 wire \i49/n103 ;
 wire \i49/n104 ;
 wire \i49/n105 ;
 wire \i49/n106 ;
 wire \i49/n107 ;
 wire \i49/n108 ;
 wire \i49/n109 ;
 wire \i49/n11 ;
 wire \i49/n110 ;
 wire \i49/n111 ;
 wire \i49/n112 ;
 wire \i49/n113 ;
 wire \i49/n114 ;
 wire \i49/n115 ;
 wire \i49/n116 ;
 wire \i49/n117 ;
 wire \i49/n118 ;
 wire \i49/n119 ;
 wire \i49/n12 ;
 wire \i49/n120 ;
 wire \i49/n121 ;
 wire \i49/n122 ;
 wire \i49/n123 ;
 wire \i49/n124 ;
 wire \i49/n125 ;
 wire \i49/n126 ;
 wire \i49/n127 ;
 wire \i49/n128 ;
 wire \i49/n129 ;
 wire \i49/n13 ;
 wire \i49/n130 ;
 wire \i49/n131 ;
 wire \i49/n132 ;
 wire \i49/n133 ;
 wire \i49/n134 ;
 wire \i49/n135 ;
 wire \i49/n136 ;
 wire \i49/n137 ;
 wire \i49/n138 ;
 wire \i49/n139 ;
 wire \i49/n14 ;
 wire \i49/n140 ;
 wire \i49/n141 ;
 wire \i49/n142 ;
 wire \i49/n143 ;
 wire \i49/n144 ;
 wire \i49/n145 ;
 wire \i49/n146 ;
 wire \i49/n147 ;
 wire \i49/n148 ;
 wire \i49/n149 ;
 wire \i49/n15 ;
 wire \i49/n150 ;
 wire \i49/n151 ;
 wire \i49/n152 ;
 wire \i49/n153 ;
 wire \i49/n154 ;
 wire \i49/n155 ;
 wire \i49/n156 ;
 wire \i49/n157 ;
 wire \i49/n158 ;
 wire \i49/n159 ;
 wire \i49/n16 ;
 wire \i49/n160 ;
 wire \i49/n161 ;
 wire \i49/n162 ;
 wire \i49/n163 ;
 wire \i49/n164 ;
 wire \i49/n165 ;
 wire \i49/n166 ;
 wire \i49/n167 ;
 wire \i49/n168 ;
 wire \i49/n169 ;
 wire \i49/n17 ;
 wire \i49/n170 ;
 wire \i49/n171 ;
 wire \i49/n172 ;
 wire \i49/n173 ;
 wire \i49/n174 ;
 wire \i49/n175 ;
 wire \i49/n176 ;
 wire \i49/n177 ;
 wire \i49/n178 ;
 wire \i49/n179 ;
 wire \i49/n18 ;
 wire \i49/n180 ;
 wire \i49/n181 ;
 wire \i49/n182 ;
 wire \i49/n183 ;
 wire \i49/n184 ;
 wire \i49/n185 ;
 wire \i49/n186 ;
 wire \i49/n187 ;
 wire \i49/n188 ;
 wire \i49/n189 ;
 wire \i49/n19 ;
 wire \i49/n190 ;
 wire \i49/n191 ;
 wire \i49/n192 ;
 wire \i49/n193 ;
 wire \i49/n194 ;
 wire \i49/n195 ;
 wire \i49/n196 ;
 wire \i49/n197 ;
 wire \i49/n198 ;
 wire \i49/n199 ;
 wire \i49/n2 ;
 wire \i49/n20 ;
 wire \i49/n200 ;
 wire \i49/n201 ;
 wire \i49/n202 ;
 wire \i49/n203 ;
 wire \i49/n204 ;
 wire \i49/n205 ;
 wire \i49/n206 ;
 wire \i49/n207 ;
 wire \i49/n208 ;
 wire \i49/n209 ;
 wire \i49/n21 ;
 wire \i49/n210 ;
 wire \i49/n211 ;
 wire \i49/n212 ;
 wire \i49/n213 ;
 wire \i49/n214 ;
 wire \i49/n215 ;
 wire \i49/n216 ;
 wire \i49/n217 ;
 wire \i49/n218 ;
 wire \i49/n219 ;
 wire \i49/n22 ;
 wire \i49/n220 ;
 wire \i49/n221 ;
 wire \i49/n222 ;
 wire \i49/n223 ;
 wire \i49/n224 ;
 wire \i49/n225 ;
 wire \i49/n226 ;
 wire \i49/n227 ;
 wire \i49/n228 ;
 wire \i49/n229 ;
 wire \i49/n23 ;
 wire \i49/n230 ;
 wire \i49/n231 ;
 wire \i49/n232 ;
 wire \i49/n233 ;
 wire \i49/n234 ;
 wire \i49/n235 ;
 wire \i49/n236 ;
 wire \i49/n237 ;
 wire \i49/n238 ;
 wire \i49/n239 ;
 wire \i49/n24 ;
 wire \i49/n240 ;
 wire \i49/n241 ;
 wire \i49/n242 ;
 wire \i49/n243 ;
 wire \i49/n244 ;
 wire \i49/n245 ;
 wire \i49/n246 ;
 wire \i49/n247 ;
 wire \i49/n248 ;
 wire \i49/n249 ;
 wire \i49/n25 ;
 wire \i49/n250 ;
 wire \i49/n251 ;
 wire \i49/n252 ;
 wire \i49/n253 ;
 wire \i49/n254 ;
 wire \i49/n255 ;
 wire \i49/n256 ;
 wire \i49/n257 ;
 wire \i49/n258 ;
 wire \i49/n259 ;
 wire \i49/n26 ;
 wire \i49/n260 ;
 wire \i49/n261 ;
 wire \i49/n262 ;
 wire \i49/n263 ;
 wire \i49/n264 ;
 wire \i49/n265 ;
 wire \i49/n266 ;
 wire \i49/n267 ;
 wire \i49/n268 ;
 wire \i49/n269 ;
 wire \i49/n27 ;
 wire \i49/n270 ;
 wire \i49/n271 ;
 wire \i49/n272 ;
 wire \i49/n273 ;
 wire \i49/n274 ;
 wire \i49/n275 ;
 wire \i49/n276 ;
 wire \i49/n277 ;
 wire \i49/n278 ;
 wire \i49/n279 ;
 wire \i49/n28 ;
 wire \i49/n280 ;
 wire \i49/n281 ;
 wire \i49/n282 ;
 wire \i49/n283 ;
 wire \i49/n284 ;
 wire \i49/n285 ;
 wire \i49/n286 ;
 wire \i49/n287 ;
 wire \i49/n288 ;
 wire \i49/n289 ;
 wire \i49/n29 ;
 wire \i49/n290 ;
 wire \i49/n291 ;
 wire \i49/n292 ;
 wire \i49/n293 ;
 wire \i49/n294 ;
 wire \i49/n295 ;
 wire \i49/n296 ;
 wire \i49/n297 ;
 wire \i49/n298 ;
 wire \i49/n299 ;
 wire \i49/n3 ;
 wire \i49/n30 ;
 wire \i49/n300 ;
 wire \i49/n301 ;
 wire \i49/n302 ;
 wire \i49/n303 ;
 wire \i49/n304 ;
 wire \i49/n305 ;
 wire \i49/n306 ;
 wire \i49/n307 ;
 wire \i49/n308 ;
 wire \i49/n309 ;
 wire \i49/n31 ;
 wire \i49/n310 ;
 wire \i49/n311 ;
 wire \i49/n312 ;
 wire \i49/n313 ;
 wire \i49/n314 ;
 wire \i49/n315 ;
 wire \i49/n316 ;
 wire \i49/n317 ;
 wire \i49/n318 ;
 wire \i49/n319 ;
 wire \i49/n32 ;
 wire \i49/n320 ;
 wire \i49/n321 ;
 wire \i49/n322 ;
 wire \i49/n323 ;
 wire \i49/n324 ;
 wire \i49/n325 ;
 wire \i49/n326 ;
 wire \i49/n327 ;
 wire \i49/n328 ;
 wire \i49/n329 ;
 wire \i49/n33 ;
 wire \i49/n330 ;
 wire \i49/n331 ;
 wire \i49/n332 ;
 wire \i49/n333 ;
 wire \i49/n334 ;
 wire \i49/n335 ;
 wire \i49/n336 ;
 wire \i49/n337 ;
 wire \i49/n338 ;
 wire \i49/n339 ;
 wire \i49/n34 ;
 wire \i49/n340 ;
 wire \i49/n341 ;
 wire \i49/n342 ;
 wire \i49/n343 ;
 wire \i49/n344 ;
 wire \i49/n345 ;
 wire \i49/n346 ;
 wire \i49/n347 ;
 wire \i49/n348 ;
 wire \i49/n349 ;
 wire \i49/n35 ;
 wire \i49/n350 ;
 wire \i49/n351 ;
 wire \i49/n352 ;
 wire \i49/n353 ;
 wire \i49/n354 ;
 wire \i49/n355 ;
 wire \i49/n356 ;
 wire \i49/n357 ;
 wire \i49/n358 ;
 wire \i49/n359 ;
 wire \i49/n36 ;
 wire \i49/n360 ;
 wire \i49/n361 ;
 wire \i49/n362 ;
 wire \i49/n363 ;
 wire \i49/n364 ;
 wire \i49/n365 ;
 wire \i49/n366 ;
 wire \i49/n367 ;
 wire \i49/n368 ;
 wire \i49/n369 ;
 wire \i49/n37 ;
 wire \i49/n370 ;
 wire \i49/n371 ;
 wire \i49/n372 ;
 wire \i49/n373 ;
 wire \i49/n374 ;
 wire \i49/n375 ;
 wire \i49/n376 ;
 wire \i49/n377 ;
 wire \i49/n378 ;
 wire \i49/n379 ;
 wire \i49/n38 ;
 wire \i49/n380 ;
 wire \i49/n381 ;
 wire \i49/n382 ;
 wire \i49/n383 ;
 wire \i49/n384 ;
 wire \i49/n385 ;
 wire \i49/n386 ;
 wire \i49/n387 ;
 wire \i49/n388 ;
 wire \i49/n389 ;
 wire \i49/n39 ;
 wire \i49/n390 ;
 wire \i49/n391 ;
 wire \i49/n392 ;
 wire \i49/n393 ;
 wire \i49/n394 ;
 wire \i49/n395 ;
 wire \i49/n396 ;
 wire \i49/n397 ;
 wire \i49/n398 ;
 wire \i49/n399 ;
 wire \i49/n4 ;
 wire \i49/n40 ;
 wire \i49/n400 ;
 wire \i49/n401 ;
 wire \i49/n402 ;
 wire \i49/n403 ;
 wire \i49/n404 ;
 wire \i49/n405 ;
 wire \i49/n406 ;
 wire \i49/n407 ;
 wire \i49/n408 ;
 wire \i49/n409 ;
 wire \i49/n41 ;
 wire \i49/n410 ;
 wire \i49/n411 ;
 wire \i49/n412 ;
 wire \i49/n413 ;
 wire \i49/n414 ;
 wire \i49/n415 ;
 wire \i49/n416 ;
 wire \i49/n417 ;
 wire \i49/n418 ;
 wire \i49/n419 ;
 wire \i49/n42 ;
 wire \i49/n420 ;
 wire \i49/n421 ;
 wire \i49/n422 ;
 wire \i49/n423 ;
 wire \i49/n424 ;
 wire \i49/n425 ;
 wire \i49/n426 ;
 wire \i49/n427 ;
 wire \i49/n428 ;
 wire \i49/n429 ;
 wire \i49/n43 ;
 wire \i49/n430 ;
 wire \i49/n431 ;
 wire \i49/n432 ;
 wire \i49/n433 ;
 wire \i49/n434 ;
 wire \i49/n435 ;
 wire \i49/n436 ;
 wire \i49/n437 ;
 wire \i49/n438 ;
 wire \i49/n439 ;
 wire \i49/n44 ;
 wire \i49/n440 ;
 wire \i49/n441 ;
 wire \i49/n442 ;
 wire \i49/n443 ;
 wire \i49/n444 ;
 wire \i49/n445 ;
 wire \i49/n446 ;
 wire \i49/n447 ;
 wire \i49/n448 ;
 wire \i49/n449 ;
 wire \i49/n45 ;
 wire \i49/n450 ;
 wire \i49/n451 ;
 wire \i49/n452 ;
 wire \i49/n453 ;
 wire \i49/n454 ;
 wire \i49/n455 ;
 wire \i49/n456 ;
 wire \i49/n457 ;
 wire \i49/n458 ;
 wire \i49/n459 ;
 wire \i49/n46 ;
 wire \i49/n460 ;
 wire \i49/n461 ;
 wire \i49/n462 ;
 wire \i49/n463 ;
 wire \i49/n464 ;
 wire \i49/n465 ;
 wire \i49/n466 ;
 wire \i49/n467 ;
 wire \i49/n468 ;
 wire \i49/n469 ;
 wire \i49/n47 ;
 wire \i49/n470 ;
 wire \i49/n471 ;
 wire \i49/n472 ;
 wire \i49/n473 ;
 wire \i49/n474 ;
 wire \i49/n475 ;
 wire \i49/n476 ;
 wire \i49/n477 ;
 wire \i49/n478 ;
 wire \i49/n479 ;
 wire \i49/n48 ;
 wire \i49/n480 ;
 wire \i49/n481 ;
 wire \i49/n482 ;
 wire \i49/n483 ;
 wire \i49/n484 ;
 wire \i49/n485 ;
 wire \i49/n486 ;
 wire \i49/n487 ;
 wire \i49/n488 ;
 wire \i49/n489 ;
 wire \i49/n49 ;
 wire \i49/n490 ;
 wire \i49/n491 ;
 wire \i49/n492 ;
 wire \i49/n493 ;
 wire \i49/n494 ;
 wire \i49/n495 ;
 wire \i49/n496 ;
 wire \i49/n497 ;
 wire \i49/n498 ;
 wire \i49/n499 ;
 wire \i49/n5 ;
 wire \i49/n50 ;
 wire \i49/n500 ;
 wire \i49/n501 ;
 wire \i49/n502 ;
 wire \i49/n503 ;
 wire \i49/n504 ;
 wire \i49/n505 ;
 wire \i49/n506 ;
 wire \i49/n507 ;
 wire \i49/n508 ;
 wire \i49/n509 ;
 wire \i49/n51 ;
 wire \i49/n510 ;
 wire \i49/n511 ;
 wire \i49/n512 ;
 wire \i49/n513 ;
 wire \i49/n514 ;
 wire \i49/n515 ;
 wire \i49/n516 ;
 wire \i49/n517 ;
 wire \i49/n518 ;
 wire \i49/n519 ;
 wire \i49/n52 ;
 wire \i49/n520 ;
 wire \i49/n521 ;
 wire \i49/n522 ;
 wire \i49/n523 ;
 wire \i49/n524 ;
 wire \i49/n525 ;
 wire \i49/n526 ;
 wire \i49/n527 ;
 wire \i49/n528 ;
 wire \i49/n529 ;
 wire \i49/n53 ;
 wire \i49/n530 ;
 wire \i49/n531 ;
 wire \i49/n532 ;
 wire \i49/n533 ;
 wire \i49/n534 ;
 wire \i49/n535 ;
 wire \i49/n536 ;
 wire \i49/n537 ;
 wire \i49/n538 ;
 wire \i49/n539 ;
 wire \i49/n54 ;
 wire \i49/n540 ;
 wire \i49/n541 ;
 wire \i49/n542 ;
 wire \i49/n543 ;
 wire \i49/n544 ;
 wire \i49/n545 ;
 wire \i49/n546 ;
 wire \i49/n547 ;
 wire \i49/n548 ;
 wire \i49/n549 ;
 wire \i49/n55 ;
 wire \i49/n550 ;
 wire \i49/n551 ;
 wire \i49/n552 ;
 wire \i49/n553 ;
 wire \i49/n554 ;
 wire \i49/n555 ;
 wire \i49/n556 ;
 wire \i49/n557 ;
 wire \i49/n558 ;
 wire \i49/n559 ;
 wire \i49/n56 ;
 wire \i49/n560 ;
 wire \i49/n561 ;
 wire \i49/n562 ;
 wire \i49/n563 ;
 wire \i49/n564 ;
 wire \i49/n565 ;
 wire \i49/n566 ;
 wire \i49/n567 ;
 wire \i49/n568 ;
 wire \i49/n569 ;
 wire \i49/n57 ;
 wire \i49/n570 ;
 wire \i49/n571 ;
 wire \i49/n572 ;
 wire \i49/n573 ;
 wire \i49/n574 ;
 wire \i49/n575 ;
 wire \i49/n576 ;
 wire \i49/n577 ;
 wire \i49/n578 ;
 wire \i49/n579 ;
 wire \i49/n58 ;
 wire \i49/n580 ;
 wire \i49/n581 ;
 wire \i49/n59 ;
 wire \i49/n6 ;
 wire \i49/n60 ;
 wire \i49/n61 ;
 wire \i49/n62 ;
 wire \i49/n63 ;
 wire \i49/n64 ;
 wire \i49/n65 ;
 wire \i49/n66 ;
 wire \i49/n67 ;
 wire \i49/n68 ;
 wire \i49/n69 ;
 wire \i49/n7 ;
 wire \i49/n70 ;
 wire \i49/n71 ;
 wire \i49/n72 ;
 wire \i49/n73 ;
 wire \i49/n74 ;
 wire \i49/n75 ;
 wire \i49/n76 ;
 wire \i49/n77 ;
 wire \i49/n78 ;
 wire \i49/n79 ;
 wire \i49/n8 ;
 wire \i49/n80 ;
 wire \i49/n81 ;
 wire \i49/n82 ;
 wire \i49/n83 ;
 wire \i49/n84 ;
 wire \i49/n85 ;
 wire \i49/n86 ;
 wire \i49/n87 ;
 wire \i49/n88 ;
 wire \i49/n89 ;
 wire \i49/n9 ;
 wire \i49/n90 ;
 wire \i49/n91 ;
 wire \i49/n92 ;
 wire \i49/n93 ;
 wire \i49/n94 ;
 wire \i49/n95 ;
 wire \i49/n96 ;
 wire \i49/n97 ;
 wire \i49/n98 ;
 wire \i49/n99 ;
 wire \i50/n0 ;
 wire \i50/n1 ;
 wire \i50/n10 ;
 wire \i50/n100 ;
 wire \i50/n101 ;
 wire \i50/n102 ;
 wire \i50/n103 ;
 wire \i50/n104 ;
 wire \i50/n105 ;
 wire \i50/n106 ;
 wire \i50/n107 ;
 wire \i50/n108 ;
 wire \i50/n109 ;
 wire \i50/n11 ;
 wire \i50/n110 ;
 wire \i50/n111 ;
 wire \i50/n112 ;
 wire \i50/n113 ;
 wire \i50/n114 ;
 wire \i50/n115 ;
 wire \i50/n116 ;
 wire \i50/n117 ;
 wire \i50/n118 ;
 wire \i50/n119 ;
 wire \i50/n12 ;
 wire \i50/n120 ;
 wire \i50/n121 ;
 wire \i50/n122 ;
 wire \i50/n123 ;
 wire \i50/n124 ;
 wire \i50/n125 ;
 wire \i50/n126 ;
 wire \i50/n127 ;
 wire \i50/n128 ;
 wire \i50/n129 ;
 wire \i50/n13 ;
 wire \i50/n130 ;
 wire \i50/n131 ;
 wire \i50/n132 ;
 wire \i50/n133 ;
 wire \i50/n134 ;
 wire \i50/n135 ;
 wire \i50/n136 ;
 wire \i50/n137 ;
 wire \i50/n138 ;
 wire \i50/n139 ;
 wire \i50/n14 ;
 wire \i50/n140 ;
 wire \i50/n141 ;
 wire \i50/n142 ;
 wire \i50/n143 ;
 wire \i50/n144 ;
 wire \i50/n145 ;
 wire \i50/n146 ;
 wire \i50/n147 ;
 wire \i50/n148 ;
 wire \i50/n149 ;
 wire \i50/n15 ;
 wire \i50/n150 ;
 wire \i50/n151 ;
 wire \i50/n152 ;
 wire \i50/n153 ;
 wire \i50/n154 ;
 wire \i50/n155 ;
 wire \i50/n156 ;
 wire \i50/n157 ;
 wire \i50/n158 ;
 wire \i50/n159 ;
 wire \i50/n16 ;
 wire \i50/n160 ;
 wire \i50/n161 ;
 wire \i50/n162 ;
 wire \i50/n163 ;
 wire \i50/n164 ;
 wire \i50/n165 ;
 wire \i50/n166 ;
 wire \i50/n167 ;
 wire \i50/n168 ;
 wire \i50/n169 ;
 wire \i50/n17 ;
 wire \i50/n170 ;
 wire \i50/n171 ;
 wire \i50/n172 ;
 wire \i50/n173 ;
 wire \i50/n174 ;
 wire \i50/n175 ;
 wire \i50/n176 ;
 wire \i50/n177 ;
 wire \i50/n178 ;
 wire \i50/n179 ;
 wire \i50/n18 ;
 wire \i50/n180 ;
 wire \i50/n181 ;
 wire \i50/n182 ;
 wire \i50/n183 ;
 wire \i50/n184 ;
 wire \i50/n185 ;
 wire \i50/n186 ;
 wire \i50/n187 ;
 wire \i50/n188 ;
 wire \i50/n189 ;
 wire \i50/n19 ;
 wire \i50/n190 ;
 wire \i50/n191 ;
 wire \i50/n192 ;
 wire \i50/n193 ;
 wire \i50/n194 ;
 wire \i50/n195 ;
 wire \i50/n196 ;
 wire \i50/n197 ;
 wire \i50/n198 ;
 wire \i50/n199 ;
 wire \i50/n2 ;
 wire \i50/n20 ;
 wire \i50/n200 ;
 wire \i50/n201 ;
 wire \i50/n202 ;
 wire \i50/n203 ;
 wire \i50/n204 ;
 wire \i50/n205 ;
 wire \i50/n206 ;
 wire \i50/n207 ;
 wire \i50/n208 ;
 wire \i50/n209 ;
 wire \i50/n21 ;
 wire \i50/n210 ;
 wire \i50/n211 ;
 wire \i50/n212 ;
 wire \i50/n213 ;
 wire \i50/n214 ;
 wire \i50/n215 ;
 wire \i50/n216 ;
 wire \i50/n217 ;
 wire \i50/n218 ;
 wire \i50/n219 ;
 wire \i50/n22 ;
 wire \i50/n220 ;
 wire \i50/n221 ;
 wire \i50/n222 ;
 wire \i50/n223 ;
 wire \i50/n224 ;
 wire \i50/n225 ;
 wire \i50/n226 ;
 wire \i50/n227 ;
 wire \i50/n228 ;
 wire \i50/n229 ;
 wire \i50/n23 ;
 wire \i50/n230 ;
 wire \i50/n231 ;
 wire \i50/n232 ;
 wire \i50/n233 ;
 wire \i50/n234 ;
 wire \i50/n235 ;
 wire \i50/n236 ;
 wire \i50/n237 ;
 wire \i50/n238 ;
 wire \i50/n239 ;
 wire \i50/n24 ;
 wire \i50/n240 ;
 wire \i50/n241 ;
 wire \i50/n242 ;
 wire \i50/n243 ;
 wire \i50/n244 ;
 wire \i50/n245 ;
 wire \i50/n246 ;
 wire \i50/n247 ;
 wire \i50/n248 ;
 wire \i50/n249 ;
 wire \i50/n25 ;
 wire \i50/n250 ;
 wire \i50/n251 ;
 wire \i50/n252 ;
 wire \i50/n253 ;
 wire \i50/n254 ;
 wire \i50/n255 ;
 wire \i50/n256 ;
 wire \i50/n257 ;
 wire \i50/n258 ;
 wire \i50/n259 ;
 wire \i50/n26 ;
 wire \i50/n260 ;
 wire \i50/n261 ;
 wire \i50/n262 ;
 wire \i50/n263 ;
 wire \i50/n264 ;
 wire \i50/n265 ;
 wire \i50/n266 ;
 wire \i50/n267 ;
 wire \i50/n268 ;
 wire \i50/n269 ;
 wire \i50/n27 ;
 wire \i50/n270 ;
 wire \i50/n271 ;
 wire \i50/n272 ;
 wire \i50/n273 ;
 wire \i50/n274 ;
 wire \i50/n275 ;
 wire \i50/n276 ;
 wire \i50/n277 ;
 wire \i50/n278 ;
 wire \i50/n279 ;
 wire \i50/n28 ;
 wire \i50/n280 ;
 wire \i50/n281 ;
 wire \i50/n282 ;
 wire \i50/n283 ;
 wire \i50/n284 ;
 wire \i50/n285 ;
 wire \i50/n286 ;
 wire \i50/n287 ;
 wire \i50/n288 ;
 wire \i50/n289 ;
 wire \i50/n29 ;
 wire \i50/n290 ;
 wire \i50/n291 ;
 wire \i50/n292 ;
 wire \i50/n293 ;
 wire \i50/n294 ;
 wire \i50/n295 ;
 wire \i50/n296 ;
 wire \i50/n297 ;
 wire \i50/n298 ;
 wire \i50/n299 ;
 wire \i50/n3 ;
 wire \i50/n30 ;
 wire \i50/n300 ;
 wire \i50/n301 ;
 wire \i50/n302 ;
 wire \i50/n303 ;
 wire \i50/n304 ;
 wire \i50/n305 ;
 wire \i50/n306 ;
 wire \i50/n307 ;
 wire \i50/n308 ;
 wire \i50/n309 ;
 wire \i50/n31 ;
 wire \i50/n310 ;
 wire \i50/n311 ;
 wire \i50/n312 ;
 wire \i50/n313 ;
 wire \i50/n314 ;
 wire \i50/n315 ;
 wire \i50/n316 ;
 wire \i50/n317 ;
 wire \i50/n318 ;
 wire \i50/n319 ;
 wire \i50/n32 ;
 wire \i50/n320 ;
 wire \i50/n321 ;
 wire \i50/n322 ;
 wire \i50/n323 ;
 wire \i50/n324 ;
 wire \i50/n325 ;
 wire \i50/n326 ;
 wire \i50/n327 ;
 wire \i50/n328 ;
 wire \i50/n329 ;
 wire \i50/n33 ;
 wire \i50/n330 ;
 wire \i50/n331 ;
 wire \i50/n332 ;
 wire \i50/n333 ;
 wire \i50/n334 ;
 wire \i50/n335 ;
 wire \i50/n336 ;
 wire \i50/n337 ;
 wire \i50/n338 ;
 wire \i50/n339 ;
 wire \i50/n34 ;
 wire \i50/n340 ;
 wire \i50/n341 ;
 wire \i50/n342 ;
 wire \i50/n343 ;
 wire \i50/n344 ;
 wire \i50/n345 ;
 wire \i50/n346 ;
 wire \i50/n347 ;
 wire \i50/n348 ;
 wire \i50/n349 ;
 wire \i50/n35 ;
 wire \i50/n350 ;
 wire \i50/n351 ;
 wire \i50/n352 ;
 wire \i50/n353 ;
 wire \i50/n354 ;
 wire \i50/n355 ;
 wire \i50/n356 ;
 wire \i50/n357 ;
 wire \i50/n358 ;
 wire \i50/n359 ;
 wire \i50/n36 ;
 wire \i50/n360 ;
 wire \i50/n361 ;
 wire \i50/n362 ;
 wire \i50/n363 ;
 wire \i50/n364 ;
 wire \i50/n365 ;
 wire \i50/n366 ;
 wire \i50/n367 ;
 wire \i50/n368 ;
 wire \i50/n369 ;
 wire \i50/n37 ;
 wire \i50/n370 ;
 wire \i50/n371 ;
 wire \i50/n372 ;
 wire \i50/n373 ;
 wire \i50/n374 ;
 wire \i50/n375 ;
 wire \i50/n376 ;
 wire \i50/n377 ;
 wire \i50/n378 ;
 wire \i50/n379 ;
 wire \i50/n38 ;
 wire \i50/n380 ;
 wire \i50/n381 ;
 wire \i50/n382 ;
 wire \i50/n383 ;
 wire \i50/n384 ;
 wire \i50/n385 ;
 wire \i50/n386 ;
 wire \i50/n387 ;
 wire \i50/n388 ;
 wire \i50/n389 ;
 wire \i50/n39 ;
 wire \i50/n390 ;
 wire \i50/n391 ;
 wire \i50/n392 ;
 wire \i50/n393 ;
 wire \i50/n394 ;
 wire \i50/n395 ;
 wire \i50/n396 ;
 wire \i50/n397 ;
 wire \i50/n398 ;
 wire \i50/n399 ;
 wire \i50/n4 ;
 wire \i50/n40 ;
 wire \i50/n400 ;
 wire \i50/n401 ;
 wire \i50/n402 ;
 wire \i50/n403 ;
 wire \i50/n404 ;
 wire \i50/n405 ;
 wire \i50/n406 ;
 wire \i50/n407 ;
 wire \i50/n408 ;
 wire \i50/n409 ;
 wire \i50/n41 ;
 wire \i50/n410 ;
 wire \i50/n411 ;
 wire \i50/n412 ;
 wire \i50/n413 ;
 wire \i50/n414 ;
 wire \i50/n415 ;
 wire \i50/n416 ;
 wire \i50/n417 ;
 wire \i50/n418 ;
 wire \i50/n419 ;
 wire \i50/n42 ;
 wire \i50/n420 ;
 wire \i50/n421 ;
 wire \i50/n422 ;
 wire \i50/n423 ;
 wire \i50/n424 ;
 wire \i50/n425 ;
 wire \i50/n426 ;
 wire \i50/n427 ;
 wire \i50/n428 ;
 wire \i50/n429 ;
 wire \i50/n43 ;
 wire \i50/n430 ;
 wire \i50/n431 ;
 wire \i50/n432 ;
 wire \i50/n433 ;
 wire \i50/n434 ;
 wire \i50/n435 ;
 wire \i50/n436 ;
 wire \i50/n437 ;
 wire \i50/n438 ;
 wire \i50/n439 ;
 wire \i50/n44 ;
 wire \i50/n440 ;
 wire \i50/n441 ;
 wire \i50/n442 ;
 wire \i50/n443 ;
 wire \i50/n444 ;
 wire \i50/n445 ;
 wire \i50/n446 ;
 wire \i50/n447 ;
 wire \i50/n448 ;
 wire \i50/n449 ;
 wire \i50/n45 ;
 wire \i50/n450 ;
 wire \i50/n451 ;
 wire \i50/n452 ;
 wire \i50/n453 ;
 wire \i50/n454 ;
 wire \i50/n455 ;
 wire \i50/n456 ;
 wire \i50/n457 ;
 wire \i50/n458 ;
 wire \i50/n459 ;
 wire \i50/n46 ;
 wire \i50/n460 ;
 wire \i50/n461 ;
 wire \i50/n462 ;
 wire \i50/n463 ;
 wire \i50/n464 ;
 wire \i50/n465 ;
 wire \i50/n466 ;
 wire \i50/n467 ;
 wire \i50/n468 ;
 wire \i50/n469 ;
 wire \i50/n47 ;
 wire \i50/n470 ;
 wire \i50/n471 ;
 wire \i50/n472 ;
 wire \i50/n473 ;
 wire \i50/n474 ;
 wire \i50/n475 ;
 wire \i50/n476 ;
 wire \i50/n477 ;
 wire \i50/n478 ;
 wire \i50/n479 ;
 wire \i50/n48 ;
 wire \i50/n480 ;
 wire \i50/n481 ;
 wire \i50/n482 ;
 wire \i50/n483 ;
 wire \i50/n484 ;
 wire \i50/n485 ;
 wire \i50/n486 ;
 wire \i50/n487 ;
 wire \i50/n488 ;
 wire \i50/n489 ;
 wire \i50/n49 ;
 wire \i50/n490 ;
 wire \i50/n491 ;
 wire \i50/n492 ;
 wire \i50/n493 ;
 wire \i50/n494 ;
 wire \i50/n495 ;
 wire \i50/n496 ;
 wire \i50/n497 ;
 wire \i50/n498 ;
 wire \i50/n499 ;
 wire \i50/n5 ;
 wire \i50/n50 ;
 wire \i50/n500 ;
 wire \i50/n501 ;
 wire \i50/n502 ;
 wire \i50/n503 ;
 wire \i50/n504 ;
 wire \i50/n505 ;
 wire \i50/n506 ;
 wire \i50/n507 ;
 wire \i50/n508 ;
 wire \i50/n509 ;
 wire \i50/n51 ;
 wire \i50/n510 ;
 wire \i50/n511 ;
 wire \i50/n512 ;
 wire \i50/n513 ;
 wire \i50/n514 ;
 wire \i50/n515 ;
 wire \i50/n516 ;
 wire \i50/n517 ;
 wire \i50/n518 ;
 wire \i50/n519 ;
 wire \i50/n52 ;
 wire \i50/n520 ;
 wire \i50/n521 ;
 wire \i50/n522 ;
 wire \i50/n523 ;
 wire \i50/n524 ;
 wire \i50/n525 ;
 wire \i50/n526 ;
 wire \i50/n527 ;
 wire \i50/n528 ;
 wire \i50/n529 ;
 wire \i50/n53 ;
 wire \i50/n530 ;
 wire \i50/n531 ;
 wire \i50/n532 ;
 wire \i50/n533 ;
 wire \i50/n534 ;
 wire \i50/n535 ;
 wire \i50/n536 ;
 wire \i50/n537 ;
 wire \i50/n538 ;
 wire \i50/n539 ;
 wire \i50/n54 ;
 wire \i50/n540 ;
 wire \i50/n541 ;
 wire \i50/n542 ;
 wire \i50/n543 ;
 wire \i50/n544 ;
 wire \i50/n545 ;
 wire \i50/n546 ;
 wire \i50/n547 ;
 wire \i50/n548 ;
 wire \i50/n549 ;
 wire \i50/n55 ;
 wire \i50/n550 ;
 wire \i50/n551 ;
 wire \i50/n552 ;
 wire \i50/n553 ;
 wire \i50/n554 ;
 wire \i50/n555 ;
 wire \i50/n556 ;
 wire \i50/n557 ;
 wire \i50/n558 ;
 wire \i50/n559 ;
 wire \i50/n56 ;
 wire \i50/n560 ;
 wire \i50/n561 ;
 wire \i50/n562 ;
 wire \i50/n563 ;
 wire \i50/n564 ;
 wire \i50/n565 ;
 wire \i50/n566 ;
 wire \i50/n567 ;
 wire \i50/n568 ;
 wire \i50/n569 ;
 wire \i50/n57 ;
 wire \i50/n570 ;
 wire \i50/n571 ;
 wire \i50/n572 ;
 wire \i50/n573 ;
 wire \i50/n574 ;
 wire \i50/n575 ;
 wire \i50/n576 ;
 wire \i50/n577 ;
 wire \i50/n578 ;
 wire \i50/n579 ;
 wire \i50/n58 ;
 wire \i50/n580 ;
 wire \i50/n59 ;
 wire \i50/n6 ;
 wire \i50/n60 ;
 wire \i50/n61 ;
 wire \i50/n62 ;
 wire \i50/n63 ;
 wire \i50/n64 ;
 wire \i50/n65 ;
 wire \i50/n66 ;
 wire \i50/n67 ;
 wire \i50/n68 ;
 wire \i50/n69 ;
 wire \i50/n7 ;
 wire \i50/n70 ;
 wire \i50/n71 ;
 wire \i50/n72 ;
 wire \i50/n73 ;
 wire \i50/n74 ;
 wire \i50/n75 ;
 wire \i50/n76 ;
 wire \i50/n77 ;
 wire \i50/n78 ;
 wire \i50/n79 ;
 wire \i50/n8 ;
 wire \i50/n80 ;
 wire \i50/n81 ;
 wire \i50/n82 ;
 wire \i50/n83 ;
 wire \i50/n84 ;
 wire \i50/n85 ;
 wire \i50/n86 ;
 wire \i50/n87 ;
 wire \i50/n88 ;
 wire \i50/n89 ;
 wire \i50/n9 ;
 wire \i50/n90 ;
 wire \i50/n91 ;
 wire \i50/n92 ;
 wire \i50/n93 ;
 wire \i50/n94 ;
 wire \i50/n95 ;
 wire \i50/n96 ;
 wire \i50/n97 ;
 wire \i50/n98 ;
 wire \i50/n99 ;
 wire \i51/n0 ;
 wire \i51/n1 ;
 wire \i51/n10 ;
 wire \i51/n100 ;
 wire \i51/n101 ;
 wire \i51/n102 ;
 wire \i51/n103 ;
 wire \i51/n104 ;
 wire \i51/n105 ;
 wire \i51/n106 ;
 wire \i51/n107 ;
 wire \i51/n108 ;
 wire \i51/n109 ;
 wire \i51/n11 ;
 wire \i51/n110 ;
 wire \i51/n111 ;
 wire \i51/n112 ;
 wire \i51/n113 ;
 wire \i51/n114 ;
 wire \i51/n115 ;
 wire \i51/n116 ;
 wire \i51/n117 ;
 wire \i51/n118 ;
 wire \i51/n119 ;
 wire \i51/n12 ;
 wire \i51/n120 ;
 wire \i51/n121 ;
 wire \i51/n122 ;
 wire \i51/n123 ;
 wire \i51/n124 ;
 wire \i51/n125 ;
 wire \i51/n126 ;
 wire \i51/n127 ;
 wire \i51/n128 ;
 wire \i51/n129 ;
 wire \i51/n13 ;
 wire \i51/n130 ;
 wire \i51/n131 ;
 wire \i51/n132 ;
 wire \i51/n133 ;
 wire \i51/n134 ;
 wire \i51/n135 ;
 wire \i51/n136 ;
 wire \i51/n137 ;
 wire \i51/n138 ;
 wire \i51/n139 ;
 wire \i51/n14 ;
 wire \i51/n140 ;
 wire \i51/n141 ;
 wire \i51/n142 ;
 wire \i51/n143 ;
 wire \i51/n144 ;
 wire \i51/n145 ;
 wire \i51/n146 ;
 wire \i51/n147 ;
 wire \i51/n148 ;
 wire \i51/n149 ;
 wire \i51/n15 ;
 wire \i51/n150 ;
 wire \i51/n151 ;
 wire \i51/n152 ;
 wire \i51/n153 ;
 wire \i51/n154 ;
 wire \i51/n155 ;
 wire \i51/n156 ;
 wire \i51/n157 ;
 wire \i51/n158 ;
 wire \i51/n159 ;
 wire \i51/n16 ;
 wire \i51/n160 ;
 wire \i51/n161 ;
 wire \i51/n162 ;
 wire \i51/n163 ;
 wire \i51/n164 ;
 wire \i51/n165 ;
 wire \i51/n166 ;
 wire \i51/n167 ;
 wire \i51/n168 ;
 wire \i51/n169 ;
 wire \i51/n17 ;
 wire \i51/n170 ;
 wire \i51/n171 ;
 wire \i51/n172 ;
 wire \i51/n173 ;
 wire \i51/n174 ;
 wire \i51/n175 ;
 wire \i51/n176 ;
 wire \i51/n177 ;
 wire \i51/n178 ;
 wire \i51/n179 ;
 wire \i51/n18 ;
 wire \i51/n180 ;
 wire \i51/n181 ;
 wire \i51/n182 ;
 wire \i51/n183 ;
 wire \i51/n184 ;
 wire \i51/n185 ;
 wire \i51/n186 ;
 wire \i51/n187 ;
 wire \i51/n188 ;
 wire \i51/n189 ;
 wire \i51/n19 ;
 wire \i51/n190 ;
 wire \i51/n191 ;
 wire \i51/n192 ;
 wire \i51/n193 ;
 wire \i51/n194 ;
 wire \i51/n195 ;
 wire \i51/n196 ;
 wire \i51/n197 ;
 wire \i51/n198 ;
 wire \i51/n199 ;
 wire \i51/n2 ;
 wire \i51/n20 ;
 wire \i51/n200 ;
 wire \i51/n201 ;
 wire \i51/n202 ;
 wire \i51/n203 ;
 wire \i51/n204 ;
 wire \i51/n205 ;
 wire \i51/n206 ;
 wire \i51/n207 ;
 wire \i51/n208 ;
 wire \i51/n209 ;
 wire \i51/n21 ;
 wire \i51/n210 ;
 wire \i51/n211 ;
 wire \i51/n212 ;
 wire \i51/n213 ;
 wire \i51/n214 ;
 wire \i51/n215 ;
 wire \i51/n216 ;
 wire \i51/n217 ;
 wire \i51/n218 ;
 wire \i51/n219 ;
 wire \i51/n22 ;
 wire \i51/n220 ;
 wire \i51/n221 ;
 wire \i51/n222 ;
 wire \i51/n223 ;
 wire \i51/n224 ;
 wire \i51/n225 ;
 wire \i51/n226 ;
 wire \i51/n227 ;
 wire \i51/n228 ;
 wire \i51/n229 ;
 wire \i51/n23 ;
 wire \i51/n230 ;
 wire \i51/n231 ;
 wire \i51/n232 ;
 wire \i51/n233 ;
 wire \i51/n234 ;
 wire \i51/n235 ;
 wire \i51/n236 ;
 wire \i51/n237 ;
 wire \i51/n238 ;
 wire \i51/n239 ;
 wire \i51/n24 ;
 wire \i51/n240 ;
 wire \i51/n241 ;
 wire \i51/n242 ;
 wire \i51/n243 ;
 wire \i51/n244 ;
 wire \i51/n245 ;
 wire \i51/n246 ;
 wire \i51/n247 ;
 wire \i51/n248 ;
 wire \i51/n249 ;
 wire \i51/n25 ;
 wire \i51/n250 ;
 wire \i51/n251 ;
 wire \i51/n252 ;
 wire \i51/n253 ;
 wire \i51/n254 ;
 wire \i51/n255 ;
 wire \i51/n256 ;
 wire \i51/n257 ;
 wire \i51/n258 ;
 wire \i51/n259 ;
 wire \i51/n26 ;
 wire \i51/n260 ;
 wire \i51/n261 ;
 wire \i51/n262 ;
 wire \i51/n263 ;
 wire \i51/n264 ;
 wire \i51/n265 ;
 wire \i51/n266 ;
 wire \i51/n267 ;
 wire \i51/n268 ;
 wire \i51/n269 ;
 wire \i51/n27 ;
 wire \i51/n270 ;
 wire \i51/n271 ;
 wire \i51/n272 ;
 wire \i51/n273 ;
 wire \i51/n274 ;
 wire \i51/n275 ;
 wire \i51/n276 ;
 wire \i51/n277 ;
 wire \i51/n278 ;
 wire \i51/n279 ;
 wire \i51/n28 ;
 wire \i51/n280 ;
 wire \i51/n281 ;
 wire \i51/n282 ;
 wire \i51/n283 ;
 wire \i51/n284 ;
 wire \i51/n285 ;
 wire \i51/n286 ;
 wire \i51/n287 ;
 wire \i51/n288 ;
 wire \i51/n289 ;
 wire \i51/n29 ;
 wire \i51/n290 ;
 wire \i51/n291 ;
 wire \i51/n292 ;
 wire \i51/n293 ;
 wire \i51/n294 ;
 wire \i51/n295 ;
 wire \i51/n296 ;
 wire \i51/n297 ;
 wire \i51/n298 ;
 wire \i51/n299 ;
 wire \i51/n3 ;
 wire \i51/n30 ;
 wire \i51/n300 ;
 wire \i51/n301 ;
 wire \i51/n302 ;
 wire \i51/n303 ;
 wire \i51/n304 ;
 wire \i51/n305 ;
 wire \i51/n306 ;
 wire \i51/n307 ;
 wire \i51/n308 ;
 wire \i51/n309 ;
 wire \i51/n31 ;
 wire \i51/n310 ;
 wire \i51/n311 ;
 wire \i51/n312 ;
 wire \i51/n313 ;
 wire \i51/n314 ;
 wire \i51/n315 ;
 wire \i51/n316 ;
 wire \i51/n317 ;
 wire \i51/n318 ;
 wire \i51/n319 ;
 wire \i51/n32 ;
 wire \i51/n320 ;
 wire \i51/n321 ;
 wire \i51/n322 ;
 wire \i51/n323 ;
 wire \i51/n324 ;
 wire \i51/n325 ;
 wire \i51/n326 ;
 wire \i51/n327 ;
 wire \i51/n328 ;
 wire \i51/n329 ;
 wire \i51/n33 ;
 wire \i51/n330 ;
 wire \i51/n331 ;
 wire \i51/n332 ;
 wire \i51/n333 ;
 wire \i51/n334 ;
 wire \i51/n335 ;
 wire \i51/n336 ;
 wire \i51/n337 ;
 wire \i51/n338 ;
 wire \i51/n339 ;
 wire \i51/n34 ;
 wire \i51/n340 ;
 wire \i51/n341 ;
 wire \i51/n342 ;
 wire \i51/n343 ;
 wire \i51/n344 ;
 wire \i51/n345 ;
 wire \i51/n346 ;
 wire \i51/n347 ;
 wire \i51/n348 ;
 wire \i51/n349 ;
 wire \i51/n35 ;
 wire \i51/n350 ;
 wire \i51/n351 ;
 wire \i51/n352 ;
 wire \i51/n353 ;
 wire \i51/n354 ;
 wire \i51/n355 ;
 wire \i51/n356 ;
 wire \i51/n357 ;
 wire \i51/n358 ;
 wire \i51/n359 ;
 wire \i51/n36 ;
 wire \i51/n360 ;
 wire \i51/n361 ;
 wire \i51/n362 ;
 wire \i51/n363 ;
 wire \i51/n364 ;
 wire \i51/n365 ;
 wire \i51/n366 ;
 wire \i51/n367 ;
 wire \i51/n368 ;
 wire \i51/n369 ;
 wire \i51/n37 ;
 wire \i51/n370 ;
 wire \i51/n371 ;
 wire \i51/n372 ;
 wire \i51/n373 ;
 wire \i51/n374 ;
 wire \i51/n375 ;
 wire \i51/n376 ;
 wire \i51/n377 ;
 wire \i51/n378 ;
 wire \i51/n379 ;
 wire \i51/n38 ;
 wire \i51/n380 ;
 wire \i51/n381 ;
 wire \i51/n382 ;
 wire \i51/n383 ;
 wire \i51/n384 ;
 wire \i51/n385 ;
 wire \i51/n386 ;
 wire \i51/n387 ;
 wire \i51/n388 ;
 wire \i51/n389 ;
 wire \i51/n39 ;
 wire \i51/n390 ;
 wire \i51/n391 ;
 wire \i51/n392 ;
 wire \i51/n393 ;
 wire \i51/n394 ;
 wire \i51/n395 ;
 wire \i51/n396 ;
 wire \i51/n397 ;
 wire \i51/n398 ;
 wire \i51/n399 ;
 wire \i51/n4 ;
 wire \i51/n40 ;
 wire \i51/n400 ;
 wire \i51/n401 ;
 wire \i51/n402 ;
 wire \i51/n403 ;
 wire \i51/n404 ;
 wire \i51/n405 ;
 wire \i51/n406 ;
 wire \i51/n407 ;
 wire \i51/n408 ;
 wire \i51/n409 ;
 wire \i51/n41 ;
 wire \i51/n410 ;
 wire \i51/n411 ;
 wire \i51/n412 ;
 wire \i51/n413 ;
 wire \i51/n414 ;
 wire \i51/n415 ;
 wire \i51/n416 ;
 wire \i51/n417 ;
 wire \i51/n418 ;
 wire \i51/n419 ;
 wire \i51/n42 ;
 wire \i51/n420 ;
 wire \i51/n421 ;
 wire \i51/n422 ;
 wire \i51/n423 ;
 wire \i51/n424 ;
 wire \i51/n425 ;
 wire \i51/n426 ;
 wire \i51/n427 ;
 wire \i51/n428 ;
 wire \i51/n429 ;
 wire \i51/n43 ;
 wire \i51/n430 ;
 wire \i51/n431 ;
 wire \i51/n432 ;
 wire \i51/n433 ;
 wire \i51/n434 ;
 wire \i51/n435 ;
 wire \i51/n436 ;
 wire \i51/n437 ;
 wire \i51/n438 ;
 wire \i51/n439 ;
 wire \i51/n44 ;
 wire \i51/n440 ;
 wire \i51/n441 ;
 wire \i51/n442 ;
 wire \i51/n443 ;
 wire \i51/n444 ;
 wire \i51/n445 ;
 wire \i51/n446 ;
 wire \i51/n447 ;
 wire \i51/n448 ;
 wire \i51/n449 ;
 wire \i51/n45 ;
 wire \i51/n450 ;
 wire \i51/n451 ;
 wire \i51/n452 ;
 wire \i51/n453 ;
 wire \i51/n454 ;
 wire \i51/n455 ;
 wire \i51/n456 ;
 wire \i51/n457 ;
 wire \i51/n458 ;
 wire \i51/n459 ;
 wire \i51/n46 ;
 wire \i51/n460 ;
 wire \i51/n461 ;
 wire \i51/n462 ;
 wire \i51/n463 ;
 wire \i51/n464 ;
 wire \i51/n465 ;
 wire \i51/n466 ;
 wire \i51/n467 ;
 wire \i51/n468 ;
 wire \i51/n469 ;
 wire \i51/n47 ;
 wire \i51/n470 ;
 wire \i51/n471 ;
 wire \i51/n472 ;
 wire \i51/n473 ;
 wire \i51/n474 ;
 wire \i51/n475 ;
 wire \i51/n476 ;
 wire \i51/n477 ;
 wire \i51/n478 ;
 wire \i51/n479 ;
 wire \i51/n48 ;
 wire \i51/n480 ;
 wire \i51/n481 ;
 wire \i51/n482 ;
 wire \i51/n483 ;
 wire \i51/n484 ;
 wire \i51/n485 ;
 wire \i51/n486 ;
 wire \i51/n487 ;
 wire \i51/n488 ;
 wire \i51/n489 ;
 wire \i51/n49 ;
 wire \i51/n490 ;
 wire \i51/n491 ;
 wire \i51/n492 ;
 wire \i51/n493 ;
 wire \i51/n494 ;
 wire \i51/n495 ;
 wire \i51/n496 ;
 wire \i51/n497 ;
 wire \i51/n498 ;
 wire \i51/n499 ;
 wire \i51/n5 ;
 wire \i51/n50 ;
 wire \i51/n500 ;
 wire \i51/n501 ;
 wire \i51/n502 ;
 wire \i51/n503 ;
 wire \i51/n504 ;
 wire \i51/n505 ;
 wire \i51/n506 ;
 wire \i51/n507 ;
 wire \i51/n508 ;
 wire \i51/n509 ;
 wire \i51/n51 ;
 wire \i51/n510 ;
 wire \i51/n511 ;
 wire \i51/n512 ;
 wire \i51/n513 ;
 wire \i51/n514 ;
 wire \i51/n515 ;
 wire \i51/n516 ;
 wire \i51/n517 ;
 wire \i51/n518 ;
 wire \i51/n519 ;
 wire \i51/n52 ;
 wire \i51/n520 ;
 wire \i51/n521 ;
 wire \i51/n522 ;
 wire \i51/n523 ;
 wire \i51/n524 ;
 wire \i51/n525 ;
 wire \i51/n526 ;
 wire \i51/n527 ;
 wire \i51/n528 ;
 wire \i51/n529 ;
 wire \i51/n53 ;
 wire \i51/n530 ;
 wire \i51/n531 ;
 wire \i51/n532 ;
 wire \i51/n533 ;
 wire \i51/n534 ;
 wire \i51/n535 ;
 wire \i51/n536 ;
 wire \i51/n537 ;
 wire \i51/n538 ;
 wire \i51/n539 ;
 wire \i51/n54 ;
 wire \i51/n540 ;
 wire \i51/n541 ;
 wire \i51/n542 ;
 wire \i51/n543 ;
 wire \i51/n544 ;
 wire \i51/n545 ;
 wire \i51/n546 ;
 wire \i51/n547 ;
 wire \i51/n548 ;
 wire \i51/n549 ;
 wire \i51/n55 ;
 wire \i51/n550 ;
 wire \i51/n551 ;
 wire \i51/n552 ;
 wire \i51/n553 ;
 wire \i51/n554 ;
 wire \i51/n555 ;
 wire \i51/n556 ;
 wire \i51/n557 ;
 wire \i51/n558 ;
 wire \i51/n559 ;
 wire \i51/n56 ;
 wire \i51/n560 ;
 wire \i51/n561 ;
 wire \i51/n562 ;
 wire \i51/n563 ;
 wire \i51/n564 ;
 wire \i51/n565 ;
 wire \i51/n566 ;
 wire \i51/n567 ;
 wire \i51/n568 ;
 wire \i51/n569 ;
 wire \i51/n57 ;
 wire \i51/n570 ;
 wire \i51/n571 ;
 wire \i51/n572 ;
 wire \i51/n573 ;
 wire \i51/n574 ;
 wire \i51/n575 ;
 wire \i51/n576 ;
 wire \i51/n577 ;
 wire \i51/n578 ;
 wire \i51/n579 ;
 wire \i51/n58 ;
 wire \i51/n580 ;
 wire \i51/n581 ;
 wire \i51/n582 ;
 wire \i51/n583 ;
 wire \i51/n59 ;
 wire \i51/n6 ;
 wire \i51/n60 ;
 wire \i51/n61 ;
 wire \i51/n62 ;
 wire \i51/n63 ;
 wire \i51/n64 ;
 wire \i51/n65 ;
 wire \i51/n66 ;
 wire \i51/n67 ;
 wire \i51/n68 ;
 wire \i51/n69 ;
 wire \i51/n7 ;
 wire \i51/n70 ;
 wire \i51/n71 ;
 wire \i51/n72 ;
 wire \i51/n73 ;
 wire \i51/n74 ;
 wire \i51/n75 ;
 wire \i51/n76 ;
 wire \i51/n77 ;
 wire \i51/n78 ;
 wire \i51/n79 ;
 wire \i51/n8 ;
 wire \i51/n80 ;
 wire \i51/n81 ;
 wire \i51/n82 ;
 wire \i51/n83 ;
 wire \i51/n84 ;
 wire \i51/n85 ;
 wire \i51/n86 ;
 wire \i51/n87 ;
 wire \i51/n88 ;
 wire \i51/n89 ;
 wire \i51/n9 ;
 wire \i51/n90 ;
 wire \i51/n91 ;
 wire \i51/n92 ;
 wire \i51/n93 ;
 wire \i51/n94 ;
 wire \i51/n95 ;
 wire \i51/n96 ;
 wire \i51/n97 ;
 wire \i51/n98 ;
 wire \i51/n99 ;
 wire \i52/n0 ;
 wire \i52/n1 ;
 wire \i52/n10 ;
 wire \i52/n100 ;
 wire \i52/n101 ;
 wire \i52/n102 ;
 wire \i52/n103 ;
 wire \i52/n104 ;
 wire \i52/n105 ;
 wire \i52/n106 ;
 wire \i52/n107 ;
 wire \i52/n108 ;
 wire \i52/n109 ;
 wire \i52/n11 ;
 wire \i52/n110 ;
 wire \i52/n111 ;
 wire \i52/n112 ;
 wire \i52/n113 ;
 wire \i52/n114 ;
 wire \i52/n115 ;
 wire \i52/n116 ;
 wire \i52/n117 ;
 wire \i52/n118 ;
 wire \i52/n119 ;
 wire \i52/n12 ;
 wire \i52/n120 ;
 wire \i52/n121 ;
 wire \i52/n122 ;
 wire \i52/n123 ;
 wire \i52/n124 ;
 wire \i52/n125 ;
 wire \i52/n126 ;
 wire \i52/n127 ;
 wire \i52/n128 ;
 wire \i52/n129 ;
 wire \i52/n13 ;
 wire \i52/n130 ;
 wire \i52/n131 ;
 wire \i52/n132 ;
 wire \i52/n133 ;
 wire \i52/n134 ;
 wire \i52/n135 ;
 wire \i52/n136 ;
 wire \i52/n137 ;
 wire \i52/n138 ;
 wire \i52/n139 ;
 wire \i52/n14 ;
 wire \i52/n140 ;
 wire \i52/n141 ;
 wire \i52/n142 ;
 wire \i52/n143 ;
 wire \i52/n144 ;
 wire \i52/n145 ;
 wire \i52/n146 ;
 wire \i52/n147 ;
 wire \i52/n148 ;
 wire \i52/n149 ;
 wire \i52/n15 ;
 wire \i52/n150 ;
 wire \i52/n151 ;
 wire \i52/n152 ;
 wire \i52/n153 ;
 wire \i52/n154 ;
 wire \i52/n155 ;
 wire \i52/n156 ;
 wire \i52/n157 ;
 wire \i52/n158 ;
 wire \i52/n159 ;
 wire \i52/n16 ;
 wire \i52/n160 ;
 wire \i52/n161 ;
 wire \i52/n162 ;
 wire \i52/n163 ;
 wire \i52/n164 ;
 wire \i52/n165 ;
 wire \i52/n166 ;
 wire \i52/n167 ;
 wire \i52/n168 ;
 wire \i52/n169 ;
 wire \i52/n17 ;
 wire \i52/n170 ;
 wire \i52/n171 ;
 wire \i52/n172 ;
 wire \i52/n173 ;
 wire \i52/n174 ;
 wire \i52/n175 ;
 wire \i52/n176 ;
 wire \i52/n177 ;
 wire \i52/n178 ;
 wire \i52/n179 ;
 wire \i52/n18 ;
 wire \i52/n180 ;
 wire \i52/n181 ;
 wire \i52/n182 ;
 wire \i52/n183 ;
 wire \i52/n184 ;
 wire \i52/n185 ;
 wire \i52/n186 ;
 wire \i52/n187 ;
 wire \i52/n188 ;
 wire \i52/n189 ;
 wire \i52/n19 ;
 wire \i52/n190 ;
 wire \i52/n191 ;
 wire \i52/n192 ;
 wire \i52/n193 ;
 wire \i52/n194 ;
 wire \i52/n195 ;
 wire \i52/n196 ;
 wire \i52/n197 ;
 wire \i52/n198 ;
 wire \i52/n199 ;
 wire \i52/n2 ;
 wire \i52/n20 ;
 wire \i52/n200 ;
 wire \i52/n201 ;
 wire \i52/n202 ;
 wire \i52/n203 ;
 wire \i52/n204 ;
 wire \i52/n205 ;
 wire \i52/n206 ;
 wire \i52/n207 ;
 wire \i52/n208 ;
 wire \i52/n209 ;
 wire \i52/n21 ;
 wire \i52/n210 ;
 wire \i52/n211 ;
 wire \i52/n212 ;
 wire \i52/n213 ;
 wire \i52/n214 ;
 wire \i52/n215 ;
 wire \i52/n216 ;
 wire \i52/n217 ;
 wire \i52/n218 ;
 wire \i52/n219 ;
 wire \i52/n22 ;
 wire \i52/n220 ;
 wire \i52/n221 ;
 wire \i52/n222 ;
 wire \i52/n223 ;
 wire \i52/n224 ;
 wire \i52/n225 ;
 wire \i52/n226 ;
 wire \i52/n227 ;
 wire \i52/n228 ;
 wire \i52/n229 ;
 wire \i52/n23 ;
 wire \i52/n230 ;
 wire \i52/n231 ;
 wire \i52/n232 ;
 wire \i52/n233 ;
 wire \i52/n234 ;
 wire \i52/n235 ;
 wire \i52/n236 ;
 wire \i52/n237 ;
 wire \i52/n238 ;
 wire \i52/n239 ;
 wire \i52/n24 ;
 wire \i52/n240 ;
 wire \i52/n241 ;
 wire \i52/n242 ;
 wire \i52/n243 ;
 wire \i52/n244 ;
 wire \i52/n245 ;
 wire \i52/n246 ;
 wire \i52/n247 ;
 wire \i52/n248 ;
 wire \i52/n249 ;
 wire \i52/n25 ;
 wire \i52/n250 ;
 wire \i52/n251 ;
 wire \i52/n252 ;
 wire \i52/n253 ;
 wire \i52/n254 ;
 wire \i52/n255 ;
 wire \i52/n256 ;
 wire \i52/n257 ;
 wire \i52/n258 ;
 wire \i52/n259 ;
 wire \i52/n26 ;
 wire \i52/n260 ;
 wire \i52/n261 ;
 wire \i52/n262 ;
 wire \i52/n263 ;
 wire \i52/n264 ;
 wire \i52/n265 ;
 wire \i52/n266 ;
 wire \i52/n267 ;
 wire \i52/n268 ;
 wire \i52/n269 ;
 wire \i52/n27 ;
 wire \i52/n270 ;
 wire \i52/n271 ;
 wire \i52/n272 ;
 wire \i52/n273 ;
 wire \i52/n274 ;
 wire \i52/n275 ;
 wire \i52/n276 ;
 wire \i52/n277 ;
 wire \i52/n278 ;
 wire \i52/n279 ;
 wire \i52/n28 ;
 wire \i52/n280 ;
 wire \i52/n281 ;
 wire \i52/n282 ;
 wire \i52/n283 ;
 wire \i52/n284 ;
 wire \i52/n285 ;
 wire \i52/n286 ;
 wire \i52/n287 ;
 wire \i52/n288 ;
 wire \i52/n289 ;
 wire \i52/n29 ;
 wire \i52/n290 ;
 wire \i52/n291 ;
 wire \i52/n292 ;
 wire \i52/n293 ;
 wire \i52/n294 ;
 wire \i52/n295 ;
 wire \i52/n296 ;
 wire \i52/n297 ;
 wire \i52/n298 ;
 wire \i52/n299 ;
 wire \i52/n3 ;
 wire \i52/n30 ;
 wire \i52/n300 ;
 wire \i52/n301 ;
 wire \i52/n302 ;
 wire \i52/n303 ;
 wire \i52/n304 ;
 wire \i52/n305 ;
 wire \i52/n306 ;
 wire \i52/n307 ;
 wire \i52/n308 ;
 wire \i52/n309 ;
 wire \i52/n31 ;
 wire \i52/n310 ;
 wire \i52/n311 ;
 wire \i52/n312 ;
 wire \i52/n313 ;
 wire \i52/n314 ;
 wire \i52/n315 ;
 wire \i52/n316 ;
 wire \i52/n317 ;
 wire \i52/n318 ;
 wire \i52/n319 ;
 wire \i52/n32 ;
 wire \i52/n320 ;
 wire \i52/n321 ;
 wire \i52/n322 ;
 wire \i52/n323 ;
 wire \i52/n324 ;
 wire \i52/n325 ;
 wire \i52/n326 ;
 wire \i52/n327 ;
 wire \i52/n328 ;
 wire \i52/n329 ;
 wire \i52/n33 ;
 wire \i52/n330 ;
 wire \i52/n331 ;
 wire \i52/n332 ;
 wire \i52/n333 ;
 wire \i52/n334 ;
 wire \i52/n335 ;
 wire \i52/n336 ;
 wire \i52/n337 ;
 wire \i52/n338 ;
 wire \i52/n339 ;
 wire \i52/n34 ;
 wire \i52/n340 ;
 wire \i52/n341 ;
 wire \i52/n342 ;
 wire \i52/n343 ;
 wire \i52/n344 ;
 wire \i52/n345 ;
 wire \i52/n346 ;
 wire \i52/n347 ;
 wire \i52/n348 ;
 wire \i52/n349 ;
 wire \i52/n35 ;
 wire \i52/n350 ;
 wire \i52/n351 ;
 wire \i52/n352 ;
 wire \i52/n353 ;
 wire \i52/n354 ;
 wire \i52/n355 ;
 wire \i52/n356 ;
 wire \i52/n357 ;
 wire \i52/n358 ;
 wire \i52/n359 ;
 wire \i52/n36 ;
 wire \i52/n360 ;
 wire \i52/n361 ;
 wire \i52/n362 ;
 wire \i52/n363 ;
 wire \i52/n364 ;
 wire \i52/n365 ;
 wire \i52/n366 ;
 wire \i52/n367 ;
 wire \i52/n368 ;
 wire \i52/n369 ;
 wire \i52/n37 ;
 wire \i52/n370 ;
 wire \i52/n371 ;
 wire \i52/n372 ;
 wire \i52/n373 ;
 wire \i52/n374 ;
 wire \i52/n375 ;
 wire \i52/n376 ;
 wire \i52/n377 ;
 wire \i52/n378 ;
 wire \i52/n379 ;
 wire \i52/n38 ;
 wire \i52/n380 ;
 wire \i52/n381 ;
 wire \i52/n382 ;
 wire \i52/n383 ;
 wire \i52/n384 ;
 wire \i52/n385 ;
 wire \i52/n386 ;
 wire \i52/n387 ;
 wire \i52/n388 ;
 wire \i52/n389 ;
 wire \i52/n39 ;
 wire \i52/n390 ;
 wire \i52/n391 ;
 wire \i52/n392 ;
 wire \i52/n393 ;
 wire \i52/n394 ;
 wire \i52/n395 ;
 wire \i52/n396 ;
 wire \i52/n397 ;
 wire \i52/n398 ;
 wire \i52/n399 ;
 wire \i52/n4 ;
 wire \i52/n40 ;
 wire \i52/n400 ;
 wire \i52/n401 ;
 wire \i52/n402 ;
 wire \i52/n403 ;
 wire \i52/n404 ;
 wire \i52/n405 ;
 wire \i52/n406 ;
 wire \i52/n407 ;
 wire \i52/n408 ;
 wire \i52/n409 ;
 wire \i52/n41 ;
 wire \i52/n410 ;
 wire \i52/n411 ;
 wire \i52/n412 ;
 wire \i52/n413 ;
 wire \i52/n414 ;
 wire \i52/n415 ;
 wire \i52/n416 ;
 wire \i52/n417 ;
 wire \i52/n418 ;
 wire \i52/n419 ;
 wire \i52/n42 ;
 wire \i52/n420 ;
 wire \i52/n421 ;
 wire \i52/n422 ;
 wire \i52/n423 ;
 wire \i52/n424 ;
 wire \i52/n425 ;
 wire \i52/n426 ;
 wire \i52/n427 ;
 wire \i52/n428 ;
 wire \i52/n429 ;
 wire \i52/n43 ;
 wire \i52/n430 ;
 wire \i52/n431 ;
 wire \i52/n432 ;
 wire \i52/n433 ;
 wire \i52/n434 ;
 wire \i52/n435 ;
 wire \i52/n436 ;
 wire \i52/n437 ;
 wire \i52/n438 ;
 wire \i52/n439 ;
 wire \i52/n44 ;
 wire \i52/n440 ;
 wire \i52/n441 ;
 wire \i52/n442 ;
 wire \i52/n443 ;
 wire \i52/n444 ;
 wire \i52/n445 ;
 wire \i52/n446 ;
 wire \i52/n447 ;
 wire \i52/n448 ;
 wire \i52/n449 ;
 wire \i52/n45 ;
 wire \i52/n450 ;
 wire \i52/n451 ;
 wire \i52/n452 ;
 wire \i52/n453 ;
 wire \i52/n454 ;
 wire \i52/n455 ;
 wire \i52/n456 ;
 wire \i52/n457 ;
 wire \i52/n458 ;
 wire \i52/n459 ;
 wire \i52/n46 ;
 wire \i52/n460 ;
 wire \i52/n461 ;
 wire \i52/n462 ;
 wire \i52/n463 ;
 wire \i52/n464 ;
 wire \i52/n465 ;
 wire \i52/n466 ;
 wire \i52/n467 ;
 wire \i52/n468 ;
 wire \i52/n469 ;
 wire \i52/n47 ;
 wire \i52/n470 ;
 wire \i52/n471 ;
 wire \i52/n472 ;
 wire \i52/n473 ;
 wire \i52/n474 ;
 wire \i52/n475 ;
 wire \i52/n476 ;
 wire \i52/n477 ;
 wire \i52/n478 ;
 wire \i52/n479 ;
 wire \i52/n48 ;
 wire \i52/n480 ;
 wire \i52/n481 ;
 wire \i52/n482 ;
 wire \i52/n483 ;
 wire \i52/n484 ;
 wire \i52/n485 ;
 wire \i52/n486 ;
 wire \i52/n487 ;
 wire \i52/n488 ;
 wire \i52/n489 ;
 wire \i52/n49 ;
 wire \i52/n490 ;
 wire \i52/n491 ;
 wire \i52/n492 ;
 wire \i52/n493 ;
 wire \i52/n494 ;
 wire \i52/n495 ;
 wire \i52/n496 ;
 wire \i52/n497 ;
 wire \i52/n498 ;
 wire \i52/n499 ;
 wire \i52/n5 ;
 wire \i52/n50 ;
 wire \i52/n500 ;
 wire \i52/n501 ;
 wire \i52/n502 ;
 wire \i52/n503 ;
 wire \i52/n504 ;
 wire \i52/n505 ;
 wire \i52/n506 ;
 wire \i52/n507 ;
 wire \i52/n508 ;
 wire \i52/n509 ;
 wire \i52/n51 ;
 wire \i52/n510 ;
 wire \i52/n511 ;
 wire \i52/n512 ;
 wire \i52/n513 ;
 wire \i52/n514 ;
 wire \i52/n515 ;
 wire \i52/n516 ;
 wire \i52/n517 ;
 wire \i52/n518 ;
 wire \i52/n519 ;
 wire \i52/n52 ;
 wire \i52/n520 ;
 wire \i52/n521 ;
 wire \i52/n522 ;
 wire \i52/n523 ;
 wire \i52/n524 ;
 wire \i52/n525 ;
 wire \i52/n526 ;
 wire \i52/n527 ;
 wire \i52/n528 ;
 wire \i52/n529 ;
 wire \i52/n53 ;
 wire \i52/n530 ;
 wire \i52/n531 ;
 wire \i52/n532 ;
 wire \i52/n533 ;
 wire \i52/n534 ;
 wire \i52/n535 ;
 wire \i52/n536 ;
 wire \i52/n537 ;
 wire \i52/n538 ;
 wire \i52/n539 ;
 wire \i52/n54 ;
 wire \i52/n540 ;
 wire \i52/n541 ;
 wire \i52/n542 ;
 wire \i52/n543 ;
 wire \i52/n544 ;
 wire \i52/n545 ;
 wire \i52/n546 ;
 wire \i52/n547 ;
 wire \i52/n548 ;
 wire \i52/n549 ;
 wire \i52/n55 ;
 wire \i52/n550 ;
 wire \i52/n551 ;
 wire \i52/n552 ;
 wire \i52/n553 ;
 wire \i52/n554 ;
 wire \i52/n555 ;
 wire \i52/n556 ;
 wire \i52/n557 ;
 wire \i52/n558 ;
 wire \i52/n559 ;
 wire \i52/n56 ;
 wire \i52/n560 ;
 wire \i52/n561 ;
 wire \i52/n562 ;
 wire \i52/n563 ;
 wire \i52/n564 ;
 wire \i52/n565 ;
 wire \i52/n566 ;
 wire \i52/n567 ;
 wire \i52/n568 ;
 wire \i52/n569 ;
 wire \i52/n57 ;
 wire \i52/n570 ;
 wire \i52/n571 ;
 wire \i52/n572 ;
 wire \i52/n573 ;
 wire \i52/n574 ;
 wire \i52/n575 ;
 wire \i52/n576 ;
 wire \i52/n577 ;
 wire \i52/n578 ;
 wire \i52/n579 ;
 wire \i52/n58 ;
 wire \i52/n580 ;
 wire \i52/n581 ;
 wire \i52/n59 ;
 wire \i52/n6 ;
 wire \i52/n60 ;
 wire \i52/n61 ;
 wire \i52/n62 ;
 wire \i52/n63 ;
 wire \i52/n64 ;
 wire \i52/n65 ;
 wire \i52/n66 ;
 wire \i52/n67 ;
 wire \i52/n68 ;
 wire \i52/n69 ;
 wire \i52/n7 ;
 wire \i52/n70 ;
 wire \i52/n71 ;
 wire \i52/n72 ;
 wire \i52/n73 ;
 wire \i52/n74 ;
 wire \i52/n75 ;
 wire \i52/n76 ;
 wire \i52/n77 ;
 wire \i52/n78 ;
 wire \i52/n79 ;
 wire \i52/n8 ;
 wire \i52/n80 ;
 wire \i52/n81 ;
 wire \i52/n82 ;
 wire \i52/n83 ;
 wire \i52/n84 ;
 wire \i52/n85 ;
 wire \i52/n86 ;
 wire \i52/n87 ;
 wire \i52/n88 ;
 wire \i52/n89 ;
 wire \i52/n9 ;
 wire \i52/n90 ;
 wire \i52/n91 ;
 wire \i52/n92 ;
 wire \i52/n93 ;
 wire \i52/n94 ;
 wire \i52/n95 ;
 wire \i52/n96 ;
 wire \i52/n97 ;
 wire \i52/n98 ;
 wire \i52/n99 ;
 wire \i53/n0 ;
 wire \i53/n1 ;
 wire \i53/n10 ;
 wire \i53/n100 ;
 wire \i53/n101 ;
 wire \i53/n102 ;
 wire \i53/n103 ;
 wire \i53/n104 ;
 wire \i53/n105 ;
 wire \i53/n106 ;
 wire \i53/n107 ;
 wire \i53/n108 ;
 wire \i53/n109 ;
 wire \i53/n11 ;
 wire \i53/n110 ;
 wire \i53/n111 ;
 wire \i53/n112 ;
 wire \i53/n113 ;
 wire \i53/n114 ;
 wire \i53/n115 ;
 wire \i53/n116 ;
 wire \i53/n117 ;
 wire \i53/n118 ;
 wire \i53/n119 ;
 wire \i53/n12 ;
 wire \i53/n120 ;
 wire \i53/n121 ;
 wire \i53/n122 ;
 wire \i53/n123 ;
 wire \i53/n124 ;
 wire \i53/n125 ;
 wire \i53/n126 ;
 wire \i53/n127 ;
 wire \i53/n128 ;
 wire \i53/n129 ;
 wire \i53/n13 ;
 wire \i53/n130 ;
 wire \i53/n131 ;
 wire \i53/n132 ;
 wire \i53/n133 ;
 wire \i53/n134 ;
 wire \i53/n135 ;
 wire \i53/n136 ;
 wire \i53/n137 ;
 wire \i53/n138 ;
 wire \i53/n139 ;
 wire \i53/n14 ;
 wire \i53/n140 ;
 wire \i53/n141 ;
 wire \i53/n142 ;
 wire \i53/n143 ;
 wire \i53/n144 ;
 wire \i53/n145 ;
 wire \i53/n146 ;
 wire \i53/n147 ;
 wire \i53/n148 ;
 wire \i53/n149 ;
 wire \i53/n15 ;
 wire \i53/n150 ;
 wire \i53/n151 ;
 wire \i53/n152 ;
 wire \i53/n153 ;
 wire \i53/n154 ;
 wire \i53/n155 ;
 wire \i53/n156 ;
 wire \i53/n157 ;
 wire \i53/n158 ;
 wire \i53/n159 ;
 wire \i53/n16 ;
 wire \i53/n160 ;
 wire \i53/n161 ;
 wire \i53/n162 ;
 wire \i53/n163 ;
 wire \i53/n164 ;
 wire \i53/n165 ;
 wire \i53/n166 ;
 wire \i53/n167 ;
 wire \i53/n168 ;
 wire \i53/n169 ;
 wire \i53/n17 ;
 wire \i53/n170 ;
 wire \i53/n171 ;
 wire \i53/n172 ;
 wire \i53/n173 ;
 wire \i53/n174 ;
 wire \i53/n175 ;
 wire \i53/n176 ;
 wire \i53/n177 ;
 wire \i53/n178 ;
 wire \i53/n179 ;
 wire \i53/n18 ;
 wire \i53/n180 ;
 wire \i53/n181 ;
 wire \i53/n182 ;
 wire \i53/n183 ;
 wire \i53/n184 ;
 wire \i53/n185 ;
 wire \i53/n186 ;
 wire \i53/n187 ;
 wire \i53/n188 ;
 wire \i53/n189 ;
 wire \i53/n19 ;
 wire \i53/n190 ;
 wire \i53/n191 ;
 wire \i53/n192 ;
 wire \i53/n193 ;
 wire \i53/n194 ;
 wire \i53/n195 ;
 wire \i53/n196 ;
 wire \i53/n197 ;
 wire \i53/n198 ;
 wire \i53/n199 ;
 wire \i53/n2 ;
 wire \i53/n20 ;
 wire \i53/n200 ;
 wire \i53/n201 ;
 wire \i53/n202 ;
 wire \i53/n203 ;
 wire \i53/n204 ;
 wire \i53/n205 ;
 wire \i53/n206 ;
 wire \i53/n207 ;
 wire \i53/n208 ;
 wire \i53/n209 ;
 wire \i53/n21 ;
 wire \i53/n210 ;
 wire \i53/n211 ;
 wire \i53/n212 ;
 wire \i53/n213 ;
 wire \i53/n214 ;
 wire \i53/n215 ;
 wire \i53/n216 ;
 wire \i53/n217 ;
 wire \i53/n218 ;
 wire \i53/n219 ;
 wire \i53/n22 ;
 wire \i53/n220 ;
 wire \i53/n221 ;
 wire \i53/n222 ;
 wire \i53/n223 ;
 wire \i53/n224 ;
 wire \i53/n225 ;
 wire \i53/n226 ;
 wire \i53/n227 ;
 wire \i53/n228 ;
 wire \i53/n229 ;
 wire \i53/n23 ;
 wire \i53/n230 ;
 wire \i53/n231 ;
 wire \i53/n232 ;
 wire \i53/n233 ;
 wire \i53/n234 ;
 wire \i53/n235 ;
 wire \i53/n236 ;
 wire \i53/n237 ;
 wire \i53/n238 ;
 wire \i53/n239 ;
 wire \i53/n24 ;
 wire \i53/n240 ;
 wire \i53/n241 ;
 wire \i53/n242 ;
 wire \i53/n243 ;
 wire \i53/n244 ;
 wire \i53/n245 ;
 wire \i53/n246 ;
 wire \i53/n247 ;
 wire \i53/n248 ;
 wire \i53/n249 ;
 wire \i53/n25 ;
 wire \i53/n250 ;
 wire \i53/n251 ;
 wire \i53/n252 ;
 wire \i53/n253 ;
 wire \i53/n254 ;
 wire \i53/n255 ;
 wire \i53/n256 ;
 wire \i53/n257 ;
 wire \i53/n258 ;
 wire \i53/n259 ;
 wire \i53/n26 ;
 wire \i53/n260 ;
 wire \i53/n261 ;
 wire \i53/n262 ;
 wire \i53/n263 ;
 wire \i53/n264 ;
 wire \i53/n265 ;
 wire \i53/n266 ;
 wire \i53/n267 ;
 wire \i53/n268 ;
 wire \i53/n269 ;
 wire \i53/n27 ;
 wire \i53/n270 ;
 wire \i53/n271 ;
 wire \i53/n272 ;
 wire \i53/n273 ;
 wire \i53/n274 ;
 wire \i53/n275 ;
 wire \i53/n276 ;
 wire \i53/n277 ;
 wire \i53/n278 ;
 wire \i53/n279 ;
 wire \i53/n28 ;
 wire \i53/n280 ;
 wire \i53/n281 ;
 wire \i53/n282 ;
 wire \i53/n283 ;
 wire \i53/n284 ;
 wire \i53/n285 ;
 wire \i53/n286 ;
 wire \i53/n287 ;
 wire \i53/n288 ;
 wire \i53/n289 ;
 wire \i53/n29 ;
 wire \i53/n290 ;
 wire \i53/n291 ;
 wire \i53/n292 ;
 wire \i53/n293 ;
 wire \i53/n294 ;
 wire \i53/n295 ;
 wire \i53/n296 ;
 wire \i53/n297 ;
 wire \i53/n298 ;
 wire \i53/n299 ;
 wire \i53/n3 ;
 wire \i53/n30 ;
 wire \i53/n300 ;
 wire \i53/n301 ;
 wire \i53/n302 ;
 wire \i53/n303 ;
 wire \i53/n304 ;
 wire \i53/n305 ;
 wire \i53/n306 ;
 wire \i53/n307 ;
 wire \i53/n308 ;
 wire \i53/n309 ;
 wire \i53/n31 ;
 wire \i53/n310 ;
 wire \i53/n311 ;
 wire \i53/n312 ;
 wire \i53/n313 ;
 wire \i53/n314 ;
 wire \i53/n315 ;
 wire \i53/n316 ;
 wire \i53/n317 ;
 wire \i53/n318 ;
 wire \i53/n319 ;
 wire \i53/n32 ;
 wire \i53/n320 ;
 wire \i53/n321 ;
 wire \i53/n322 ;
 wire \i53/n323 ;
 wire \i53/n324 ;
 wire \i53/n325 ;
 wire \i53/n326 ;
 wire \i53/n327 ;
 wire \i53/n328 ;
 wire \i53/n329 ;
 wire \i53/n33 ;
 wire \i53/n330 ;
 wire \i53/n331 ;
 wire \i53/n332 ;
 wire \i53/n333 ;
 wire \i53/n334 ;
 wire \i53/n335 ;
 wire \i53/n336 ;
 wire \i53/n337 ;
 wire \i53/n338 ;
 wire \i53/n339 ;
 wire \i53/n34 ;
 wire \i53/n340 ;
 wire \i53/n341 ;
 wire \i53/n342 ;
 wire \i53/n343 ;
 wire \i53/n344 ;
 wire \i53/n345 ;
 wire \i53/n346 ;
 wire \i53/n347 ;
 wire \i53/n348 ;
 wire \i53/n349 ;
 wire \i53/n35 ;
 wire \i53/n350 ;
 wire \i53/n351 ;
 wire \i53/n352 ;
 wire \i53/n353 ;
 wire \i53/n354 ;
 wire \i53/n355 ;
 wire \i53/n356 ;
 wire \i53/n357 ;
 wire \i53/n358 ;
 wire \i53/n359 ;
 wire \i53/n36 ;
 wire \i53/n360 ;
 wire \i53/n361 ;
 wire \i53/n362 ;
 wire \i53/n363 ;
 wire \i53/n364 ;
 wire \i53/n365 ;
 wire \i53/n366 ;
 wire \i53/n367 ;
 wire \i53/n368 ;
 wire \i53/n369 ;
 wire \i53/n37 ;
 wire \i53/n370 ;
 wire \i53/n371 ;
 wire \i53/n372 ;
 wire \i53/n373 ;
 wire \i53/n374 ;
 wire \i53/n375 ;
 wire \i53/n376 ;
 wire \i53/n377 ;
 wire \i53/n378 ;
 wire \i53/n379 ;
 wire \i53/n38 ;
 wire \i53/n380 ;
 wire \i53/n381 ;
 wire \i53/n382 ;
 wire \i53/n383 ;
 wire \i53/n384 ;
 wire \i53/n385 ;
 wire \i53/n386 ;
 wire \i53/n387 ;
 wire \i53/n388 ;
 wire \i53/n389 ;
 wire \i53/n39 ;
 wire \i53/n390 ;
 wire \i53/n391 ;
 wire \i53/n392 ;
 wire \i53/n393 ;
 wire \i53/n394 ;
 wire \i53/n395 ;
 wire \i53/n396 ;
 wire \i53/n397 ;
 wire \i53/n398 ;
 wire \i53/n399 ;
 wire \i53/n4 ;
 wire \i53/n40 ;
 wire \i53/n400 ;
 wire \i53/n401 ;
 wire \i53/n402 ;
 wire \i53/n403 ;
 wire \i53/n404 ;
 wire \i53/n405 ;
 wire \i53/n406 ;
 wire \i53/n407 ;
 wire \i53/n408 ;
 wire \i53/n409 ;
 wire \i53/n41 ;
 wire \i53/n410 ;
 wire \i53/n411 ;
 wire \i53/n412 ;
 wire \i53/n413 ;
 wire \i53/n414 ;
 wire \i53/n415 ;
 wire \i53/n416 ;
 wire \i53/n417 ;
 wire \i53/n418 ;
 wire \i53/n419 ;
 wire \i53/n42 ;
 wire \i53/n420 ;
 wire \i53/n421 ;
 wire \i53/n422 ;
 wire \i53/n423 ;
 wire \i53/n424 ;
 wire \i53/n425 ;
 wire \i53/n426 ;
 wire \i53/n427 ;
 wire \i53/n428 ;
 wire \i53/n429 ;
 wire \i53/n43 ;
 wire \i53/n430 ;
 wire \i53/n431 ;
 wire \i53/n432 ;
 wire \i53/n433 ;
 wire \i53/n434 ;
 wire \i53/n435 ;
 wire \i53/n436 ;
 wire \i53/n437 ;
 wire \i53/n438 ;
 wire \i53/n439 ;
 wire \i53/n44 ;
 wire \i53/n440 ;
 wire \i53/n441 ;
 wire \i53/n442 ;
 wire \i53/n443 ;
 wire \i53/n444 ;
 wire \i53/n445 ;
 wire \i53/n446 ;
 wire \i53/n447 ;
 wire \i53/n448 ;
 wire \i53/n449 ;
 wire \i53/n45 ;
 wire \i53/n450 ;
 wire \i53/n451 ;
 wire \i53/n452 ;
 wire \i53/n453 ;
 wire \i53/n454 ;
 wire \i53/n455 ;
 wire \i53/n456 ;
 wire \i53/n457 ;
 wire \i53/n458 ;
 wire \i53/n459 ;
 wire \i53/n46 ;
 wire \i53/n460 ;
 wire \i53/n461 ;
 wire \i53/n462 ;
 wire \i53/n463 ;
 wire \i53/n464 ;
 wire \i53/n465 ;
 wire \i53/n466 ;
 wire \i53/n467 ;
 wire \i53/n468 ;
 wire \i53/n469 ;
 wire \i53/n47 ;
 wire \i53/n470 ;
 wire \i53/n471 ;
 wire \i53/n472 ;
 wire \i53/n473 ;
 wire \i53/n474 ;
 wire \i53/n475 ;
 wire \i53/n476 ;
 wire \i53/n477 ;
 wire \i53/n478 ;
 wire \i53/n479 ;
 wire \i53/n48 ;
 wire \i53/n480 ;
 wire \i53/n481 ;
 wire \i53/n482 ;
 wire \i53/n483 ;
 wire \i53/n484 ;
 wire \i53/n485 ;
 wire \i53/n486 ;
 wire \i53/n487 ;
 wire \i53/n488 ;
 wire \i53/n489 ;
 wire \i53/n49 ;
 wire \i53/n490 ;
 wire \i53/n491 ;
 wire \i53/n492 ;
 wire \i53/n493 ;
 wire \i53/n494 ;
 wire \i53/n495 ;
 wire \i53/n496 ;
 wire \i53/n497 ;
 wire \i53/n498 ;
 wire \i53/n499 ;
 wire \i53/n5 ;
 wire \i53/n50 ;
 wire \i53/n500 ;
 wire \i53/n501 ;
 wire \i53/n502 ;
 wire \i53/n503 ;
 wire \i53/n504 ;
 wire \i53/n505 ;
 wire \i53/n506 ;
 wire \i53/n507 ;
 wire \i53/n508 ;
 wire \i53/n509 ;
 wire \i53/n51 ;
 wire \i53/n510 ;
 wire \i53/n511 ;
 wire \i53/n512 ;
 wire \i53/n513 ;
 wire \i53/n514 ;
 wire \i53/n515 ;
 wire \i53/n516 ;
 wire \i53/n517 ;
 wire \i53/n518 ;
 wire \i53/n519 ;
 wire \i53/n52 ;
 wire \i53/n520 ;
 wire \i53/n521 ;
 wire \i53/n522 ;
 wire \i53/n523 ;
 wire \i53/n524 ;
 wire \i53/n525 ;
 wire \i53/n526 ;
 wire \i53/n527 ;
 wire \i53/n528 ;
 wire \i53/n529 ;
 wire \i53/n53 ;
 wire \i53/n530 ;
 wire \i53/n531 ;
 wire \i53/n532 ;
 wire \i53/n533 ;
 wire \i53/n534 ;
 wire \i53/n535 ;
 wire \i53/n536 ;
 wire \i53/n537 ;
 wire \i53/n538 ;
 wire \i53/n539 ;
 wire \i53/n54 ;
 wire \i53/n540 ;
 wire \i53/n541 ;
 wire \i53/n542 ;
 wire \i53/n543 ;
 wire \i53/n544 ;
 wire \i53/n545 ;
 wire \i53/n546 ;
 wire \i53/n547 ;
 wire \i53/n548 ;
 wire \i53/n549 ;
 wire \i53/n55 ;
 wire \i53/n550 ;
 wire \i53/n551 ;
 wire \i53/n552 ;
 wire \i53/n553 ;
 wire \i53/n554 ;
 wire \i53/n555 ;
 wire \i53/n556 ;
 wire \i53/n557 ;
 wire \i53/n558 ;
 wire \i53/n559 ;
 wire \i53/n56 ;
 wire \i53/n560 ;
 wire \i53/n561 ;
 wire \i53/n562 ;
 wire \i53/n563 ;
 wire \i53/n564 ;
 wire \i53/n565 ;
 wire \i53/n566 ;
 wire \i53/n567 ;
 wire \i53/n568 ;
 wire \i53/n569 ;
 wire \i53/n57 ;
 wire \i53/n570 ;
 wire \i53/n571 ;
 wire \i53/n572 ;
 wire \i53/n573 ;
 wire \i53/n574 ;
 wire \i53/n575 ;
 wire \i53/n576 ;
 wire \i53/n577 ;
 wire \i53/n578 ;
 wire \i53/n579 ;
 wire \i53/n58 ;
 wire \i53/n580 ;
 wire \i53/n581 ;
 wire \i53/n582 ;
 wire \i53/n583 ;
 wire \i53/n584 ;
 wire \i53/n59 ;
 wire \i53/n6 ;
 wire \i53/n60 ;
 wire \i53/n61 ;
 wire \i53/n62 ;
 wire \i53/n63 ;
 wire \i53/n64 ;
 wire \i53/n65 ;
 wire \i53/n66 ;
 wire \i53/n67 ;
 wire \i53/n68 ;
 wire \i53/n69 ;
 wire \i53/n7 ;
 wire \i53/n70 ;
 wire \i53/n71 ;
 wire \i53/n72 ;
 wire \i53/n73 ;
 wire \i53/n74 ;
 wire \i53/n75 ;
 wire \i53/n76 ;
 wire \i53/n77 ;
 wire \i53/n78 ;
 wire \i53/n79 ;
 wire \i53/n8 ;
 wire \i53/n80 ;
 wire \i53/n81 ;
 wire \i53/n82 ;
 wire \i53/n83 ;
 wire \i53/n84 ;
 wire \i53/n85 ;
 wire \i53/n86 ;
 wire \i53/n87 ;
 wire \i53/n88 ;
 wire \i53/n89 ;
 wire \i53/n9 ;
 wire \i53/n90 ;
 wire \i53/n91 ;
 wire \i53/n92 ;
 wire \i53/n93 ;
 wire \i53/n94 ;
 wire \i53/n95 ;
 wire \i53/n96 ;
 wire \i53/n97 ;
 wire \i53/n98 ;
 wire \i53/n99 ;
 wire \i54/n0 ;
 wire \i54/n1 ;
 wire \i54/n10 ;
 wire \i54/n100 ;
 wire \i54/n101 ;
 wire \i54/n102 ;
 wire \i54/n103 ;
 wire \i54/n104 ;
 wire \i54/n105 ;
 wire \i54/n106 ;
 wire \i54/n107 ;
 wire \i54/n108 ;
 wire \i54/n109 ;
 wire \i54/n11 ;
 wire \i54/n110 ;
 wire \i54/n111 ;
 wire \i54/n112 ;
 wire \i54/n113 ;
 wire \i54/n114 ;
 wire \i54/n115 ;
 wire \i54/n116 ;
 wire \i54/n117 ;
 wire \i54/n118 ;
 wire \i54/n119 ;
 wire \i54/n12 ;
 wire \i54/n120 ;
 wire \i54/n121 ;
 wire \i54/n122 ;
 wire \i54/n123 ;
 wire \i54/n124 ;
 wire \i54/n125 ;
 wire \i54/n126 ;
 wire \i54/n127 ;
 wire \i54/n128 ;
 wire \i54/n129 ;
 wire \i54/n13 ;
 wire \i54/n130 ;
 wire \i54/n131 ;
 wire \i54/n132 ;
 wire \i54/n133 ;
 wire \i54/n134 ;
 wire \i54/n135 ;
 wire \i54/n136 ;
 wire \i54/n137 ;
 wire \i54/n138 ;
 wire \i54/n139 ;
 wire \i54/n14 ;
 wire \i54/n140 ;
 wire \i54/n141 ;
 wire \i54/n142 ;
 wire \i54/n143 ;
 wire \i54/n144 ;
 wire \i54/n145 ;
 wire \i54/n146 ;
 wire \i54/n147 ;
 wire \i54/n148 ;
 wire \i54/n149 ;
 wire \i54/n15 ;
 wire \i54/n150 ;
 wire \i54/n151 ;
 wire \i54/n152 ;
 wire \i54/n153 ;
 wire \i54/n154 ;
 wire \i54/n155 ;
 wire \i54/n156 ;
 wire \i54/n157 ;
 wire \i54/n158 ;
 wire \i54/n159 ;
 wire \i54/n16 ;
 wire \i54/n160 ;
 wire \i54/n161 ;
 wire \i54/n162 ;
 wire \i54/n163 ;
 wire \i54/n164 ;
 wire \i54/n165 ;
 wire \i54/n166 ;
 wire \i54/n167 ;
 wire \i54/n168 ;
 wire \i54/n169 ;
 wire \i54/n17 ;
 wire \i54/n170 ;
 wire \i54/n171 ;
 wire \i54/n172 ;
 wire \i54/n173 ;
 wire \i54/n174 ;
 wire \i54/n175 ;
 wire \i54/n176 ;
 wire \i54/n177 ;
 wire \i54/n178 ;
 wire \i54/n179 ;
 wire \i54/n18 ;
 wire \i54/n180 ;
 wire \i54/n181 ;
 wire \i54/n182 ;
 wire \i54/n183 ;
 wire \i54/n184 ;
 wire \i54/n185 ;
 wire \i54/n186 ;
 wire \i54/n187 ;
 wire \i54/n188 ;
 wire \i54/n189 ;
 wire \i54/n19 ;
 wire \i54/n190 ;
 wire \i54/n191 ;
 wire \i54/n192 ;
 wire \i54/n193 ;
 wire \i54/n194 ;
 wire \i54/n195 ;
 wire \i54/n196 ;
 wire \i54/n197 ;
 wire \i54/n198 ;
 wire \i54/n199 ;
 wire \i54/n2 ;
 wire \i54/n20 ;
 wire \i54/n200 ;
 wire \i54/n201 ;
 wire \i54/n202 ;
 wire \i54/n203 ;
 wire \i54/n204 ;
 wire \i54/n205 ;
 wire \i54/n206 ;
 wire \i54/n207 ;
 wire \i54/n208 ;
 wire \i54/n209 ;
 wire \i54/n21 ;
 wire \i54/n210 ;
 wire \i54/n211 ;
 wire \i54/n212 ;
 wire \i54/n213 ;
 wire \i54/n214 ;
 wire \i54/n215 ;
 wire \i54/n216 ;
 wire \i54/n217 ;
 wire \i54/n218 ;
 wire \i54/n219 ;
 wire \i54/n22 ;
 wire \i54/n220 ;
 wire \i54/n221 ;
 wire \i54/n222 ;
 wire \i54/n223 ;
 wire \i54/n224 ;
 wire \i54/n225 ;
 wire \i54/n226 ;
 wire \i54/n227 ;
 wire \i54/n228 ;
 wire \i54/n229 ;
 wire \i54/n23 ;
 wire \i54/n230 ;
 wire \i54/n231 ;
 wire \i54/n232 ;
 wire \i54/n233 ;
 wire \i54/n234 ;
 wire \i54/n235 ;
 wire \i54/n236 ;
 wire \i54/n237 ;
 wire \i54/n238 ;
 wire \i54/n239 ;
 wire \i54/n24 ;
 wire \i54/n240 ;
 wire \i54/n241 ;
 wire \i54/n242 ;
 wire \i54/n243 ;
 wire \i54/n244 ;
 wire \i54/n245 ;
 wire \i54/n246 ;
 wire \i54/n247 ;
 wire \i54/n248 ;
 wire \i54/n249 ;
 wire \i54/n25 ;
 wire \i54/n250 ;
 wire \i54/n251 ;
 wire \i54/n252 ;
 wire \i54/n253 ;
 wire \i54/n254 ;
 wire \i54/n255 ;
 wire \i54/n256 ;
 wire \i54/n257 ;
 wire \i54/n258 ;
 wire \i54/n259 ;
 wire \i54/n26 ;
 wire \i54/n260 ;
 wire \i54/n261 ;
 wire \i54/n262 ;
 wire \i54/n263 ;
 wire \i54/n264 ;
 wire \i54/n265 ;
 wire \i54/n266 ;
 wire \i54/n267 ;
 wire \i54/n268 ;
 wire \i54/n269 ;
 wire \i54/n27 ;
 wire \i54/n270 ;
 wire \i54/n271 ;
 wire \i54/n272 ;
 wire \i54/n273 ;
 wire \i54/n274 ;
 wire \i54/n275 ;
 wire \i54/n276 ;
 wire \i54/n277 ;
 wire \i54/n278 ;
 wire \i54/n279 ;
 wire \i54/n28 ;
 wire \i54/n280 ;
 wire \i54/n281 ;
 wire \i54/n282 ;
 wire \i54/n283 ;
 wire \i54/n284 ;
 wire \i54/n285 ;
 wire \i54/n286 ;
 wire \i54/n287 ;
 wire \i54/n288 ;
 wire \i54/n289 ;
 wire \i54/n29 ;
 wire \i54/n290 ;
 wire \i54/n291 ;
 wire \i54/n292 ;
 wire \i54/n293 ;
 wire \i54/n294 ;
 wire \i54/n295 ;
 wire \i54/n296 ;
 wire \i54/n297 ;
 wire \i54/n298 ;
 wire \i54/n299 ;
 wire \i54/n3 ;
 wire \i54/n30 ;
 wire \i54/n300 ;
 wire \i54/n301 ;
 wire \i54/n302 ;
 wire \i54/n303 ;
 wire \i54/n304 ;
 wire \i54/n305 ;
 wire \i54/n306 ;
 wire \i54/n307 ;
 wire \i54/n308 ;
 wire \i54/n309 ;
 wire \i54/n31 ;
 wire \i54/n310 ;
 wire \i54/n311 ;
 wire \i54/n312 ;
 wire \i54/n313 ;
 wire \i54/n314 ;
 wire \i54/n315 ;
 wire \i54/n316 ;
 wire \i54/n317 ;
 wire \i54/n318 ;
 wire \i54/n319 ;
 wire \i54/n32 ;
 wire \i54/n320 ;
 wire \i54/n321 ;
 wire \i54/n322 ;
 wire \i54/n323 ;
 wire \i54/n324 ;
 wire \i54/n325 ;
 wire \i54/n326 ;
 wire \i54/n327 ;
 wire \i54/n328 ;
 wire \i54/n329 ;
 wire \i54/n33 ;
 wire \i54/n330 ;
 wire \i54/n331 ;
 wire \i54/n332 ;
 wire \i54/n333 ;
 wire \i54/n334 ;
 wire \i54/n335 ;
 wire \i54/n336 ;
 wire \i54/n337 ;
 wire \i54/n338 ;
 wire \i54/n339 ;
 wire \i54/n34 ;
 wire \i54/n340 ;
 wire \i54/n341 ;
 wire \i54/n342 ;
 wire \i54/n343 ;
 wire \i54/n344 ;
 wire \i54/n345 ;
 wire \i54/n346 ;
 wire \i54/n347 ;
 wire \i54/n348 ;
 wire \i54/n349 ;
 wire \i54/n35 ;
 wire \i54/n350 ;
 wire \i54/n351 ;
 wire \i54/n352 ;
 wire \i54/n353 ;
 wire \i54/n354 ;
 wire \i54/n355 ;
 wire \i54/n356 ;
 wire \i54/n357 ;
 wire \i54/n358 ;
 wire \i54/n359 ;
 wire \i54/n36 ;
 wire \i54/n360 ;
 wire \i54/n361 ;
 wire \i54/n362 ;
 wire \i54/n363 ;
 wire \i54/n364 ;
 wire \i54/n365 ;
 wire \i54/n366 ;
 wire \i54/n367 ;
 wire \i54/n368 ;
 wire \i54/n369 ;
 wire \i54/n37 ;
 wire \i54/n370 ;
 wire \i54/n371 ;
 wire \i54/n372 ;
 wire \i54/n373 ;
 wire \i54/n374 ;
 wire \i54/n375 ;
 wire \i54/n376 ;
 wire \i54/n377 ;
 wire \i54/n378 ;
 wire \i54/n379 ;
 wire \i54/n38 ;
 wire \i54/n380 ;
 wire \i54/n381 ;
 wire \i54/n382 ;
 wire \i54/n383 ;
 wire \i54/n384 ;
 wire \i54/n385 ;
 wire \i54/n386 ;
 wire \i54/n387 ;
 wire \i54/n388 ;
 wire \i54/n389 ;
 wire \i54/n39 ;
 wire \i54/n390 ;
 wire \i54/n391 ;
 wire \i54/n392 ;
 wire \i54/n393 ;
 wire \i54/n394 ;
 wire \i54/n395 ;
 wire \i54/n396 ;
 wire \i54/n397 ;
 wire \i54/n398 ;
 wire \i54/n399 ;
 wire \i54/n4 ;
 wire \i54/n40 ;
 wire \i54/n400 ;
 wire \i54/n401 ;
 wire \i54/n402 ;
 wire \i54/n403 ;
 wire \i54/n404 ;
 wire \i54/n405 ;
 wire \i54/n406 ;
 wire \i54/n407 ;
 wire \i54/n408 ;
 wire \i54/n409 ;
 wire \i54/n41 ;
 wire \i54/n410 ;
 wire \i54/n411 ;
 wire \i54/n412 ;
 wire \i54/n413 ;
 wire \i54/n414 ;
 wire \i54/n415 ;
 wire \i54/n416 ;
 wire \i54/n417 ;
 wire \i54/n418 ;
 wire \i54/n419 ;
 wire \i54/n42 ;
 wire \i54/n420 ;
 wire \i54/n421 ;
 wire \i54/n422 ;
 wire \i54/n423 ;
 wire \i54/n424 ;
 wire \i54/n425 ;
 wire \i54/n426 ;
 wire \i54/n427 ;
 wire \i54/n428 ;
 wire \i54/n429 ;
 wire \i54/n43 ;
 wire \i54/n430 ;
 wire \i54/n431 ;
 wire \i54/n432 ;
 wire \i54/n433 ;
 wire \i54/n434 ;
 wire \i54/n435 ;
 wire \i54/n436 ;
 wire \i54/n437 ;
 wire \i54/n438 ;
 wire \i54/n439 ;
 wire \i54/n44 ;
 wire \i54/n440 ;
 wire \i54/n441 ;
 wire \i54/n442 ;
 wire \i54/n443 ;
 wire \i54/n444 ;
 wire \i54/n445 ;
 wire \i54/n446 ;
 wire \i54/n447 ;
 wire \i54/n448 ;
 wire \i54/n449 ;
 wire \i54/n45 ;
 wire \i54/n450 ;
 wire \i54/n451 ;
 wire \i54/n452 ;
 wire \i54/n453 ;
 wire \i54/n454 ;
 wire \i54/n455 ;
 wire \i54/n456 ;
 wire \i54/n457 ;
 wire \i54/n458 ;
 wire \i54/n459 ;
 wire \i54/n46 ;
 wire \i54/n460 ;
 wire \i54/n461 ;
 wire \i54/n462 ;
 wire \i54/n463 ;
 wire \i54/n464 ;
 wire \i54/n465 ;
 wire \i54/n466 ;
 wire \i54/n467 ;
 wire \i54/n468 ;
 wire \i54/n469 ;
 wire \i54/n47 ;
 wire \i54/n470 ;
 wire \i54/n471 ;
 wire \i54/n472 ;
 wire \i54/n473 ;
 wire \i54/n474 ;
 wire \i54/n475 ;
 wire \i54/n476 ;
 wire \i54/n477 ;
 wire \i54/n478 ;
 wire \i54/n479 ;
 wire \i54/n48 ;
 wire \i54/n480 ;
 wire \i54/n481 ;
 wire \i54/n482 ;
 wire \i54/n483 ;
 wire \i54/n484 ;
 wire \i54/n485 ;
 wire \i54/n486 ;
 wire \i54/n487 ;
 wire \i54/n488 ;
 wire \i54/n489 ;
 wire \i54/n49 ;
 wire \i54/n490 ;
 wire \i54/n491 ;
 wire \i54/n492 ;
 wire \i54/n493 ;
 wire \i54/n494 ;
 wire \i54/n495 ;
 wire \i54/n496 ;
 wire \i54/n497 ;
 wire \i54/n498 ;
 wire \i54/n499 ;
 wire \i54/n5 ;
 wire \i54/n50 ;
 wire \i54/n500 ;
 wire \i54/n501 ;
 wire \i54/n502 ;
 wire \i54/n503 ;
 wire \i54/n504 ;
 wire \i54/n505 ;
 wire \i54/n506 ;
 wire \i54/n507 ;
 wire \i54/n508 ;
 wire \i54/n509 ;
 wire \i54/n51 ;
 wire \i54/n510 ;
 wire \i54/n511 ;
 wire \i54/n512 ;
 wire \i54/n513 ;
 wire \i54/n514 ;
 wire \i54/n515 ;
 wire \i54/n516 ;
 wire \i54/n517 ;
 wire \i54/n518 ;
 wire \i54/n519 ;
 wire \i54/n52 ;
 wire \i54/n520 ;
 wire \i54/n521 ;
 wire \i54/n522 ;
 wire \i54/n523 ;
 wire \i54/n524 ;
 wire \i54/n525 ;
 wire \i54/n526 ;
 wire \i54/n527 ;
 wire \i54/n528 ;
 wire \i54/n529 ;
 wire \i54/n53 ;
 wire \i54/n530 ;
 wire \i54/n531 ;
 wire \i54/n532 ;
 wire \i54/n533 ;
 wire \i54/n534 ;
 wire \i54/n535 ;
 wire \i54/n536 ;
 wire \i54/n537 ;
 wire \i54/n538 ;
 wire \i54/n539 ;
 wire \i54/n54 ;
 wire \i54/n540 ;
 wire \i54/n541 ;
 wire \i54/n542 ;
 wire \i54/n543 ;
 wire \i54/n544 ;
 wire \i54/n545 ;
 wire \i54/n546 ;
 wire \i54/n547 ;
 wire \i54/n548 ;
 wire \i54/n549 ;
 wire \i54/n55 ;
 wire \i54/n550 ;
 wire \i54/n551 ;
 wire \i54/n552 ;
 wire \i54/n553 ;
 wire \i54/n554 ;
 wire \i54/n555 ;
 wire \i54/n556 ;
 wire \i54/n557 ;
 wire \i54/n558 ;
 wire \i54/n559 ;
 wire \i54/n56 ;
 wire \i54/n560 ;
 wire \i54/n561 ;
 wire \i54/n562 ;
 wire \i54/n563 ;
 wire \i54/n564 ;
 wire \i54/n565 ;
 wire \i54/n566 ;
 wire \i54/n567 ;
 wire \i54/n568 ;
 wire \i54/n569 ;
 wire \i54/n57 ;
 wire \i54/n570 ;
 wire \i54/n571 ;
 wire \i54/n572 ;
 wire \i54/n573 ;
 wire \i54/n574 ;
 wire \i54/n575 ;
 wire \i54/n576 ;
 wire \i54/n577 ;
 wire \i54/n578 ;
 wire \i54/n579 ;
 wire \i54/n58 ;
 wire \i54/n580 ;
 wire \i54/n581 ;
 wire \i54/n59 ;
 wire \i54/n6 ;
 wire \i54/n60 ;
 wire \i54/n61 ;
 wire \i54/n62 ;
 wire \i54/n63 ;
 wire \i54/n64 ;
 wire \i54/n65 ;
 wire \i54/n66 ;
 wire \i54/n67 ;
 wire \i54/n68 ;
 wire \i54/n69 ;
 wire \i54/n7 ;
 wire \i54/n70 ;
 wire \i54/n71 ;
 wire \i54/n72 ;
 wire \i54/n73 ;
 wire \i54/n74 ;
 wire \i54/n75 ;
 wire \i54/n76 ;
 wire \i54/n77 ;
 wire \i54/n78 ;
 wire \i54/n79 ;
 wire \i54/n8 ;
 wire \i54/n80 ;
 wire \i54/n81 ;
 wire \i54/n82 ;
 wire \i54/n83 ;
 wire \i54/n84 ;
 wire \i54/n85 ;
 wire \i54/n86 ;
 wire \i54/n87 ;
 wire \i54/n88 ;
 wire \i54/n89 ;
 wire \i54/n9 ;
 wire \i54/n90 ;
 wire \i54/n91 ;
 wire \i54/n92 ;
 wire \i54/n93 ;
 wire \i54/n94 ;
 wire \i54/n95 ;
 wire \i54/n96 ;
 wire \i54/n97 ;
 wire \i54/n98 ;
 wire \i54/n99 ;
 wire \i55/n0 ;
 wire \i55/n1 ;
 wire \i55/n10 ;
 wire \i55/n100 ;
 wire \i55/n101 ;
 wire \i55/n102 ;
 wire \i55/n103 ;
 wire \i55/n104 ;
 wire \i55/n105 ;
 wire \i55/n106 ;
 wire \i55/n107 ;
 wire \i55/n108 ;
 wire \i55/n109 ;
 wire \i55/n11 ;
 wire \i55/n110 ;
 wire \i55/n111 ;
 wire \i55/n112 ;
 wire \i55/n113 ;
 wire \i55/n114 ;
 wire \i55/n115 ;
 wire \i55/n116 ;
 wire \i55/n117 ;
 wire \i55/n118 ;
 wire \i55/n119 ;
 wire \i55/n12 ;
 wire \i55/n120 ;
 wire \i55/n121 ;
 wire \i55/n122 ;
 wire \i55/n123 ;
 wire \i55/n124 ;
 wire \i55/n125 ;
 wire \i55/n126 ;
 wire \i55/n127 ;
 wire \i55/n128 ;
 wire \i55/n129 ;
 wire \i55/n13 ;
 wire \i55/n130 ;
 wire \i55/n131 ;
 wire \i55/n132 ;
 wire \i55/n133 ;
 wire \i55/n134 ;
 wire \i55/n135 ;
 wire \i55/n136 ;
 wire \i55/n137 ;
 wire \i55/n138 ;
 wire \i55/n139 ;
 wire \i55/n14 ;
 wire \i55/n140 ;
 wire \i55/n141 ;
 wire \i55/n142 ;
 wire \i55/n143 ;
 wire \i55/n144 ;
 wire \i55/n145 ;
 wire \i55/n146 ;
 wire \i55/n147 ;
 wire \i55/n148 ;
 wire \i55/n149 ;
 wire \i55/n15 ;
 wire \i55/n150 ;
 wire \i55/n151 ;
 wire \i55/n152 ;
 wire \i55/n153 ;
 wire \i55/n154 ;
 wire \i55/n155 ;
 wire \i55/n156 ;
 wire \i55/n157 ;
 wire \i55/n158 ;
 wire \i55/n159 ;
 wire \i55/n16 ;
 wire \i55/n160 ;
 wire \i55/n161 ;
 wire \i55/n162 ;
 wire \i55/n163 ;
 wire \i55/n164 ;
 wire \i55/n165 ;
 wire \i55/n166 ;
 wire \i55/n167 ;
 wire \i55/n168 ;
 wire \i55/n169 ;
 wire \i55/n17 ;
 wire \i55/n170 ;
 wire \i55/n171 ;
 wire \i55/n172 ;
 wire \i55/n173 ;
 wire \i55/n174 ;
 wire \i55/n175 ;
 wire \i55/n176 ;
 wire \i55/n177 ;
 wire \i55/n178 ;
 wire \i55/n179 ;
 wire \i55/n18 ;
 wire \i55/n180 ;
 wire \i55/n181 ;
 wire \i55/n182 ;
 wire \i55/n183 ;
 wire \i55/n184 ;
 wire \i55/n185 ;
 wire \i55/n186 ;
 wire \i55/n187 ;
 wire \i55/n188 ;
 wire \i55/n189 ;
 wire \i55/n19 ;
 wire \i55/n190 ;
 wire \i55/n191 ;
 wire \i55/n192 ;
 wire \i55/n193 ;
 wire \i55/n194 ;
 wire \i55/n195 ;
 wire \i55/n196 ;
 wire \i55/n197 ;
 wire \i55/n198 ;
 wire \i55/n199 ;
 wire \i55/n2 ;
 wire \i55/n20 ;
 wire \i55/n200 ;
 wire \i55/n201 ;
 wire \i55/n202 ;
 wire \i55/n203 ;
 wire \i55/n204 ;
 wire \i55/n205 ;
 wire \i55/n206 ;
 wire \i55/n207 ;
 wire \i55/n208 ;
 wire \i55/n209 ;
 wire \i55/n21 ;
 wire \i55/n210 ;
 wire \i55/n211 ;
 wire \i55/n212 ;
 wire \i55/n213 ;
 wire \i55/n214 ;
 wire \i55/n215 ;
 wire \i55/n216 ;
 wire \i55/n217 ;
 wire \i55/n218 ;
 wire \i55/n219 ;
 wire \i55/n22 ;
 wire \i55/n220 ;
 wire \i55/n221 ;
 wire \i55/n222 ;
 wire \i55/n223 ;
 wire \i55/n224 ;
 wire \i55/n225 ;
 wire \i55/n226 ;
 wire \i55/n227 ;
 wire \i55/n228 ;
 wire \i55/n229 ;
 wire \i55/n23 ;
 wire \i55/n230 ;
 wire \i55/n231 ;
 wire \i55/n232 ;
 wire \i55/n233 ;
 wire \i55/n234 ;
 wire \i55/n235 ;
 wire \i55/n236 ;
 wire \i55/n237 ;
 wire \i55/n238 ;
 wire \i55/n239 ;
 wire \i55/n24 ;
 wire \i55/n240 ;
 wire \i55/n241 ;
 wire \i55/n242 ;
 wire \i55/n243 ;
 wire \i55/n244 ;
 wire \i55/n245 ;
 wire \i55/n246 ;
 wire \i55/n247 ;
 wire \i55/n248 ;
 wire \i55/n249 ;
 wire \i55/n25 ;
 wire \i55/n250 ;
 wire \i55/n251 ;
 wire \i55/n252 ;
 wire \i55/n253 ;
 wire \i55/n254 ;
 wire \i55/n255 ;
 wire \i55/n256 ;
 wire \i55/n257 ;
 wire \i55/n258 ;
 wire \i55/n259 ;
 wire \i55/n26 ;
 wire \i55/n260 ;
 wire \i55/n261 ;
 wire \i55/n262 ;
 wire \i55/n263 ;
 wire \i55/n264 ;
 wire \i55/n265 ;
 wire \i55/n266 ;
 wire \i55/n267 ;
 wire \i55/n268 ;
 wire \i55/n269 ;
 wire \i55/n27 ;
 wire \i55/n270 ;
 wire \i55/n271 ;
 wire \i55/n272 ;
 wire \i55/n273 ;
 wire \i55/n274 ;
 wire \i55/n275 ;
 wire \i55/n276 ;
 wire \i55/n277 ;
 wire \i55/n278 ;
 wire \i55/n279 ;
 wire \i55/n28 ;
 wire \i55/n280 ;
 wire \i55/n281 ;
 wire \i55/n282 ;
 wire \i55/n283 ;
 wire \i55/n284 ;
 wire \i55/n285 ;
 wire \i55/n286 ;
 wire \i55/n287 ;
 wire \i55/n288 ;
 wire \i55/n289 ;
 wire \i55/n29 ;
 wire \i55/n290 ;
 wire \i55/n291 ;
 wire \i55/n292 ;
 wire \i55/n293 ;
 wire \i55/n294 ;
 wire \i55/n295 ;
 wire \i55/n296 ;
 wire \i55/n297 ;
 wire \i55/n298 ;
 wire \i55/n299 ;
 wire \i55/n3 ;
 wire \i55/n30 ;
 wire \i55/n300 ;
 wire \i55/n301 ;
 wire \i55/n302 ;
 wire \i55/n303 ;
 wire \i55/n304 ;
 wire \i55/n305 ;
 wire \i55/n306 ;
 wire \i55/n307 ;
 wire \i55/n308 ;
 wire \i55/n309 ;
 wire \i55/n31 ;
 wire \i55/n310 ;
 wire \i55/n311 ;
 wire \i55/n312 ;
 wire \i55/n313 ;
 wire \i55/n314 ;
 wire \i55/n315 ;
 wire \i55/n316 ;
 wire \i55/n317 ;
 wire \i55/n318 ;
 wire \i55/n319 ;
 wire \i55/n32 ;
 wire \i55/n320 ;
 wire \i55/n321 ;
 wire \i55/n322 ;
 wire \i55/n323 ;
 wire \i55/n324 ;
 wire \i55/n325 ;
 wire \i55/n326 ;
 wire \i55/n327 ;
 wire \i55/n328 ;
 wire \i55/n329 ;
 wire \i55/n33 ;
 wire \i55/n330 ;
 wire \i55/n331 ;
 wire \i55/n332 ;
 wire \i55/n333 ;
 wire \i55/n334 ;
 wire \i55/n335 ;
 wire \i55/n336 ;
 wire \i55/n337 ;
 wire \i55/n338 ;
 wire \i55/n339 ;
 wire \i55/n34 ;
 wire \i55/n340 ;
 wire \i55/n341 ;
 wire \i55/n342 ;
 wire \i55/n343 ;
 wire \i55/n344 ;
 wire \i55/n345 ;
 wire \i55/n346 ;
 wire \i55/n347 ;
 wire \i55/n348 ;
 wire \i55/n349 ;
 wire \i55/n35 ;
 wire \i55/n350 ;
 wire \i55/n351 ;
 wire \i55/n352 ;
 wire \i55/n353 ;
 wire \i55/n354 ;
 wire \i55/n355 ;
 wire \i55/n356 ;
 wire \i55/n357 ;
 wire \i55/n358 ;
 wire \i55/n359 ;
 wire \i55/n36 ;
 wire \i55/n360 ;
 wire \i55/n361 ;
 wire \i55/n362 ;
 wire \i55/n363 ;
 wire \i55/n364 ;
 wire \i55/n365 ;
 wire \i55/n366 ;
 wire \i55/n367 ;
 wire \i55/n368 ;
 wire \i55/n369 ;
 wire \i55/n37 ;
 wire \i55/n370 ;
 wire \i55/n371 ;
 wire \i55/n372 ;
 wire \i55/n373 ;
 wire \i55/n374 ;
 wire \i55/n375 ;
 wire \i55/n376 ;
 wire \i55/n377 ;
 wire \i55/n378 ;
 wire \i55/n379 ;
 wire \i55/n38 ;
 wire \i55/n380 ;
 wire \i55/n381 ;
 wire \i55/n382 ;
 wire \i55/n383 ;
 wire \i55/n384 ;
 wire \i55/n385 ;
 wire \i55/n386 ;
 wire \i55/n387 ;
 wire \i55/n388 ;
 wire \i55/n389 ;
 wire \i55/n39 ;
 wire \i55/n390 ;
 wire \i55/n391 ;
 wire \i55/n392 ;
 wire \i55/n393 ;
 wire \i55/n394 ;
 wire \i55/n395 ;
 wire \i55/n396 ;
 wire \i55/n397 ;
 wire \i55/n398 ;
 wire \i55/n399 ;
 wire \i55/n4 ;
 wire \i55/n40 ;
 wire \i55/n400 ;
 wire \i55/n401 ;
 wire \i55/n402 ;
 wire \i55/n403 ;
 wire \i55/n404 ;
 wire \i55/n405 ;
 wire \i55/n406 ;
 wire \i55/n407 ;
 wire \i55/n408 ;
 wire \i55/n409 ;
 wire \i55/n41 ;
 wire \i55/n410 ;
 wire \i55/n411 ;
 wire \i55/n412 ;
 wire \i55/n413 ;
 wire \i55/n414 ;
 wire \i55/n415 ;
 wire \i55/n416 ;
 wire \i55/n417 ;
 wire \i55/n418 ;
 wire \i55/n419 ;
 wire \i55/n42 ;
 wire \i55/n420 ;
 wire \i55/n421 ;
 wire \i55/n422 ;
 wire \i55/n423 ;
 wire \i55/n424 ;
 wire \i55/n425 ;
 wire \i55/n426 ;
 wire \i55/n427 ;
 wire \i55/n428 ;
 wire \i55/n429 ;
 wire \i55/n43 ;
 wire \i55/n430 ;
 wire \i55/n431 ;
 wire \i55/n432 ;
 wire \i55/n433 ;
 wire \i55/n434 ;
 wire \i55/n435 ;
 wire \i55/n436 ;
 wire \i55/n437 ;
 wire \i55/n438 ;
 wire \i55/n439 ;
 wire \i55/n44 ;
 wire \i55/n440 ;
 wire \i55/n441 ;
 wire \i55/n442 ;
 wire \i55/n443 ;
 wire \i55/n444 ;
 wire \i55/n445 ;
 wire \i55/n446 ;
 wire \i55/n447 ;
 wire \i55/n448 ;
 wire \i55/n449 ;
 wire \i55/n45 ;
 wire \i55/n450 ;
 wire \i55/n451 ;
 wire \i55/n452 ;
 wire \i55/n453 ;
 wire \i55/n454 ;
 wire \i55/n455 ;
 wire \i55/n456 ;
 wire \i55/n457 ;
 wire \i55/n458 ;
 wire \i55/n459 ;
 wire \i55/n46 ;
 wire \i55/n460 ;
 wire \i55/n461 ;
 wire \i55/n462 ;
 wire \i55/n463 ;
 wire \i55/n464 ;
 wire \i55/n465 ;
 wire \i55/n466 ;
 wire \i55/n467 ;
 wire \i55/n468 ;
 wire \i55/n469 ;
 wire \i55/n47 ;
 wire \i55/n470 ;
 wire \i55/n471 ;
 wire \i55/n472 ;
 wire \i55/n473 ;
 wire \i55/n474 ;
 wire \i55/n475 ;
 wire \i55/n476 ;
 wire \i55/n477 ;
 wire \i55/n478 ;
 wire \i55/n479 ;
 wire \i55/n48 ;
 wire \i55/n480 ;
 wire \i55/n481 ;
 wire \i55/n482 ;
 wire \i55/n483 ;
 wire \i55/n484 ;
 wire \i55/n485 ;
 wire \i55/n486 ;
 wire \i55/n487 ;
 wire \i55/n488 ;
 wire \i55/n489 ;
 wire \i55/n49 ;
 wire \i55/n490 ;
 wire \i55/n491 ;
 wire \i55/n492 ;
 wire \i55/n493 ;
 wire \i55/n494 ;
 wire \i55/n495 ;
 wire \i55/n496 ;
 wire \i55/n497 ;
 wire \i55/n498 ;
 wire \i55/n499 ;
 wire \i55/n5 ;
 wire \i55/n50 ;
 wire \i55/n500 ;
 wire \i55/n501 ;
 wire \i55/n502 ;
 wire \i55/n503 ;
 wire \i55/n504 ;
 wire \i55/n505 ;
 wire \i55/n506 ;
 wire \i55/n507 ;
 wire \i55/n508 ;
 wire \i55/n509 ;
 wire \i55/n51 ;
 wire \i55/n510 ;
 wire \i55/n511 ;
 wire \i55/n512 ;
 wire \i55/n513 ;
 wire \i55/n514 ;
 wire \i55/n515 ;
 wire \i55/n516 ;
 wire \i55/n517 ;
 wire \i55/n518 ;
 wire \i55/n519 ;
 wire \i55/n52 ;
 wire \i55/n520 ;
 wire \i55/n521 ;
 wire \i55/n522 ;
 wire \i55/n523 ;
 wire \i55/n524 ;
 wire \i55/n525 ;
 wire \i55/n526 ;
 wire \i55/n527 ;
 wire \i55/n528 ;
 wire \i55/n529 ;
 wire \i55/n53 ;
 wire \i55/n530 ;
 wire \i55/n531 ;
 wire \i55/n532 ;
 wire \i55/n533 ;
 wire \i55/n534 ;
 wire \i55/n535 ;
 wire \i55/n536 ;
 wire \i55/n537 ;
 wire \i55/n538 ;
 wire \i55/n539 ;
 wire \i55/n54 ;
 wire \i55/n540 ;
 wire \i55/n541 ;
 wire \i55/n542 ;
 wire \i55/n543 ;
 wire \i55/n544 ;
 wire \i55/n545 ;
 wire \i55/n546 ;
 wire \i55/n547 ;
 wire \i55/n548 ;
 wire \i55/n549 ;
 wire \i55/n55 ;
 wire \i55/n550 ;
 wire \i55/n551 ;
 wire \i55/n552 ;
 wire \i55/n553 ;
 wire \i55/n554 ;
 wire \i55/n555 ;
 wire \i55/n556 ;
 wire \i55/n557 ;
 wire \i55/n558 ;
 wire \i55/n559 ;
 wire \i55/n56 ;
 wire \i55/n560 ;
 wire \i55/n561 ;
 wire \i55/n562 ;
 wire \i55/n563 ;
 wire \i55/n564 ;
 wire \i55/n565 ;
 wire \i55/n566 ;
 wire \i55/n567 ;
 wire \i55/n568 ;
 wire \i55/n569 ;
 wire \i55/n57 ;
 wire \i55/n570 ;
 wire \i55/n571 ;
 wire \i55/n572 ;
 wire \i55/n573 ;
 wire \i55/n574 ;
 wire \i55/n575 ;
 wire \i55/n576 ;
 wire \i55/n577 ;
 wire \i55/n578 ;
 wire \i55/n579 ;
 wire \i55/n58 ;
 wire \i55/n580 ;
 wire \i55/n581 ;
 wire \i55/n59 ;
 wire \i55/n6 ;
 wire \i55/n60 ;
 wire \i55/n61 ;
 wire \i55/n62 ;
 wire \i55/n63 ;
 wire \i55/n64 ;
 wire \i55/n65 ;
 wire \i55/n66 ;
 wire \i55/n67 ;
 wire \i55/n68 ;
 wire \i55/n69 ;
 wire \i55/n7 ;
 wire \i55/n70 ;
 wire \i55/n71 ;
 wire \i55/n72 ;
 wire \i55/n73 ;
 wire \i55/n74 ;
 wire \i55/n75 ;
 wire \i55/n76 ;
 wire \i55/n77 ;
 wire \i55/n78 ;
 wire \i55/n79 ;
 wire \i55/n8 ;
 wire \i55/n80 ;
 wire \i55/n81 ;
 wire \i55/n82 ;
 wire \i55/n83 ;
 wire \i55/n84 ;
 wire \i55/n85 ;
 wire \i55/n86 ;
 wire \i55/n87 ;
 wire \i55/n88 ;
 wire \i55/n89 ;
 wire \i55/n9 ;
 wire \i55/n90 ;
 wire \i55/n91 ;
 wire \i55/n92 ;
 wire \i55/n93 ;
 wire \i55/n94 ;
 wire \i55/n95 ;
 wire \i55/n96 ;
 wire \i55/n97 ;
 wire \i55/n98 ;
 wire \i55/n99 ;
 wire \i56/n0 ;
 wire \i56/n1 ;
 wire \i56/n10 ;
 wire \i56/n100 ;
 wire \i56/n101 ;
 wire \i56/n102 ;
 wire \i56/n103 ;
 wire \i56/n104 ;
 wire \i56/n105 ;
 wire \i56/n106 ;
 wire \i56/n107 ;
 wire \i56/n108 ;
 wire \i56/n109 ;
 wire \i56/n11 ;
 wire \i56/n110 ;
 wire \i56/n111 ;
 wire \i56/n112 ;
 wire \i56/n113 ;
 wire \i56/n114 ;
 wire \i56/n115 ;
 wire \i56/n116 ;
 wire \i56/n117 ;
 wire \i56/n118 ;
 wire \i56/n119 ;
 wire \i56/n12 ;
 wire \i56/n120 ;
 wire \i56/n121 ;
 wire \i56/n122 ;
 wire \i56/n123 ;
 wire \i56/n124 ;
 wire \i56/n125 ;
 wire \i56/n126 ;
 wire \i56/n127 ;
 wire \i56/n128 ;
 wire \i56/n129 ;
 wire \i56/n13 ;
 wire \i56/n130 ;
 wire \i56/n131 ;
 wire \i56/n132 ;
 wire \i56/n133 ;
 wire \i56/n134 ;
 wire \i56/n135 ;
 wire \i56/n136 ;
 wire \i56/n137 ;
 wire \i56/n138 ;
 wire \i56/n139 ;
 wire \i56/n14 ;
 wire \i56/n140 ;
 wire \i56/n141 ;
 wire \i56/n142 ;
 wire \i56/n143 ;
 wire \i56/n144 ;
 wire \i56/n145 ;
 wire \i56/n146 ;
 wire \i56/n147 ;
 wire \i56/n148 ;
 wire \i56/n149 ;
 wire \i56/n15 ;
 wire \i56/n150 ;
 wire \i56/n151 ;
 wire \i56/n152 ;
 wire \i56/n153 ;
 wire \i56/n154 ;
 wire \i56/n155 ;
 wire \i56/n156 ;
 wire \i56/n157 ;
 wire \i56/n158 ;
 wire \i56/n159 ;
 wire \i56/n16 ;
 wire \i56/n160 ;
 wire \i56/n161 ;
 wire \i56/n162 ;
 wire \i56/n163 ;
 wire \i56/n164 ;
 wire \i56/n165 ;
 wire \i56/n166 ;
 wire \i56/n167 ;
 wire \i56/n168 ;
 wire \i56/n169 ;
 wire \i56/n17 ;
 wire \i56/n170 ;
 wire \i56/n171 ;
 wire \i56/n172 ;
 wire \i56/n173 ;
 wire \i56/n174 ;
 wire \i56/n175 ;
 wire \i56/n176 ;
 wire \i56/n177 ;
 wire \i56/n178 ;
 wire \i56/n179 ;
 wire \i56/n18 ;
 wire \i56/n180 ;
 wire \i56/n181 ;
 wire \i56/n182 ;
 wire \i56/n183 ;
 wire \i56/n184 ;
 wire \i56/n185 ;
 wire \i56/n186 ;
 wire \i56/n187 ;
 wire \i56/n188 ;
 wire \i56/n189 ;
 wire \i56/n19 ;
 wire \i56/n190 ;
 wire \i56/n191 ;
 wire \i56/n192 ;
 wire \i56/n193 ;
 wire \i56/n194 ;
 wire \i56/n195 ;
 wire \i56/n196 ;
 wire \i56/n197 ;
 wire \i56/n198 ;
 wire \i56/n199 ;
 wire \i56/n2 ;
 wire \i56/n20 ;
 wire \i56/n200 ;
 wire \i56/n201 ;
 wire \i56/n202 ;
 wire \i56/n203 ;
 wire \i56/n204 ;
 wire \i56/n205 ;
 wire \i56/n206 ;
 wire \i56/n207 ;
 wire \i56/n208 ;
 wire \i56/n209 ;
 wire \i56/n21 ;
 wire \i56/n210 ;
 wire \i56/n211 ;
 wire \i56/n212 ;
 wire \i56/n213 ;
 wire \i56/n214 ;
 wire \i56/n215 ;
 wire \i56/n216 ;
 wire \i56/n217 ;
 wire \i56/n218 ;
 wire \i56/n219 ;
 wire \i56/n22 ;
 wire \i56/n220 ;
 wire \i56/n221 ;
 wire \i56/n222 ;
 wire \i56/n223 ;
 wire \i56/n224 ;
 wire \i56/n225 ;
 wire \i56/n226 ;
 wire \i56/n227 ;
 wire \i56/n228 ;
 wire \i56/n229 ;
 wire \i56/n23 ;
 wire \i56/n230 ;
 wire \i56/n231 ;
 wire \i56/n232 ;
 wire \i56/n233 ;
 wire \i56/n234 ;
 wire \i56/n235 ;
 wire \i56/n236 ;
 wire \i56/n237 ;
 wire \i56/n238 ;
 wire \i56/n239 ;
 wire \i56/n24 ;
 wire \i56/n240 ;
 wire \i56/n241 ;
 wire \i56/n242 ;
 wire \i56/n243 ;
 wire \i56/n244 ;
 wire \i56/n245 ;
 wire \i56/n246 ;
 wire \i56/n247 ;
 wire \i56/n248 ;
 wire \i56/n249 ;
 wire \i56/n25 ;
 wire \i56/n250 ;
 wire \i56/n251 ;
 wire \i56/n252 ;
 wire \i56/n253 ;
 wire \i56/n254 ;
 wire \i56/n255 ;
 wire \i56/n256 ;
 wire \i56/n257 ;
 wire \i56/n258 ;
 wire \i56/n259 ;
 wire \i56/n26 ;
 wire \i56/n260 ;
 wire \i56/n261 ;
 wire \i56/n262 ;
 wire \i56/n263 ;
 wire \i56/n264 ;
 wire \i56/n265 ;
 wire \i56/n266 ;
 wire \i56/n267 ;
 wire \i56/n268 ;
 wire \i56/n269 ;
 wire \i56/n27 ;
 wire \i56/n270 ;
 wire \i56/n271 ;
 wire \i56/n272 ;
 wire \i56/n273 ;
 wire \i56/n274 ;
 wire \i56/n275 ;
 wire \i56/n276 ;
 wire \i56/n277 ;
 wire \i56/n278 ;
 wire \i56/n279 ;
 wire \i56/n28 ;
 wire \i56/n280 ;
 wire \i56/n281 ;
 wire \i56/n282 ;
 wire \i56/n283 ;
 wire \i56/n284 ;
 wire \i56/n285 ;
 wire \i56/n286 ;
 wire \i56/n287 ;
 wire \i56/n288 ;
 wire \i56/n289 ;
 wire \i56/n29 ;
 wire \i56/n290 ;
 wire \i56/n291 ;
 wire \i56/n292 ;
 wire \i56/n293 ;
 wire \i56/n294 ;
 wire \i56/n295 ;
 wire \i56/n296 ;
 wire \i56/n297 ;
 wire \i56/n298 ;
 wire \i56/n299 ;
 wire \i56/n3 ;
 wire \i56/n30 ;
 wire \i56/n300 ;
 wire \i56/n301 ;
 wire \i56/n302 ;
 wire \i56/n303 ;
 wire \i56/n304 ;
 wire \i56/n305 ;
 wire \i56/n306 ;
 wire \i56/n307 ;
 wire \i56/n308 ;
 wire \i56/n309 ;
 wire \i56/n31 ;
 wire \i56/n310 ;
 wire \i56/n311 ;
 wire \i56/n312 ;
 wire \i56/n313 ;
 wire \i56/n314 ;
 wire \i56/n315 ;
 wire \i56/n316 ;
 wire \i56/n317 ;
 wire \i56/n318 ;
 wire \i56/n319 ;
 wire \i56/n32 ;
 wire \i56/n320 ;
 wire \i56/n321 ;
 wire \i56/n322 ;
 wire \i56/n323 ;
 wire \i56/n324 ;
 wire \i56/n325 ;
 wire \i56/n326 ;
 wire \i56/n327 ;
 wire \i56/n328 ;
 wire \i56/n329 ;
 wire \i56/n33 ;
 wire \i56/n330 ;
 wire \i56/n331 ;
 wire \i56/n332 ;
 wire \i56/n333 ;
 wire \i56/n334 ;
 wire \i56/n335 ;
 wire \i56/n336 ;
 wire \i56/n337 ;
 wire \i56/n338 ;
 wire \i56/n339 ;
 wire \i56/n34 ;
 wire \i56/n340 ;
 wire \i56/n341 ;
 wire \i56/n342 ;
 wire \i56/n343 ;
 wire \i56/n344 ;
 wire \i56/n345 ;
 wire \i56/n346 ;
 wire \i56/n347 ;
 wire \i56/n348 ;
 wire \i56/n349 ;
 wire \i56/n35 ;
 wire \i56/n350 ;
 wire \i56/n351 ;
 wire \i56/n352 ;
 wire \i56/n353 ;
 wire \i56/n354 ;
 wire \i56/n355 ;
 wire \i56/n356 ;
 wire \i56/n357 ;
 wire \i56/n358 ;
 wire \i56/n359 ;
 wire \i56/n36 ;
 wire \i56/n360 ;
 wire \i56/n361 ;
 wire \i56/n362 ;
 wire \i56/n363 ;
 wire \i56/n364 ;
 wire \i56/n365 ;
 wire \i56/n366 ;
 wire \i56/n367 ;
 wire \i56/n368 ;
 wire \i56/n369 ;
 wire \i56/n37 ;
 wire \i56/n370 ;
 wire \i56/n371 ;
 wire \i56/n372 ;
 wire \i56/n373 ;
 wire \i56/n374 ;
 wire \i56/n375 ;
 wire \i56/n376 ;
 wire \i56/n377 ;
 wire \i56/n378 ;
 wire \i56/n379 ;
 wire \i56/n38 ;
 wire \i56/n380 ;
 wire \i56/n381 ;
 wire \i56/n382 ;
 wire \i56/n383 ;
 wire \i56/n384 ;
 wire \i56/n385 ;
 wire \i56/n386 ;
 wire \i56/n387 ;
 wire \i56/n388 ;
 wire \i56/n389 ;
 wire \i56/n39 ;
 wire \i56/n390 ;
 wire \i56/n391 ;
 wire \i56/n392 ;
 wire \i56/n393 ;
 wire \i56/n394 ;
 wire \i56/n395 ;
 wire \i56/n396 ;
 wire \i56/n397 ;
 wire \i56/n398 ;
 wire \i56/n399 ;
 wire \i56/n4 ;
 wire \i56/n40 ;
 wire \i56/n400 ;
 wire \i56/n401 ;
 wire \i56/n402 ;
 wire \i56/n403 ;
 wire \i56/n404 ;
 wire \i56/n405 ;
 wire \i56/n406 ;
 wire \i56/n407 ;
 wire \i56/n408 ;
 wire \i56/n409 ;
 wire \i56/n41 ;
 wire \i56/n410 ;
 wire \i56/n411 ;
 wire \i56/n412 ;
 wire \i56/n413 ;
 wire \i56/n414 ;
 wire \i56/n415 ;
 wire \i56/n416 ;
 wire \i56/n417 ;
 wire \i56/n418 ;
 wire \i56/n419 ;
 wire \i56/n42 ;
 wire \i56/n420 ;
 wire \i56/n421 ;
 wire \i56/n422 ;
 wire \i56/n423 ;
 wire \i56/n424 ;
 wire \i56/n425 ;
 wire \i56/n426 ;
 wire \i56/n427 ;
 wire \i56/n428 ;
 wire \i56/n429 ;
 wire \i56/n43 ;
 wire \i56/n430 ;
 wire \i56/n431 ;
 wire \i56/n432 ;
 wire \i56/n433 ;
 wire \i56/n434 ;
 wire \i56/n435 ;
 wire \i56/n436 ;
 wire \i56/n437 ;
 wire \i56/n438 ;
 wire \i56/n439 ;
 wire \i56/n44 ;
 wire \i56/n440 ;
 wire \i56/n441 ;
 wire \i56/n442 ;
 wire \i56/n443 ;
 wire \i56/n444 ;
 wire \i56/n445 ;
 wire \i56/n446 ;
 wire \i56/n447 ;
 wire \i56/n448 ;
 wire \i56/n449 ;
 wire \i56/n45 ;
 wire \i56/n450 ;
 wire \i56/n451 ;
 wire \i56/n452 ;
 wire \i56/n453 ;
 wire \i56/n454 ;
 wire \i56/n455 ;
 wire \i56/n456 ;
 wire \i56/n457 ;
 wire \i56/n458 ;
 wire \i56/n459 ;
 wire \i56/n46 ;
 wire \i56/n460 ;
 wire \i56/n461 ;
 wire \i56/n462 ;
 wire \i56/n463 ;
 wire \i56/n464 ;
 wire \i56/n465 ;
 wire \i56/n466 ;
 wire \i56/n467 ;
 wire \i56/n468 ;
 wire \i56/n469 ;
 wire \i56/n47 ;
 wire \i56/n470 ;
 wire \i56/n471 ;
 wire \i56/n472 ;
 wire \i56/n473 ;
 wire \i56/n474 ;
 wire \i56/n475 ;
 wire \i56/n476 ;
 wire \i56/n477 ;
 wire \i56/n478 ;
 wire \i56/n479 ;
 wire \i56/n48 ;
 wire \i56/n480 ;
 wire \i56/n481 ;
 wire \i56/n482 ;
 wire \i56/n483 ;
 wire \i56/n484 ;
 wire \i56/n485 ;
 wire \i56/n486 ;
 wire \i56/n487 ;
 wire \i56/n488 ;
 wire \i56/n489 ;
 wire \i56/n49 ;
 wire \i56/n490 ;
 wire \i56/n491 ;
 wire \i56/n492 ;
 wire \i56/n493 ;
 wire \i56/n494 ;
 wire \i56/n495 ;
 wire \i56/n496 ;
 wire \i56/n497 ;
 wire \i56/n498 ;
 wire \i56/n499 ;
 wire \i56/n5 ;
 wire \i56/n50 ;
 wire \i56/n500 ;
 wire \i56/n501 ;
 wire \i56/n502 ;
 wire \i56/n503 ;
 wire \i56/n504 ;
 wire \i56/n505 ;
 wire \i56/n506 ;
 wire \i56/n507 ;
 wire \i56/n508 ;
 wire \i56/n509 ;
 wire \i56/n51 ;
 wire \i56/n510 ;
 wire \i56/n511 ;
 wire \i56/n512 ;
 wire \i56/n513 ;
 wire \i56/n514 ;
 wire \i56/n515 ;
 wire \i56/n516 ;
 wire \i56/n517 ;
 wire \i56/n518 ;
 wire \i56/n519 ;
 wire \i56/n52 ;
 wire \i56/n520 ;
 wire \i56/n521 ;
 wire \i56/n522 ;
 wire \i56/n523 ;
 wire \i56/n524 ;
 wire \i56/n525 ;
 wire \i56/n526 ;
 wire \i56/n527 ;
 wire \i56/n528 ;
 wire \i56/n529 ;
 wire \i56/n53 ;
 wire \i56/n530 ;
 wire \i56/n531 ;
 wire \i56/n532 ;
 wire \i56/n533 ;
 wire \i56/n534 ;
 wire \i56/n535 ;
 wire \i56/n536 ;
 wire \i56/n537 ;
 wire \i56/n538 ;
 wire \i56/n539 ;
 wire \i56/n54 ;
 wire \i56/n540 ;
 wire \i56/n541 ;
 wire \i56/n542 ;
 wire \i56/n543 ;
 wire \i56/n544 ;
 wire \i56/n545 ;
 wire \i56/n546 ;
 wire \i56/n547 ;
 wire \i56/n548 ;
 wire \i56/n549 ;
 wire \i56/n55 ;
 wire \i56/n550 ;
 wire \i56/n551 ;
 wire \i56/n552 ;
 wire \i56/n553 ;
 wire \i56/n554 ;
 wire \i56/n555 ;
 wire \i56/n556 ;
 wire \i56/n557 ;
 wire \i56/n56 ;
 wire \i56/n57 ;
 wire \i56/n58 ;
 wire \i56/n59 ;
 wire \i56/n6 ;
 wire \i56/n60 ;
 wire \i56/n61 ;
 wire \i56/n62 ;
 wire \i56/n63 ;
 wire \i56/n64 ;
 wire \i56/n65 ;
 wire \i56/n66 ;
 wire \i56/n67 ;
 wire \i56/n68 ;
 wire \i56/n69 ;
 wire \i56/n7 ;
 wire \i56/n70 ;
 wire \i56/n71 ;
 wire \i56/n72 ;
 wire \i56/n73 ;
 wire \i56/n74 ;
 wire \i56/n75 ;
 wire \i56/n76 ;
 wire \i56/n77 ;
 wire \i56/n78 ;
 wire \i56/n79 ;
 wire \i56/n8 ;
 wire \i56/n80 ;
 wire \i56/n81 ;
 wire \i56/n82 ;
 wire \i56/n83 ;
 wire \i56/n84 ;
 wire \i56/n85 ;
 wire \i56/n86 ;
 wire \i56/n87 ;
 wire \i56/n88 ;
 wire \i56/n89 ;
 wire \i56/n9 ;
 wire \i56/n90 ;
 wire \i56/n91 ;
 wire \i56/n92 ;
 wire \i56/n93 ;
 wire \i56/n94 ;
 wire \i56/n95 ;
 wire \i56/n96 ;
 wire \i56/n97 ;
 wire \i56/n98 ;
 wire \i56/n99 ;
 wire \i57/n0 ;
 wire \i57/n1 ;
 wire \i57/n10 ;
 wire \i57/n100 ;
 wire \i57/n101 ;
 wire \i57/n102 ;
 wire \i57/n103 ;
 wire \i57/n104 ;
 wire \i57/n105 ;
 wire \i57/n106 ;
 wire \i57/n107 ;
 wire \i57/n108 ;
 wire \i57/n109 ;
 wire \i57/n11 ;
 wire \i57/n110 ;
 wire \i57/n111 ;
 wire \i57/n112 ;
 wire \i57/n113 ;
 wire \i57/n114 ;
 wire \i57/n115 ;
 wire \i57/n116 ;
 wire \i57/n117 ;
 wire \i57/n118 ;
 wire \i57/n119 ;
 wire \i57/n12 ;
 wire \i57/n120 ;
 wire \i57/n121 ;
 wire \i57/n122 ;
 wire \i57/n123 ;
 wire \i57/n124 ;
 wire \i57/n125 ;
 wire \i57/n126 ;
 wire \i57/n127 ;
 wire \i57/n128 ;
 wire \i57/n129 ;
 wire \i57/n13 ;
 wire \i57/n130 ;
 wire \i57/n131 ;
 wire \i57/n132 ;
 wire \i57/n133 ;
 wire \i57/n134 ;
 wire \i57/n135 ;
 wire \i57/n136 ;
 wire \i57/n137 ;
 wire \i57/n138 ;
 wire \i57/n139 ;
 wire \i57/n14 ;
 wire \i57/n140 ;
 wire \i57/n141 ;
 wire \i57/n142 ;
 wire \i57/n143 ;
 wire \i57/n144 ;
 wire \i57/n145 ;
 wire \i57/n146 ;
 wire \i57/n147 ;
 wire \i57/n148 ;
 wire \i57/n149 ;
 wire \i57/n15 ;
 wire \i57/n150 ;
 wire \i57/n151 ;
 wire \i57/n152 ;
 wire \i57/n153 ;
 wire \i57/n154 ;
 wire \i57/n155 ;
 wire \i57/n156 ;
 wire \i57/n157 ;
 wire \i57/n158 ;
 wire \i57/n159 ;
 wire \i57/n16 ;
 wire \i57/n160 ;
 wire \i57/n161 ;
 wire \i57/n162 ;
 wire \i57/n163 ;
 wire \i57/n164 ;
 wire \i57/n165 ;
 wire \i57/n166 ;
 wire \i57/n167 ;
 wire \i57/n168 ;
 wire \i57/n169 ;
 wire \i57/n17 ;
 wire \i57/n170 ;
 wire \i57/n171 ;
 wire \i57/n172 ;
 wire \i57/n173 ;
 wire \i57/n174 ;
 wire \i57/n175 ;
 wire \i57/n176 ;
 wire \i57/n177 ;
 wire \i57/n178 ;
 wire \i57/n179 ;
 wire \i57/n18 ;
 wire \i57/n180 ;
 wire \i57/n181 ;
 wire \i57/n182 ;
 wire \i57/n183 ;
 wire \i57/n184 ;
 wire \i57/n185 ;
 wire \i57/n186 ;
 wire \i57/n187 ;
 wire \i57/n188 ;
 wire \i57/n189 ;
 wire \i57/n19 ;
 wire \i57/n190 ;
 wire \i57/n191 ;
 wire \i57/n192 ;
 wire \i57/n193 ;
 wire \i57/n194 ;
 wire \i57/n195 ;
 wire \i57/n196 ;
 wire \i57/n197 ;
 wire \i57/n198 ;
 wire \i57/n199 ;
 wire \i57/n2 ;
 wire \i57/n20 ;
 wire \i57/n200 ;
 wire \i57/n201 ;
 wire \i57/n202 ;
 wire \i57/n203 ;
 wire \i57/n204 ;
 wire \i57/n205 ;
 wire \i57/n206 ;
 wire \i57/n207 ;
 wire \i57/n208 ;
 wire \i57/n209 ;
 wire \i57/n21 ;
 wire \i57/n210 ;
 wire \i57/n211 ;
 wire \i57/n212 ;
 wire \i57/n213 ;
 wire \i57/n214 ;
 wire \i57/n215 ;
 wire \i57/n216 ;
 wire \i57/n217 ;
 wire \i57/n218 ;
 wire \i57/n219 ;
 wire \i57/n22 ;
 wire \i57/n220 ;
 wire \i57/n221 ;
 wire \i57/n222 ;
 wire \i57/n223 ;
 wire \i57/n224 ;
 wire \i57/n225 ;
 wire \i57/n226 ;
 wire \i57/n227 ;
 wire \i57/n228 ;
 wire \i57/n229 ;
 wire \i57/n23 ;
 wire \i57/n230 ;
 wire \i57/n231 ;
 wire \i57/n232 ;
 wire \i57/n233 ;
 wire \i57/n234 ;
 wire \i57/n235 ;
 wire \i57/n236 ;
 wire \i57/n237 ;
 wire \i57/n238 ;
 wire \i57/n239 ;
 wire \i57/n24 ;
 wire \i57/n240 ;
 wire \i57/n241 ;
 wire \i57/n242 ;
 wire \i57/n243 ;
 wire \i57/n244 ;
 wire \i57/n245 ;
 wire \i57/n246 ;
 wire \i57/n247 ;
 wire \i57/n248 ;
 wire \i57/n249 ;
 wire \i57/n25 ;
 wire \i57/n250 ;
 wire \i57/n251 ;
 wire \i57/n252 ;
 wire \i57/n253 ;
 wire \i57/n254 ;
 wire \i57/n255 ;
 wire \i57/n256 ;
 wire \i57/n257 ;
 wire \i57/n258 ;
 wire \i57/n259 ;
 wire \i57/n26 ;
 wire \i57/n260 ;
 wire \i57/n261 ;
 wire \i57/n262 ;
 wire \i57/n263 ;
 wire \i57/n264 ;
 wire \i57/n265 ;
 wire \i57/n266 ;
 wire \i57/n267 ;
 wire \i57/n268 ;
 wire \i57/n269 ;
 wire \i57/n27 ;
 wire \i57/n270 ;
 wire \i57/n271 ;
 wire \i57/n272 ;
 wire \i57/n273 ;
 wire \i57/n274 ;
 wire \i57/n275 ;
 wire \i57/n276 ;
 wire \i57/n277 ;
 wire \i57/n278 ;
 wire \i57/n279 ;
 wire \i57/n28 ;
 wire \i57/n280 ;
 wire \i57/n281 ;
 wire \i57/n282 ;
 wire \i57/n283 ;
 wire \i57/n284 ;
 wire \i57/n285 ;
 wire \i57/n286 ;
 wire \i57/n287 ;
 wire \i57/n288 ;
 wire \i57/n289 ;
 wire \i57/n29 ;
 wire \i57/n290 ;
 wire \i57/n291 ;
 wire \i57/n292 ;
 wire \i57/n293 ;
 wire \i57/n294 ;
 wire \i57/n295 ;
 wire \i57/n296 ;
 wire \i57/n297 ;
 wire \i57/n298 ;
 wire \i57/n299 ;
 wire \i57/n3 ;
 wire \i57/n30 ;
 wire \i57/n300 ;
 wire \i57/n301 ;
 wire \i57/n302 ;
 wire \i57/n303 ;
 wire \i57/n304 ;
 wire \i57/n305 ;
 wire \i57/n306 ;
 wire \i57/n307 ;
 wire \i57/n308 ;
 wire \i57/n309 ;
 wire \i57/n31 ;
 wire \i57/n310 ;
 wire \i57/n311 ;
 wire \i57/n312 ;
 wire \i57/n313 ;
 wire \i57/n314 ;
 wire \i57/n315 ;
 wire \i57/n316 ;
 wire \i57/n317 ;
 wire \i57/n318 ;
 wire \i57/n319 ;
 wire \i57/n32 ;
 wire \i57/n320 ;
 wire \i57/n321 ;
 wire \i57/n322 ;
 wire \i57/n323 ;
 wire \i57/n324 ;
 wire \i57/n325 ;
 wire \i57/n326 ;
 wire \i57/n327 ;
 wire \i57/n328 ;
 wire \i57/n329 ;
 wire \i57/n33 ;
 wire \i57/n330 ;
 wire \i57/n331 ;
 wire \i57/n332 ;
 wire \i57/n333 ;
 wire \i57/n334 ;
 wire \i57/n335 ;
 wire \i57/n336 ;
 wire \i57/n337 ;
 wire \i57/n338 ;
 wire \i57/n339 ;
 wire \i57/n34 ;
 wire \i57/n340 ;
 wire \i57/n341 ;
 wire \i57/n342 ;
 wire \i57/n343 ;
 wire \i57/n344 ;
 wire \i57/n345 ;
 wire \i57/n346 ;
 wire \i57/n347 ;
 wire \i57/n348 ;
 wire \i57/n349 ;
 wire \i57/n35 ;
 wire \i57/n350 ;
 wire \i57/n351 ;
 wire \i57/n352 ;
 wire \i57/n353 ;
 wire \i57/n354 ;
 wire \i57/n355 ;
 wire \i57/n356 ;
 wire \i57/n357 ;
 wire \i57/n358 ;
 wire \i57/n359 ;
 wire \i57/n36 ;
 wire \i57/n360 ;
 wire \i57/n361 ;
 wire \i57/n362 ;
 wire \i57/n363 ;
 wire \i57/n364 ;
 wire \i57/n365 ;
 wire \i57/n366 ;
 wire \i57/n367 ;
 wire \i57/n368 ;
 wire \i57/n369 ;
 wire \i57/n37 ;
 wire \i57/n370 ;
 wire \i57/n371 ;
 wire \i57/n372 ;
 wire \i57/n373 ;
 wire \i57/n374 ;
 wire \i57/n375 ;
 wire \i57/n376 ;
 wire \i57/n377 ;
 wire \i57/n378 ;
 wire \i57/n379 ;
 wire \i57/n38 ;
 wire \i57/n380 ;
 wire \i57/n381 ;
 wire \i57/n382 ;
 wire \i57/n383 ;
 wire \i57/n384 ;
 wire \i57/n385 ;
 wire \i57/n386 ;
 wire \i57/n387 ;
 wire \i57/n388 ;
 wire \i57/n389 ;
 wire \i57/n39 ;
 wire \i57/n390 ;
 wire \i57/n391 ;
 wire \i57/n392 ;
 wire \i57/n393 ;
 wire \i57/n394 ;
 wire \i57/n395 ;
 wire \i57/n396 ;
 wire \i57/n397 ;
 wire \i57/n398 ;
 wire \i57/n399 ;
 wire \i57/n4 ;
 wire \i57/n40 ;
 wire \i57/n400 ;
 wire \i57/n401 ;
 wire \i57/n402 ;
 wire \i57/n403 ;
 wire \i57/n404 ;
 wire \i57/n405 ;
 wire \i57/n406 ;
 wire \i57/n407 ;
 wire \i57/n408 ;
 wire \i57/n409 ;
 wire \i57/n41 ;
 wire \i57/n410 ;
 wire \i57/n411 ;
 wire \i57/n412 ;
 wire \i57/n413 ;
 wire \i57/n414 ;
 wire \i57/n415 ;
 wire \i57/n416 ;
 wire \i57/n417 ;
 wire \i57/n418 ;
 wire \i57/n419 ;
 wire \i57/n42 ;
 wire \i57/n420 ;
 wire \i57/n421 ;
 wire \i57/n422 ;
 wire \i57/n423 ;
 wire \i57/n424 ;
 wire \i57/n425 ;
 wire \i57/n426 ;
 wire \i57/n427 ;
 wire \i57/n428 ;
 wire \i57/n429 ;
 wire \i57/n43 ;
 wire \i57/n430 ;
 wire \i57/n431 ;
 wire \i57/n432 ;
 wire \i57/n433 ;
 wire \i57/n434 ;
 wire \i57/n435 ;
 wire \i57/n436 ;
 wire \i57/n437 ;
 wire \i57/n438 ;
 wire \i57/n439 ;
 wire \i57/n44 ;
 wire \i57/n440 ;
 wire \i57/n441 ;
 wire \i57/n442 ;
 wire \i57/n443 ;
 wire \i57/n444 ;
 wire \i57/n445 ;
 wire \i57/n446 ;
 wire \i57/n447 ;
 wire \i57/n448 ;
 wire \i57/n449 ;
 wire \i57/n45 ;
 wire \i57/n450 ;
 wire \i57/n451 ;
 wire \i57/n452 ;
 wire \i57/n453 ;
 wire \i57/n454 ;
 wire \i57/n455 ;
 wire \i57/n456 ;
 wire \i57/n457 ;
 wire \i57/n458 ;
 wire \i57/n459 ;
 wire \i57/n46 ;
 wire \i57/n460 ;
 wire \i57/n461 ;
 wire \i57/n462 ;
 wire \i57/n463 ;
 wire \i57/n464 ;
 wire \i57/n465 ;
 wire \i57/n466 ;
 wire \i57/n467 ;
 wire \i57/n468 ;
 wire \i57/n469 ;
 wire \i57/n47 ;
 wire \i57/n470 ;
 wire \i57/n471 ;
 wire \i57/n472 ;
 wire \i57/n473 ;
 wire \i57/n474 ;
 wire \i57/n475 ;
 wire \i57/n476 ;
 wire \i57/n477 ;
 wire \i57/n478 ;
 wire \i57/n479 ;
 wire \i57/n48 ;
 wire \i57/n480 ;
 wire \i57/n481 ;
 wire \i57/n482 ;
 wire \i57/n483 ;
 wire \i57/n484 ;
 wire \i57/n485 ;
 wire \i57/n486 ;
 wire \i57/n487 ;
 wire \i57/n488 ;
 wire \i57/n489 ;
 wire \i57/n49 ;
 wire \i57/n490 ;
 wire \i57/n491 ;
 wire \i57/n492 ;
 wire \i57/n493 ;
 wire \i57/n494 ;
 wire \i57/n495 ;
 wire \i57/n496 ;
 wire \i57/n497 ;
 wire \i57/n498 ;
 wire \i57/n499 ;
 wire \i57/n5 ;
 wire \i57/n50 ;
 wire \i57/n500 ;
 wire \i57/n501 ;
 wire \i57/n502 ;
 wire \i57/n503 ;
 wire \i57/n504 ;
 wire \i57/n505 ;
 wire \i57/n506 ;
 wire \i57/n507 ;
 wire \i57/n508 ;
 wire \i57/n509 ;
 wire \i57/n51 ;
 wire \i57/n510 ;
 wire \i57/n511 ;
 wire \i57/n512 ;
 wire \i57/n513 ;
 wire \i57/n514 ;
 wire \i57/n515 ;
 wire \i57/n516 ;
 wire \i57/n517 ;
 wire \i57/n518 ;
 wire \i57/n519 ;
 wire \i57/n52 ;
 wire \i57/n520 ;
 wire \i57/n521 ;
 wire \i57/n522 ;
 wire \i57/n523 ;
 wire \i57/n524 ;
 wire \i57/n525 ;
 wire \i57/n526 ;
 wire \i57/n527 ;
 wire \i57/n528 ;
 wire \i57/n529 ;
 wire \i57/n53 ;
 wire \i57/n530 ;
 wire \i57/n531 ;
 wire \i57/n532 ;
 wire \i57/n533 ;
 wire \i57/n534 ;
 wire \i57/n535 ;
 wire \i57/n536 ;
 wire \i57/n537 ;
 wire \i57/n538 ;
 wire \i57/n539 ;
 wire \i57/n54 ;
 wire \i57/n540 ;
 wire \i57/n541 ;
 wire \i57/n542 ;
 wire \i57/n543 ;
 wire \i57/n544 ;
 wire \i57/n545 ;
 wire \i57/n546 ;
 wire \i57/n547 ;
 wire \i57/n548 ;
 wire \i57/n549 ;
 wire \i57/n55 ;
 wire \i57/n550 ;
 wire \i57/n551 ;
 wire \i57/n552 ;
 wire \i57/n553 ;
 wire \i57/n554 ;
 wire \i57/n555 ;
 wire \i57/n556 ;
 wire \i57/n557 ;
 wire \i57/n558 ;
 wire \i57/n56 ;
 wire \i57/n57 ;
 wire \i57/n58 ;
 wire \i57/n59 ;
 wire \i57/n6 ;
 wire \i57/n60 ;
 wire \i57/n61 ;
 wire \i57/n62 ;
 wire \i57/n63 ;
 wire \i57/n64 ;
 wire \i57/n65 ;
 wire \i57/n66 ;
 wire \i57/n67 ;
 wire \i57/n68 ;
 wire \i57/n69 ;
 wire \i57/n7 ;
 wire \i57/n70 ;
 wire \i57/n71 ;
 wire \i57/n72 ;
 wire \i57/n73 ;
 wire \i57/n74 ;
 wire \i57/n75 ;
 wire \i57/n76 ;
 wire \i57/n77 ;
 wire \i57/n78 ;
 wire \i57/n79 ;
 wire \i57/n8 ;
 wire \i57/n80 ;
 wire \i57/n81 ;
 wire \i57/n82 ;
 wire \i57/n83 ;
 wire \i57/n84 ;
 wire \i57/n85 ;
 wire \i57/n86 ;
 wire \i57/n87 ;
 wire \i57/n88 ;
 wire \i57/n89 ;
 wire \i57/n9 ;
 wire \i57/n90 ;
 wire \i57/n91 ;
 wire \i57/n92 ;
 wire \i57/n93 ;
 wire \i57/n94 ;
 wire \i57/n95 ;
 wire \i57/n96 ;
 wire \i57/n97 ;
 wire \i57/n98 ;
 wire \i57/n99 ;
 wire \i58/n0 ;
 wire \i58/n1 ;
 wire \i58/n10 ;
 wire \i58/n100 ;
 wire \i58/n101 ;
 wire \i58/n102 ;
 wire \i58/n103 ;
 wire \i58/n104 ;
 wire \i58/n105 ;
 wire \i58/n106 ;
 wire \i58/n107 ;
 wire \i58/n108 ;
 wire \i58/n109 ;
 wire \i58/n11 ;
 wire \i58/n110 ;
 wire \i58/n111 ;
 wire \i58/n112 ;
 wire \i58/n113 ;
 wire \i58/n114 ;
 wire \i58/n115 ;
 wire \i58/n116 ;
 wire \i58/n117 ;
 wire \i58/n118 ;
 wire \i58/n119 ;
 wire \i58/n12 ;
 wire \i58/n120 ;
 wire \i58/n121 ;
 wire \i58/n122 ;
 wire \i58/n123 ;
 wire \i58/n124 ;
 wire \i58/n125 ;
 wire \i58/n126 ;
 wire \i58/n127 ;
 wire \i58/n128 ;
 wire \i58/n129 ;
 wire \i58/n13 ;
 wire \i58/n130 ;
 wire \i58/n131 ;
 wire \i58/n132 ;
 wire \i58/n133 ;
 wire \i58/n134 ;
 wire \i58/n135 ;
 wire \i58/n136 ;
 wire \i58/n137 ;
 wire \i58/n138 ;
 wire \i58/n139 ;
 wire \i58/n14 ;
 wire \i58/n140 ;
 wire \i58/n141 ;
 wire \i58/n142 ;
 wire \i58/n143 ;
 wire \i58/n144 ;
 wire \i58/n145 ;
 wire \i58/n146 ;
 wire \i58/n147 ;
 wire \i58/n148 ;
 wire \i58/n149 ;
 wire \i58/n15 ;
 wire \i58/n150 ;
 wire \i58/n151 ;
 wire \i58/n152 ;
 wire \i58/n153 ;
 wire \i58/n154 ;
 wire \i58/n155 ;
 wire \i58/n156 ;
 wire \i58/n157 ;
 wire \i58/n158 ;
 wire \i58/n159 ;
 wire \i58/n16 ;
 wire \i58/n160 ;
 wire \i58/n161 ;
 wire \i58/n162 ;
 wire \i58/n163 ;
 wire \i58/n164 ;
 wire \i58/n165 ;
 wire \i58/n166 ;
 wire \i58/n167 ;
 wire \i58/n168 ;
 wire \i58/n169 ;
 wire \i58/n17 ;
 wire \i58/n170 ;
 wire \i58/n171 ;
 wire \i58/n172 ;
 wire \i58/n173 ;
 wire \i58/n174 ;
 wire \i58/n175 ;
 wire \i58/n176 ;
 wire \i58/n177 ;
 wire \i58/n178 ;
 wire \i58/n179 ;
 wire \i58/n18 ;
 wire \i58/n180 ;
 wire \i58/n181 ;
 wire \i58/n182 ;
 wire \i58/n183 ;
 wire \i58/n184 ;
 wire \i58/n185 ;
 wire \i58/n186 ;
 wire \i58/n187 ;
 wire \i58/n188 ;
 wire \i58/n189 ;
 wire \i58/n19 ;
 wire \i58/n190 ;
 wire \i58/n191 ;
 wire \i58/n192 ;
 wire \i58/n193 ;
 wire \i58/n194 ;
 wire \i58/n195 ;
 wire \i58/n196 ;
 wire \i58/n197 ;
 wire \i58/n198 ;
 wire \i58/n199 ;
 wire \i58/n2 ;
 wire \i58/n20 ;
 wire \i58/n200 ;
 wire \i58/n201 ;
 wire \i58/n202 ;
 wire \i58/n203 ;
 wire \i58/n204 ;
 wire \i58/n205 ;
 wire \i58/n206 ;
 wire \i58/n207 ;
 wire \i58/n208 ;
 wire \i58/n209 ;
 wire \i58/n21 ;
 wire \i58/n210 ;
 wire \i58/n211 ;
 wire \i58/n212 ;
 wire \i58/n213 ;
 wire \i58/n214 ;
 wire \i58/n215 ;
 wire \i58/n216 ;
 wire \i58/n217 ;
 wire \i58/n218 ;
 wire \i58/n219 ;
 wire \i58/n22 ;
 wire \i58/n220 ;
 wire \i58/n221 ;
 wire \i58/n222 ;
 wire \i58/n223 ;
 wire \i58/n224 ;
 wire \i58/n225 ;
 wire \i58/n226 ;
 wire \i58/n227 ;
 wire \i58/n228 ;
 wire \i58/n229 ;
 wire \i58/n23 ;
 wire \i58/n230 ;
 wire \i58/n231 ;
 wire \i58/n232 ;
 wire \i58/n233 ;
 wire \i58/n234 ;
 wire \i58/n235 ;
 wire \i58/n236 ;
 wire \i58/n237 ;
 wire \i58/n238 ;
 wire \i58/n239 ;
 wire \i58/n24 ;
 wire \i58/n240 ;
 wire \i58/n241 ;
 wire \i58/n242 ;
 wire \i58/n243 ;
 wire \i58/n244 ;
 wire \i58/n245 ;
 wire \i58/n246 ;
 wire \i58/n247 ;
 wire \i58/n248 ;
 wire \i58/n249 ;
 wire \i58/n25 ;
 wire \i58/n250 ;
 wire \i58/n251 ;
 wire \i58/n252 ;
 wire \i58/n253 ;
 wire \i58/n254 ;
 wire \i58/n255 ;
 wire \i58/n256 ;
 wire \i58/n257 ;
 wire \i58/n258 ;
 wire \i58/n259 ;
 wire \i58/n26 ;
 wire \i58/n260 ;
 wire \i58/n261 ;
 wire \i58/n262 ;
 wire \i58/n263 ;
 wire \i58/n264 ;
 wire \i58/n265 ;
 wire \i58/n266 ;
 wire \i58/n267 ;
 wire \i58/n268 ;
 wire \i58/n269 ;
 wire \i58/n27 ;
 wire \i58/n270 ;
 wire \i58/n271 ;
 wire \i58/n272 ;
 wire \i58/n273 ;
 wire \i58/n274 ;
 wire \i58/n275 ;
 wire \i58/n276 ;
 wire \i58/n277 ;
 wire \i58/n278 ;
 wire \i58/n279 ;
 wire \i58/n28 ;
 wire \i58/n280 ;
 wire \i58/n281 ;
 wire \i58/n282 ;
 wire \i58/n283 ;
 wire \i58/n284 ;
 wire \i58/n285 ;
 wire \i58/n286 ;
 wire \i58/n287 ;
 wire \i58/n288 ;
 wire \i58/n289 ;
 wire \i58/n29 ;
 wire \i58/n290 ;
 wire \i58/n291 ;
 wire \i58/n292 ;
 wire \i58/n293 ;
 wire \i58/n294 ;
 wire \i58/n295 ;
 wire \i58/n296 ;
 wire \i58/n297 ;
 wire \i58/n298 ;
 wire \i58/n299 ;
 wire \i58/n3 ;
 wire \i58/n30 ;
 wire \i58/n300 ;
 wire \i58/n301 ;
 wire \i58/n302 ;
 wire \i58/n303 ;
 wire \i58/n304 ;
 wire \i58/n305 ;
 wire \i58/n306 ;
 wire \i58/n307 ;
 wire \i58/n308 ;
 wire \i58/n309 ;
 wire \i58/n31 ;
 wire \i58/n310 ;
 wire \i58/n311 ;
 wire \i58/n312 ;
 wire \i58/n313 ;
 wire \i58/n314 ;
 wire \i58/n315 ;
 wire \i58/n316 ;
 wire \i58/n317 ;
 wire \i58/n318 ;
 wire \i58/n319 ;
 wire \i58/n32 ;
 wire \i58/n320 ;
 wire \i58/n321 ;
 wire \i58/n322 ;
 wire \i58/n323 ;
 wire \i58/n324 ;
 wire \i58/n325 ;
 wire \i58/n326 ;
 wire \i58/n327 ;
 wire \i58/n328 ;
 wire \i58/n329 ;
 wire \i58/n33 ;
 wire \i58/n330 ;
 wire \i58/n331 ;
 wire \i58/n332 ;
 wire \i58/n333 ;
 wire \i58/n334 ;
 wire \i58/n335 ;
 wire \i58/n336 ;
 wire \i58/n337 ;
 wire \i58/n338 ;
 wire \i58/n339 ;
 wire \i58/n34 ;
 wire \i58/n340 ;
 wire \i58/n341 ;
 wire \i58/n342 ;
 wire \i58/n343 ;
 wire \i58/n344 ;
 wire \i58/n345 ;
 wire \i58/n346 ;
 wire \i58/n347 ;
 wire \i58/n348 ;
 wire \i58/n349 ;
 wire \i58/n35 ;
 wire \i58/n350 ;
 wire \i58/n351 ;
 wire \i58/n352 ;
 wire \i58/n353 ;
 wire \i58/n354 ;
 wire \i58/n355 ;
 wire \i58/n356 ;
 wire \i58/n357 ;
 wire \i58/n358 ;
 wire \i58/n359 ;
 wire \i58/n36 ;
 wire \i58/n360 ;
 wire \i58/n361 ;
 wire \i58/n362 ;
 wire \i58/n363 ;
 wire \i58/n364 ;
 wire \i58/n365 ;
 wire \i58/n366 ;
 wire \i58/n367 ;
 wire \i58/n368 ;
 wire \i58/n369 ;
 wire \i58/n37 ;
 wire \i58/n370 ;
 wire \i58/n371 ;
 wire \i58/n372 ;
 wire \i58/n373 ;
 wire \i58/n374 ;
 wire \i58/n375 ;
 wire \i58/n376 ;
 wire \i58/n377 ;
 wire \i58/n378 ;
 wire \i58/n379 ;
 wire \i58/n38 ;
 wire \i58/n380 ;
 wire \i58/n381 ;
 wire \i58/n382 ;
 wire \i58/n383 ;
 wire \i58/n384 ;
 wire \i58/n385 ;
 wire \i58/n386 ;
 wire \i58/n387 ;
 wire \i58/n388 ;
 wire \i58/n389 ;
 wire \i58/n39 ;
 wire \i58/n390 ;
 wire \i58/n391 ;
 wire \i58/n392 ;
 wire \i58/n393 ;
 wire \i58/n394 ;
 wire \i58/n395 ;
 wire \i58/n396 ;
 wire \i58/n397 ;
 wire \i58/n398 ;
 wire \i58/n399 ;
 wire \i58/n4 ;
 wire \i58/n40 ;
 wire \i58/n400 ;
 wire \i58/n401 ;
 wire \i58/n402 ;
 wire \i58/n403 ;
 wire \i58/n404 ;
 wire \i58/n405 ;
 wire \i58/n406 ;
 wire \i58/n407 ;
 wire \i58/n408 ;
 wire \i58/n409 ;
 wire \i58/n41 ;
 wire \i58/n410 ;
 wire \i58/n411 ;
 wire \i58/n412 ;
 wire \i58/n413 ;
 wire \i58/n414 ;
 wire \i58/n415 ;
 wire \i58/n416 ;
 wire \i58/n417 ;
 wire \i58/n418 ;
 wire \i58/n419 ;
 wire \i58/n42 ;
 wire \i58/n420 ;
 wire \i58/n421 ;
 wire \i58/n422 ;
 wire \i58/n423 ;
 wire \i58/n424 ;
 wire \i58/n425 ;
 wire \i58/n426 ;
 wire \i58/n427 ;
 wire \i58/n428 ;
 wire \i58/n429 ;
 wire \i58/n43 ;
 wire \i58/n430 ;
 wire \i58/n431 ;
 wire \i58/n432 ;
 wire \i58/n433 ;
 wire \i58/n434 ;
 wire \i58/n435 ;
 wire \i58/n436 ;
 wire \i58/n437 ;
 wire \i58/n438 ;
 wire \i58/n439 ;
 wire \i58/n44 ;
 wire \i58/n440 ;
 wire \i58/n441 ;
 wire \i58/n442 ;
 wire \i58/n443 ;
 wire \i58/n444 ;
 wire \i58/n445 ;
 wire \i58/n446 ;
 wire \i58/n447 ;
 wire \i58/n448 ;
 wire \i58/n449 ;
 wire \i58/n45 ;
 wire \i58/n450 ;
 wire \i58/n451 ;
 wire \i58/n452 ;
 wire \i58/n453 ;
 wire \i58/n454 ;
 wire \i58/n455 ;
 wire \i58/n456 ;
 wire \i58/n457 ;
 wire \i58/n458 ;
 wire \i58/n459 ;
 wire \i58/n46 ;
 wire \i58/n460 ;
 wire \i58/n461 ;
 wire \i58/n462 ;
 wire \i58/n463 ;
 wire \i58/n464 ;
 wire \i58/n465 ;
 wire \i58/n466 ;
 wire \i58/n467 ;
 wire \i58/n468 ;
 wire \i58/n469 ;
 wire \i58/n47 ;
 wire \i58/n470 ;
 wire \i58/n471 ;
 wire \i58/n472 ;
 wire \i58/n473 ;
 wire \i58/n474 ;
 wire \i58/n475 ;
 wire \i58/n476 ;
 wire \i58/n477 ;
 wire \i58/n478 ;
 wire \i58/n479 ;
 wire \i58/n48 ;
 wire \i58/n480 ;
 wire \i58/n481 ;
 wire \i58/n482 ;
 wire \i58/n483 ;
 wire \i58/n484 ;
 wire \i58/n485 ;
 wire \i58/n486 ;
 wire \i58/n487 ;
 wire \i58/n488 ;
 wire \i58/n489 ;
 wire \i58/n49 ;
 wire \i58/n490 ;
 wire \i58/n491 ;
 wire \i58/n492 ;
 wire \i58/n493 ;
 wire \i58/n494 ;
 wire \i58/n495 ;
 wire \i58/n496 ;
 wire \i58/n497 ;
 wire \i58/n498 ;
 wire \i58/n499 ;
 wire \i58/n5 ;
 wire \i58/n50 ;
 wire \i58/n500 ;
 wire \i58/n501 ;
 wire \i58/n502 ;
 wire \i58/n503 ;
 wire \i58/n504 ;
 wire \i58/n505 ;
 wire \i58/n506 ;
 wire \i58/n507 ;
 wire \i58/n508 ;
 wire \i58/n509 ;
 wire \i58/n51 ;
 wire \i58/n510 ;
 wire \i58/n511 ;
 wire \i58/n512 ;
 wire \i58/n513 ;
 wire \i58/n514 ;
 wire \i58/n515 ;
 wire \i58/n516 ;
 wire \i58/n517 ;
 wire \i58/n518 ;
 wire \i58/n519 ;
 wire \i58/n52 ;
 wire \i58/n520 ;
 wire \i58/n521 ;
 wire \i58/n522 ;
 wire \i58/n523 ;
 wire \i58/n524 ;
 wire \i58/n525 ;
 wire \i58/n526 ;
 wire \i58/n527 ;
 wire \i58/n528 ;
 wire \i58/n529 ;
 wire \i58/n53 ;
 wire \i58/n530 ;
 wire \i58/n531 ;
 wire \i58/n532 ;
 wire \i58/n533 ;
 wire \i58/n534 ;
 wire \i58/n535 ;
 wire \i58/n536 ;
 wire \i58/n537 ;
 wire \i58/n538 ;
 wire \i58/n539 ;
 wire \i58/n54 ;
 wire \i58/n540 ;
 wire \i58/n541 ;
 wire \i58/n542 ;
 wire \i58/n543 ;
 wire \i58/n544 ;
 wire \i58/n545 ;
 wire \i58/n546 ;
 wire \i58/n547 ;
 wire \i58/n548 ;
 wire \i58/n549 ;
 wire \i58/n55 ;
 wire \i58/n550 ;
 wire \i58/n551 ;
 wire \i58/n552 ;
 wire \i58/n553 ;
 wire \i58/n554 ;
 wire \i58/n555 ;
 wire \i58/n556 ;
 wire \i58/n557 ;
 wire \i58/n558 ;
 wire \i58/n56 ;
 wire \i58/n57 ;
 wire \i58/n58 ;
 wire \i58/n59 ;
 wire \i58/n6 ;
 wire \i58/n60 ;
 wire \i58/n61 ;
 wire \i58/n62 ;
 wire \i58/n63 ;
 wire \i58/n64 ;
 wire \i58/n65 ;
 wire \i58/n66 ;
 wire \i58/n67 ;
 wire \i58/n68 ;
 wire \i58/n69 ;
 wire \i58/n7 ;
 wire \i58/n70 ;
 wire \i58/n71 ;
 wire \i58/n72 ;
 wire \i58/n73 ;
 wire \i58/n74 ;
 wire \i58/n75 ;
 wire \i58/n76 ;
 wire \i58/n77 ;
 wire \i58/n78 ;
 wire \i58/n79 ;
 wire \i58/n8 ;
 wire \i58/n80 ;
 wire \i58/n81 ;
 wire \i58/n82 ;
 wire \i58/n83 ;
 wire \i58/n84 ;
 wire \i58/n85 ;
 wire \i58/n86 ;
 wire \i58/n87 ;
 wire \i58/n88 ;
 wire \i58/n89 ;
 wire \i58/n9 ;
 wire \i58/n90 ;
 wire \i58/n91 ;
 wire \i58/n92 ;
 wire \i58/n93 ;
 wire \i58/n94 ;
 wire \i58/n95 ;
 wire \i58/n96 ;
 wire \i58/n97 ;
 wire \i58/n98 ;
 wire \i58/n99 ;
 wire \i59/n0 ;
 wire \i59/n1 ;
 wire \i59/n10 ;
 wire \i59/n100 ;
 wire \i59/n101 ;
 wire \i59/n102 ;
 wire \i59/n103 ;
 wire \i59/n104 ;
 wire \i59/n105 ;
 wire \i59/n106 ;
 wire \i59/n107 ;
 wire \i59/n108 ;
 wire \i59/n109 ;
 wire \i59/n11 ;
 wire \i59/n110 ;
 wire \i59/n111 ;
 wire \i59/n112 ;
 wire \i59/n113 ;
 wire \i59/n114 ;
 wire \i59/n115 ;
 wire \i59/n116 ;
 wire \i59/n117 ;
 wire \i59/n118 ;
 wire \i59/n119 ;
 wire \i59/n12 ;
 wire \i59/n120 ;
 wire \i59/n121 ;
 wire \i59/n122 ;
 wire \i59/n123 ;
 wire \i59/n124 ;
 wire \i59/n125 ;
 wire \i59/n126 ;
 wire \i59/n127 ;
 wire \i59/n128 ;
 wire \i59/n129 ;
 wire \i59/n13 ;
 wire \i59/n130 ;
 wire \i59/n131 ;
 wire \i59/n132 ;
 wire \i59/n133 ;
 wire \i59/n134 ;
 wire \i59/n135 ;
 wire \i59/n136 ;
 wire \i59/n137 ;
 wire \i59/n138 ;
 wire \i59/n139 ;
 wire \i59/n14 ;
 wire \i59/n140 ;
 wire \i59/n141 ;
 wire \i59/n142 ;
 wire \i59/n143 ;
 wire \i59/n144 ;
 wire \i59/n145 ;
 wire \i59/n146 ;
 wire \i59/n147 ;
 wire \i59/n148 ;
 wire \i59/n149 ;
 wire \i59/n15 ;
 wire \i59/n150 ;
 wire \i59/n151 ;
 wire \i59/n152 ;
 wire \i59/n153 ;
 wire \i59/n154 ;
 wire \i59/n155 ;
 wire \i59/n156 ;
 wire \i59/n157 ;
 wire \i59/n158 ;
 wire \i59/n159 ;
 wire \i59/n16 ;
 wire \i59/n160 ;
 wire \i59/n161 ;
 wire \i59/n162 ;
 wire \i59/n163 ;
 wire \i59/n164 ;
 wire \i59/n165 ;
 wire \i59/n166 ;
 wire \i59/n167 ;
 wire \i59/n168 ;
 wire \i59/n169 ;
 wire \i59/n17 ;
 wire \i59/n170 ;
 wire \i59/n171 ;
 wire \i59/n172 ;
 wire \i59/n173 ;
 wire \i59/n174 ;
 wire \i59/n175 ;
 wire \i59/n176 ;
 wire \i59/n177 ;
 wire \i59/n178 ;
 wire \i59/n179 ;
 wire \i59/n18 ;
 wire \i59/n180 ;
 wire \i59/n181 ;
 wire \i59/n182 ;
 wire \i59/n183 ;
 wire \i59/n184 ;
 wire \i59/n185 ;
 wire \i59/n186 ;
 wire \i59/n187 ;
 wire \i59/n188 ;
 wire \i59/n189 ;
 wire \i59/n19 ;
 wire \i59/n190 ;
 wire \i59/n191 ;
 wire \i59/n192 ;
 wire \i59/n193 ;
 wire \i59/n194 ;
 wire \i59/n195 ;
 wire \i59/n196 ;
 wire \i59/n197 ;
 wire \i59/n198 ;
 wire \i59/n199 ;
 wire \i59/n2 ;
 wire \i59/n20 ;
 wire \i59/n200 ;
 wire \i59/n201 ;
 wire \i59/n202 ;
 wire \i59/n203 ;
 wire \i59/n204 ;
 wire \i59/n205 ;
 wire \i59/n206 ;
 wire \i59/n207 ;
 wire \i59/n208 ;
 wire \i59/n209 ;
 wire \i59/n21 ;
 wire \i59/n210 ;
 wire \i59/n211 ;
 wire \i59/n212 ;
 wire \i59/n213 ;
 wire \i59/n214 ;
 wire \i59/n215 ;
 wire \i59/n216 ;
 wire \i59/n217 ;
 wire \i59/n218 ;
 wire \i59/n219 ;
 wire \i59/n22 ;
 wire \i59/n220 ;
 wire \i59/n221 ;
 wire \i59/n222 ;
 wire \i59/n223 ;
 wire \i59/n224 ;
 wire \i59/n225 ;
 wire \i59/n226 ;
 wire \i59/n227 ;
 wire \i59/n228 ;
 wire \i59/n229 ;
 wire \i59/n23 ;
 wire \i59/n230 ;
 wire \i59/n231 ;
 wire \i59/n232 ;
 wire \i59/n233 ;
 wire \i59/n234 ;
 wire \i59/n235 ;
 wire \i59/n236 ;
 wire \i59/n237 ;
 wire \i59/n238 ;
 wire \i59/n239 ;
 wire \i59/n24 ;
 wire \i59/n240 ;
 wire \i59/n241 ;
 wire \i59/n242 ;
 wire \i59/n243 ;
 wire \i59/n244 ;
 wire \i59/n245 ;
 wire \i59/n246 ;
 wire \i59/n247 ;
 wire \i59/n248 ;
 wire \i59/n249 ;
 wire \i59/n25 ;
 wire \i59/n250 ;
 wire \i59/n251 ;
 wire \i59/n252 ;
 wire \i59/n253 ;
 wire \i59/n254 ;
 wire \i59/n255 ;
 wire \i59/n256 ;
 wire \i59/n257 ;
 wire \i59/n258 ;
 wire \i59/n259 ;
 wire \i59/n26 ;
 wire \i59/n260 ;
 wire \i59/n261 ;
 wire \i59/n262 ;
 wire \i59/n263 ;
 wire \i59/n264 ;
 wire \i59/n265 ;
 wire \i59/n266 ;
 wire \i59/n267 ;
 wire \i59/n268 ;
 wire \i59/n269 ;
 wire \i59/n27 ;
 wire \i59/n270 ;
 wire \i59/n271 ;
 wire \i59/n272 ;
 wire \i59/n273 ;
 wire \i59/n274 ;
 wire \i59/n275 ;
 wire \i59/n276 ;
 wire \i59/n277 ;
 wire \i59/n278 ;
 wire \i59/n279 ;
 wire \i59/n28 ;
 wire \i59/n280 ;
 wire \i59/n281 ;
 wire \i59/n282 ;
 wire \i59/n283 ;
 wire \i59/n284 ;
 wire \i59/n285 ;
 wire \i59/n286 ;
 wire \i59/n287 ;
 wire \i59/n288 ;
 wire \i59/n289 ;
 wire \i59/n29 ;
 wire \i59/n290 ;
 wire \i59/n291 ;
 wire \i59/n292 ;
 wire \i59/n293 ;
 wire \i59/n294 ;
 wire \i59/n295 ;
 wire \i59/n296 ;
 wire \i59/n297 ;
 wire \i59/n298 ;
 wire \i59/n299 ;
 wire \i59/n3 ;
 wire \i59/n30 ;
 wire \i59/n300 ;
 wire \i59/n301 ;
 wire \i59/n302 ;
 wire \i59/n303 ;
 wire \i59/n304 ;
 wire \i59/n305 ;
 wire \i59/n306 ;
 wire \i59/n307 ;
 wire \i59/n308 ;
 wire \i59/n309 ;
 wire \i59/n31 ;
 wire \i59/n310 ;
 wire \i59/n311 ;
 wire \i59/n312 ;
 wire \i59/n313 ;
 wire \i59/n314 ;
 wire \i59/n315 ;
 wire \i59/n316 ;
 wire \i59/n317 ;
 wire \i59/n318 ;
 wire \i59/n319 ;
 wire \i59/n32 ;
 wire \i59/n320 ;
 wire \i59/n321 ;
 wire \i59/n322 ;
 wire \i59/n323 ;
 wire \i59/n324 ;
 wire \i59/n325 ;
 wire \i59/n326 ;
 wire \i59/n327 ;
 wire \i59/n328 ;
 wire \i59/n329 ;
 wire \i59/n33 ;
 wire \i59/n330 ;
 wire \i59/n331 ;
 wire \i59/n332 ;
 wire \i59/n333 ;
 wire \i59/n334 ;
 wire \i59/n335 ;
 wire \i59/n336 ;
 wire \i59/n337 ;
 wire \i59/n338 ;
 wire \i59/n339 ;
 wire \i59/n34 ;
 wire \i59/n340 ;
 wire \i59/n341 ;
 wire \i59/n342 ;
 wire \i59/n343 ;
 wire \i59/n344 ;
 wire \i59/n345 ;
 wire \i59/n346 ;
 wire \i59/n347 ;
 wire \i59/n348 ;
 wire \i59/n349 ;
 wire \i59/n35 ;
 wire \i59/n350 ;
 wire \i59/n351 ;
 wire \i59/n352 ;
 wire \i59/n353 ;
 wire \i59/n354 ;
 wire \i59/n355 ;
 wire \i59/n356 ;
 wire \i59/n357 ;
 wire \i59/n358 ;
 wire \i59/n359 ;
 wire \i59/n36 ;
 wire \i59/n360 ;
 wire \i59/n361 ;
 wire \i59/n362 ;
 wire \i59/n363 ;
 wire \i59/n364 ;
 wire \i59/n365 ;
 wire \i59/n366 ;
 wire \i59/n367 ;
 wire \i59/n368 ;
 wire \i59/n369 ;
 wire \i59/n37 ;
 wire \i59/n370 ;
 wire \i59/n371 ;
 wire \i59/n372 ;
 wire \i59/n373 ;
 wire \i59/n374 ;
 wire \i59/n375 ;
 wire \i59/n376 ;
 wire \i59/n377 ;
 wire \i59/n378 ;
 wire \i59/n379 ;
 wire \i59/n38 ;
 wire \i59/n380 ;
 wire \i59/n381 ;
 wire \i59/n382 ;
 wire \i59/n383 ;
 wire \i59/n384 ;
 wire \i59/n385 ;
 wire \i59/n386 ;
 wire \i59/n387 ;
 wire \i59/n388 ;
 wire \i59/n389 ;
 wire \i59/n39 ;
 wire \i59/n390 ;
 wire \i59/n391 ;
 wire \i59/n392 ;
 wire \i59/n393 ;
 wire \i59/n394 ;
 wire \i59/n395 ;
 wire \i59/n396 ;
 wire \i59/n397 ;
 wire \i59/n398 ;
 wire \i59/n399 ;
 wire \i59/n4 ;
 wire \i59/n40 ;
 wire \i59/n400 ;
 wire \i59/n401 ;
 wire \i59/n402 ;
 wire \i59/n403 ;
 wire \i59/n404 ;
 wire \i59/n405 ;
 wire \i59/n406 ;
 wire \i59/n407 ;
 wire \i59/n408 ;
 wire \i59/n409 ;
 wire \i59/n41 ;
 wire \i59/n410 ;
 wire \i59/n411 ;
 wire \i59/n412 ;
 wire \i59/n413 ;
 wire \i59/n414 ;
 wire \i59/n415 ;
 wire \i59/n416 ;
 wire \i59/n417 ;
 wire \i59/n418 ;
 wire \i59/n419 ;
 wire \i59/n42 ;
 wire \i59/n420 ;
 wire \i59/n421 ;
 wire \i59/n422 ;
 wire \i59/n423 ;
 wire \i59/n424 ;
 wire \i59/n425 ;
 wire \i59/n426 ;
 wire \i59/n427 ;
 wire \i59/n428 ;
 wire \i59/n429 ;
 wire \i59/n43 ;
 wire \i59/n430 ;
 wire \i59/n431 ;
 wire \i59/n432 ;
 wire \i59/n433 ;
 wire \i59/n434 ;
 wire \i59/n435 ;
 wire \i59/n436 ;
 wire \i59/n437 ;
 wire \i59/n438 ;
 wire \i59/n439 ;
 wire \i59/n44 ;
 wire \i59/n440 ;
 wire \i59/n441 ;
 wire \i59/n442 ;
 wire \i59/n443 ;
 wire \i59/n444 ;
 wire \i59/n445 ;
 wire \i59/n446 ;
 wire \i59/n447 ;
 wire \i59/n448 ;
 wire \i59/n449 ;
 wire \i59/n45 ;
 wire \i59/n450 ;
 wire \i59/n451 ;
 wire \i59/n452 ;
 wire \i59/n453 ;
 wire \i59/n454 ;
 wire \i59/n455 ;
 wire \i59/n456 ;
 wire \i59/n457 ;
 wire \i59/n458 ;
 wire \i59/n459 ;
 wire \i59/n46 ;
 wire \i59/n460 ;
 wire \i59/n461 ;
 wire \i59/n462 ;
 wire \i59/n463 ;
 wire \i59/n464 ;
 wire \i59/n465 ;
 wire \i59/n466 ;
 wire \i59/n467 ;
 wire \i59/n468 ;
 wire \i59/n469 ;
 wire \i59/n47 ;
 wire \i59/n470 ;
 wire \i59/n471 ;
 wire \i59/n472 ;
 wire \i59/n473 ;
 wire \i59/n474 ;
 wire \i59/n475 ;
 wire \i59/n476 ;
 wire \i59/n477 ;
 wire \i59/n478 ;
 wire \i59/n479 ;
 wire \i59/n48 ;
 wire \i59/n480 ;
 wire \i59/n481 ;
 wire \i59/n482 ;
 wire \i59/n483 ;
 wire \i59/n484 ;
 wire \i59/n485 ;
 wire \i59/n486 ;
 wire \i59/n487 ;
 wire \i59/n488 ;
 wire \i59/n489 ;
 wire \i59/n49 ;
 wire \i59/n490 ;
 wire \i59/n491 ;
 wire \i59/n492 ;
 wire \i59/n493 ;
 wire \i59/n494 ;
 wire \i59/n495 ;
 wire \i59/n496 ;
 wire \i59/n497 ;
 wire \i59/n498 ;
 wire \i59/n499 ;
 wire \i59/n5 ;
 wire \i59/n50 ;
 wire \i59/n500 ;
 wire \i59/n501 ;
 wire \i59/n502 ;
 wire \i59/n503 ;
 wire \i59/n504 ;
 wire \i59/n505 ;
 wire \i59/n506 ;
 wire \i59/n507 ;
 wire \i59/n508 ;
 wire \i59/n509 ;
 wire \i59/n51 ;
 wire \i59/n510 ;
 wire \i59/n511 ;
 wire \i59/n512 ;
 wire \i59/n513 ;
 wire \i59/n514 ;
 wire \i59/n515 ;
 wire \i59/n516 ;
 wire \i59/n517 ;
 wire \i59/n518 ;
 wire \i59/n519 ;
 wire \i59/n52 ;
 wire \i59/n520 ;
 wire \i59/n521 ;
 wire \i59/n522 ;
 wire \i59/n523 ;
 wire \i59/n524 ;
 wire \i59/n525 ;
 wire \i59/n526 ;
 wire \i59/n527 ;
 wire \i59/n528 ;
 wire \i59/n529 ;
 wire \i59/n53 ;
 wire \i59/n530 ;
 wire \i59/n531 ;
 wire \i59/n532 ;
 wire \i59/n533 ;
 wire \i59/n534 ;
 wire \i59/n535 ;
 wire \i59/n536 ;
 wire \i59/n537 ;
 wire \i59/n538 ;
 wire \i59/n539 ;
 wire \i59/n54 ;
 wire \i59/n540 ;
 wire \i59/n541 ;
 wire \i59/n542 ;
 wire \i59/n543 ;
 wire \i59/n544 ;
 wire \i59/n545 ;
 wire \i59/n546 ;
 wire \i59/n547 ;
 wire \i59/n548 ;
 wire \i59/n549 ;
 wire \i59/n55 ;
 wire \i59/n550 ;
 wire \i59/n551 ;
 wire \i59/n552 ;
 wire \i59/n553 ;
 wire \i59/n554 ;
 wire \i59/n555 ;
 wire \i59/n56 ;
 wire \i59/n57 ;
 wire \i59/n58 ;
 wire \i59/n59 ;
 wire \i59/n6 ;
 wire \i59/n60 ;
 wire \i59/n61 ;
 wire \i59/n62 ;
 wire \i59/n63 ;
 wire \i59/n64 ;
 wire \i59/n65 ;
 wire \i59/n66 ;
 wire \i59/n67 ;
 wire \i59/n68 ;
 wire \i59/n69 ;
 wire \i59/n7 ;
 wire \i59/n70 ;
 wire \i59/n71 ;
 wire \i59/n72 ;
 wire \i59/n73 ;
 wire \i59/n74 ;
 wire \i59/n75 ;
 wire \i59/n76 ;
 wire \i59/n77 ;
 wire \i59/n78 ;
 wire \i59/n79 ;
 wire \i59/n8 ;
 wire \i59/n80 ;
 wire \i59/n81 ;
 wire \i59/n82 ;
 wire \i59/n83 ;
 wire \i59/n84 ;
 wire \i59/n85 ;
 wire \i59/n86 ;
 wire \i59/n87 ;
 wire \i59/n88 ;
 wire \i59/n89 ;
 wire \i59/n9 ;
 wire \i59/n90 ;
 wire \i59/n91 ;
 wire \i59/n92 ;
 wire \i59/n93 ;
 wire \i59/n94 ;
 wire \i59/n95 ;
 wire \i59/n96 ;
 wire \i59/n97 ;
 wire \i59/n98 ;
 wire \i59/n99 ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire [3:0] \i43/i45/n0 ;
 wire [3:0] \i43/i45/n1 ;
 wire [31:0] \i43/n0 ;
 wire [31:0] \i43/n2 ;
 wire [127:0] n0;
 wire [3:0] n1;
 wire [7:0] n10;
 wire [7:0] n11;
 wire [7:0] n12;
 wire [7:0] n13;
 wire [7:0] n14;
 wire [7:0] n15;
 wire [7:0] n16;
 wire [7:0] n17;
 wire [7:0] n18;
 wire [7:0] n19;
 wire [7:0] n2;
 wire [7:0] n20;
 wire [7:0] n21;
 wire [7:0] n22;
 wire [7:0] n23;
 wire [7:0] n24;
 wire [7:0] n25;
 wire [7:0] n26;
 wire [7:0] n27;
 wire [7:0] n28;
 wire [7:0] n29;
 wire [7:0] n3;
 wire [7:0] n30;
 wire [7:0] n31;
 wire [7:0] n32;
 wire [7:0] n33;
 wire [31:0] n34;
 wire [31:0] n35;
 wire [31:0] n36;
 wire [31:0] n37;
 wire [7:0] n4;
 wire [7:0] n5;
 wire [7:0] n6;
 wire [7:0] n7;
 wire [7:0] n8;
 wire [7:0] n9;

 INVx2_ASAP7_75t_SL i0 (.A(net129),
    .Y(n38));
 INVx2_ASAP7_75t_SL i1 (.A(n32[7]),
    .Y(n84));
 INVxp67_ASAP7_75t_SL i10 (.A(n22[7]),
    .Y(n93));
 SDFHx4_ASAP7_75t_SL i100 (.CLK(clk),
    .D(n392),
    .QN(n27[6]),
    .SE(n1229),
    .SI(n1090));
 XNOR2xp5_ASAP7_75t_SL i1000 (.A(n0[117]),
    .B(n37[21]),
    .Y(n417));
 XNOR2xp5_ASAP7_75t_SL i1001 (.A(n34[19]),
    .B(n0[19]),
    .Y(n416));
 XNOR2xp5_ASAP7_75t_SL i1002 (.A(n0[126]),
    .B(n37[30]),
    .Y(n415));
 XNOR2xp5_ASAP7_75t_SL i1003 (.A(n0[68]),
    .B(n36[4]),
    .Y(n414));
 XNOR2xp5_ASAP7_75t_SL i1004 (.A(n0[3]),
    .B(n34[3]),
    .Y(n413));
 XNOR2xp5_ASAP7_75t_SL i1005 (.A(n0[67]),
    .B(n36[3]),
    .Y(n412));
 XNOR2xp5_ASAP7_75t_SL i1006 (.A(n0[116]),
    .B(n37[20]),
    .Y(n411));
 XNOR2xp5_ASAP7_75t_SL i1007 (.A(n0[66]),
    .B(n36[2]),
    .Y(n410));
 XNOR2xp5_ASAP7_75t_SL i1008 (.A(n0[65]),
    .B(n36[1]),
    .Y(n409));
 XNOR2xp5_ASAP7_75t_SL i1009 (.A(n0[115]),
    .B(n37[19]),
    .Y(n408));
 SDFHx4_ASAP7_75t_SL i101 (.CLK(clk),
    .D(n396),
    .QN(n27[7]),
    .SE(n1229),
    .SI(n1124));
 XNOR2xp5_ASAP7_75t_SL i1010 (.A(n0[64]),
    .B(n36[0]),
    .Y(n407));
 XNOR2xp5_ASAP7_75t_SL i1011 (.A(n0[125]),
    .B(n37[29]),
    .Y(n406));
 XNOR2xp5_ASAP7_75t_SL i1012 (.A(n0[103]),
    .B(n37[7]),
    .Y(n405));
 XNOR2xp5_ASAP7_75t_SL i1013 (.A(n0[113]),
    .B(n37[17]),
    .Y(n404));
 XNOR2xp5_ASAP7_75t_SL i1014 (.A(n0[102]),
    .B(n37[6]),
    .Y(n403));
 XNOR2xp5_ASAP7_75t_SL i1015 (.A(n0[101]),
    .B(n37[5]),
    .Y(n402));
 XNOR2xp5_ASAP7_75t_SL i1016 (.A(n0[55]),
    .B(n35[23]),
    .Y(n401));
 XNOR2xp5_ASAP7_75t_SL i1017 (.A(n34[4]),
    .B(n0[4]),
    .Y(n400));
 XNOR2xp5_ASAP7_75t_SL i1018 (.A(n0[112]),
    .B(n37[16]),
    .Y(n399));
 XNOR2xp5_ASAP7_75t_SL i1019 (.A(n0[100]),
    .B(n37[4]),
    .Y(n398));
 SDFHx4_ASAP7_75t_SL i102 (.CLK(clk),
    .D(n399),
    .QN(n25[0]),
    .SE(n1229),
    .SI(n1035));
 XNOR2xp5_ASAP7_75t_SL i1020 (.A(n0[99]),
    .B(n37[3]),
    .Y(n397));
 XNOR2xp5_ASAP7_75t_SL i1021 (.A(n34[31]),
    .B(n0[31]),
    .Y(n396));
 XNOR2xp5_ASAP7_75t_SL i1022 (.A(n0[124]),
    .B(n37[28]),
    .Y(n395));
 XNOR2xp5_ASAP7_75t_SL i1023 (.A(n0[98]),
    .B(n37[2]),
    .Y(n394));
 XNOR2xp5_ASAP7_75t_SL i1024 (.A(n0[97]),
    .B(n37[1]),
    .Y(n393));
 XNOR2xp5_ASAP7_75t_SL i1025 (.A(n34[30]),
    .B(n0[30]),
    .Y(n392));
 XNOR2xp5_ASAP7_75t_SL i1026 (.A(n0[96]),
    .B(n37[0]),
    .Y(n391));
 XNOR2xp5_ASAP7_75t_SL i1027 (.A(n34[15]),
    .B(n0[15]),
    .Y(n390));
 XNOR2xp5_ASAP7_75t_SL i1028 (.A(n34[14]),
    .B(n0[14]),
    .Y(n388));
 XNOR2xp5_ASAP7_75t_SL i1029 (.A(n34[29]),
    .B(n0[29]),
    .Y(n387));
 SDFHx4_ASAP7_75t_SL i103 (.CLK(clk),
    .D(n404),
    .QN(n25[1]),
    .SE(n1229),
    .SI(n1083));
 XNOR2xp5_ASAP7_75t_SL i1030 (.A(n0[123]),
    .B(n37[27]),
    .Y(n386));
 XNOR2xp5_ASAP7_75t_SL i1031 (.A(n34[13]),
    .B(n0[13]),
    .Y(n385));
 XNOR2xp5_ASAP7_75t_SL i1032 (.A(n34[12]),
    .B(n0[12]),
    .Y(n384));
 XNOR2xp5_ASAP7_75t_SL i1033 (.A(n34[28]),
    .B(n0[28]),
    .Y(n383));
 XNOR2xp5_ASAP7_75t_SL i1034 (.A(n0[11]),
    .B(n34[11]),
    .Y(n382));
 XNOR2xp5_ASAP7_75t_SL i1035 (.A(n34[10]),
    .B(n0[10]),
    .Y(n381));
 XNOR2xp5_ASAP7_75t_SL i1036 (.A(n0[85]),
    .B(n36[21]),
    .Y(n380));
 XNOR2xp5_ASAP7_75t_SL i1037 (.A(n34[9]),
    .B(n0[9]),
    .Y(n379));
 XNOR2xp5_ASAP7_75t_SL i1038 (.A(n0[122]),
    .B(n37[26]),
    .Y(n378));
 XNOR2xp5_ASAP7_75t_SL i1039 (.A(n0[27]),
    .B(n34[27]),
    .Y(n377));
 SDFHx4_ASAP7_75t_SL i104 (.CLK(clk),
    .D(n408),
    .QN(n25[3]),
    .SE(n1229),
    .SI(n1082));
 XNOR2xp5_ASAP7_75t_SL i1040 (.A(n0[8]),
    .B(n34[8]),
    .Y(n376));
 XNOR2xp5_ASAP7_75t_SL i1041 (.A(n0[47]),
    .B(n35[15]),
    .Y(n375));
 XNOR2xp5_ASAP7_75t_SL i1042 (.A(n0[46]),
    .B(n35[14]),
    .Y(n374));
 XNOR2xp5_ASAP7_75t_SL i1043 (.A(n34[26]),
    .B(n0[26]),
    .Y(n373));
 XNOR2xp5_ASAP7_75t_SL i1044 (.A(n0[45]),
    .B(n35[13]),
    .Y(n372));
 XNOR2xp5_ASAP7_75t_SL i1045 (.A(n0[44]),
    .B(n35[12]),
    .Y(n371));
 XNOR2xp5_ASAP7_75t_SL i1046 (.A(n0[121]),
    .B(n37[25]),
    .Y(n370));
 XNOR2xp5_ASAP7_75t_SL i1047 (.A(n34[25]),
    .B(n0[25]),
    .Y(n369));
 XNOR2xp5_ASAP7_75t_SL i1048 (.A(n0[43]),
    .B(n35[11]),
    .Y(n368));
 XNOR2xp5_ASAP7_75t_SL i1049 (.A(n0[90]),
    .B(n36[26]),
    .Y(n367));
 SDFHx4_ASAP7_75t_SL i105 (.CLK(clk),
    .D(n411),
    .QN(n25[4]),
    .SE(n1229),
    .SI(n1079));
 XNOR2xp5_ASAP7_75t_SL i1050 (.A(n0[42]),
    .B(n35[10]),
    .Y(n366));
 XNOR2xp5_ASAP7_75t_SL i1051 (.A(n0[41]),
    .B(n35[9]),
    .Y(n365));
 XNOR2xp5_ASAP7_75t_SL i1052 (.A(n0[111]),
    .B(n37[15]),
    .Y(n364));
 XNOR2xp5_ASAP7_75t_SL i1053 (.A(n0[60]),
    .B(n35[28]),
    .Y(n363));
 XNOR2xp5_ASAP7_75t_SL i1054 (.A(n0[72]),
    .B(n36[8]),
    .Y(n362));
 XNOR2xp5_ASAP7_75t_SL i1055 (.A(n0[73]),
    .B(n36[9]),
    .Y(n361));
 XNOR2xp5_ASAP7_75t_SL i1056 (.A(n0[61]),
    .B(n35[29]),
    .Y(n360));
 XNOR2xp5_ASAP7_75t_SL i1057 (.A(n0[74]),
    .B(n36[10]),
    .Y(n359));
 XNOR2xp5_ASAP7_75t_SL i1058 (.A(n0[75]),
    .B(n36[11]),
    .Y(n358));
 XNOR2xp5_ASAP7_75t_SL i1059 (.A(n0[76]),
    .B(n36[12]),
    .Y(n357));
 SDFHx4_ASAP7_75t_SL i106 (.CLK(clk),
    .D(n417),
    .QN(n25[5]),
    .SE(n1229),
    .SI(n1074));
 XNOR2xp5_ASAP7_75t_SL i1060 (.A(n0[62]),
    .B(n35[30]),
    .Y(n356));
 XNOR2xp5_ASAP7_75t_SL i1061 (.A(n0[77]),
    .B(n36[13]),
    .Y(n355));
 XNOR2xp5_ASAP7_75t_SL i1062 (.A(n0[86]),
    .B(n36[22]),
    .Y(n354));
 XNOR2xp5_ASAP7_75t_SL i1063 (.A(n0[78]),
    .B(n36[14]),
    .Y(n353));
 XNOR2xp5_ASAP7_75t_SL i1064 (.A(n0[120]),
    .B(n37[24]),
    .Y(n352));
 XNOR2xp5_ASAP7_75t_SL i1065 (.A(n0[63]),
    .B(n35[31]),
    .Y(n351));
 XNOR2xp5_ASAP7_75t_SL i1066 (.A(n0[79]),
    .B(n36[15]),
    .Y(n350));
 XNOR2xp5_ASAP7_75t_SL i1067 (.A(n0[40]),
    .B(n35[8]),
    .Y(n349));
 OAI22xp5_ASAP7_75t_SL i1068 (.A1(n259),
    .A2(n6[1]),
    .B1(n35[9]),
    .B2(n166),
    .Y(n582));
 OAI22xp5_ASAP7_75t_SL i1069 (.A1(n273),
    .A2(n2[6]),
    .B1(n37[14]),
    .B2(n122),
    .Y(n348));
 SDFHx4_ASAP7_75t_SL i107 (.CLK(clk),
    .D(n471),
    .QN(n25[6]),
    .SE(n1229),
    .SI(n1072));
 OAI22xp5_ASAP7_75t_SL i1070 (.A1(n62),
    .A2(n24[0]),
    .B1(n34[24]),
    .B2(n130),
    .Y(n579));
 AOI22xp5_ASAP7_75t_R i1071 (.A1(n8[2]),
    .A2(n198),
    .B1(n113),
    .B2(n30[2]),
    .Y(n347));
 OAI22xp5_ASAP7_75t_SL i1072 (.A1(n46),
    .A2(n22[3]),
    .B1(n37[20]),
    .B2(n1166),
    .Y(n346));
 AOI22xp5_ASAP7_75t_SL i1073 (.A1(n2[5]),
    .A2(n184),
    .B1(n181),
    .B2(n2[4]),
    .Y(n578));
 OAI22xp5_ASAP7_75t_SL i1074 (.A1(n286),
    .A2(n18[2]),
    .B1(n35[26]),
    .B2(n189),
    .Y(n575));
 OAI22xp5_ASAP7_75t_SL i1075 (.A1(n116),
    .A2(n28[3]),
    .B1(n6[3]),
    .B2(n182),
    .Y(n345));
 OAI22xp5_ASAP7_75t_SL i1076 (.A1(n253),
    .A2(n2[3]),
    .B1(n37[11]),
    .B2(n123),
    .Y(n573));
 OAI22xp5_ASAP7_75t_SL i1077 (.A1(n44),
    .A2(n22[1]),
    .B1(n37[25]),
    .B2(n176),
    .Y(n571));
 OAI22xp5_ASAP7_75t_SL i1078 (.A1(n280),
    .A2(n18[7]),
    .B1(n35[15]),
    .B2(n1160),
    .Y(n569));
 OAI22xp33_ASAP7_75t_SL i1079 (.A1(n112),
    .A2(n30[3]),
    .B1(n8[3]),
    .B2(n165),
    .Y(n344));
 SDFHx4_ASAP7_75t_SL i108 (.CLK(clk),
    .D(n423),
    .QN(n25[7]),
    .SE(n1229),
    .SI(n1139));
 OAI22xp5_ASAP7_75t_SL i1080 (.A1(n16[1]),
    .A2(n186),
    .B1(n28[2]),
    .B2(n191),
    .Y(n567));
 OAI22xp5_ASAP7_75t_SL i1081 (.A1(n275),
    .A2(n2[1]),
    .B1(n37[9]),
    .B2(n192),
    .Y(n565));
 OAI22xp5_ASAP7_75t_SL i1082 (.A1(n248),
    .A2(n18[1]),
    .B1(n35[25]),
    .B2(n228),
    .Y(n563));
 OAI22xp5_ASAP7_75t_SL i1083 (.A1(n75),
    .A2(n4[1]),
    .B1(n34[9]),
    .B2(n164),
    .Y(n561));
 AOI22xp5_ASAP7_75t_SL i1084 (.A1(n157),
    .A2(n37[21]),
    .B1(n45),
    .B2(n32[5]),
    .Y(n343));
 OAI22xp5_ASAP7_75t_SL i1085 (.A1(n251),
    .A2(n2[0]),
    .B1(n37[8]),
    .B2(n194),
    .Y(n559));
 OAI22xp5_ASAP7_75t_SL i1086 (.A1(n289),
    .A2(n30[5]),
    .B1(n36[6]),
    .B2(n1164),
    .Y(n342));
 OAI22xp5_ASAP7_75t_SL i1087 (.A1(n40),
    .A2(n22[6]),
    .B1(n37[30]),
    .B2(n152),
    .Y(n341));
 OAI22xp5_ASAP7_75t_SL i1088 (.A1(n14[6]),
    .A2(n1157),
    .B1(n100),
    .B2(n14[7]),
    .Y(n557));
 OAI22xp5_ASAP7_75t_R i1089 (.A1(n63),
    .A2(n24[6]),
    .B1(n34[23]),
    .B2(n92),
    .Y(n340));
 SDFHx4_ASAP7_75t_SL i109 (.CLK(clk),
    .D(n426),
    .QN(n23[0]),
    .SE(n1229),
    .SI(n1032));
 OAI22xp5_ASAP7_75t_SL i1090 (.A1(n49),
    .A2(n2[2]),
    .B1(n37[10]),
    .B2(n187),
    .Y(n555));
 AOI22xp5_ASAP7_75t_SL i1091 (.A1(n195),
    .A2(n34[22]),
    .B1(n64),
    .B2(n24[5]),
    .Y(n339));
 AOI22xp5_ASAP7_75t_SL i1092 (.A1(n26[6]),
    .A2(n190),
    .B1(n14[5]),
    .B2(n91),
    .Y(n338));
 OAI22xp5_ASAP7_75t_SL i1093 (.A1(n134),
    .A2(n30[6]),
    .B1(n8[6]),
    .B2(n135),
    .Y(n337));
 OAI22xp5_ASAP7_75t_SL i1094 (.A1(n70),
    .A2(n24[7]),
    .B1(n34[15]),
    .B2(n1156),
    .Y(n553));
 OAI22xp5_ASAP7_75t_SL i1095 (.A1(n65),
    .A2(n26[5]),
    .B1(n140),
    .B2(n34[21]),
    .Y(n551));
 OAI22xp5_ASAP7_75t_SL i1096 (.A1(n241),
    .A2(n30[7]),
    .B1(n36[7]),
    .B2(n86),
    .Y(n336));
 OAI22xp5_ASAP7_75t_SL i1097 (.A1(n66),
    .A2(n24[3]),
    .B1(n34[20]),
    .B2(n1222),
    .Y(n335));
 OAI22xp5_ASAP7_75t_SL i1098 (.A1(n288),
    .A2(n12[1]),
    .B1(n37[1]),
    .B2(n177),
    .Y(n334));
 OAI22xp5_ASAP7_75t_SL i1099 (.A1(n14[3]),
    .A2(n101),
    .B1(n14[4]),
    .B2(n102),
    .Y(n333));
 INVxp33_ASAP7_75t_SL i11 (.A(n22[5]),
    .Y(n94));
 SDFHx4_ASAP7_75t_SL i110 (.CLK(clk),
    .D(n465),
    .QN(n23[1]),
    .SE(n1229),
    .SI(n1065));
 OAI22xp5_ASAP7_75t_SL i1100 (.A1(n67),
    .A2(n26[3]),
    .B1(n34[19]),
    .B2(n1227),
    .Y(n332));
 AOI22xp5_ASAP7_75t_SL i1101 (.A1(n32[6]),
    .A2(n105),
    .B1(n12[5]),
    .B2(n85),
    .Y(n331));
 AOI22xp5_ASAP7_75t_SL i1102 (.A1(n2[2]),
    .A2(n131),
    .B1(n32[2]),
    .B2(n187),
    .Y(n330));
 AOI22xp5_ASAP7_75t_SL i1103 (.A1(n94),
    .A2(n37[22]),
    .B1(n267),
    .B2(n22[5]),
    .Y(n329));
 OAI22xp5_ASAP7_75t_SL i1104 (.A1(n264),
    .A2(n18[0]),
    .B1(n35[24]),
    .B2(n133),
    .Y(n548));
 OAI22xp5_ASAP7_75t_SL i1105 (.A1(n69),
    .A2(n26[0]),
    .B1(n34[16]),
    .B2(n136),
    .Y(n546));
 AOI22xp5_ASAP7_75t_SL i1106 (.A1(n6[0]),
    .A2(n146),
    .B1(n169),
    .B2(n28[0]),
    .Y(n328));
 AOI22xp5_ASAP7_75t_SL i1107 (.A1(n20[5]),
    .A2(n162),
    .B1(n143),
    .B2(n20[4]),
    .Y(n327));
 OAI22xp5_ASAP7_75t_R i1108 (.A1(n272),
    .A2(n22[6]),
    .B1(n37[23]),
    .B2(n152),
    .Y(n326));
 AOI22xp5_ASAP7_75t_SL i1109 (.A1(n144),
    .A2(n35[22]),
    .B1(n254),
    .B2(n18[5]),
    .Y(n325));
 SDFHx4_ASAP7_75t_SL i111 (.CLK(clk),
    .D(n431),
    .QN(n23[2]),
    .SE(n1229),
    .SI(n1138));
 AOI22xp5_ASAP7_75t_SL i1110 (.A1(n200),
    .A2(n28[6]),
    .B1(n16[5]),
    .B2(n1220),
    .Y(n324));
 OAI22xp5_ASAP7_75t_SL i1111 (.A1(n53),
    .A2(n8[4]),
    .B1(n36[28]),
    .B2(n111),
    .Y(n323));
 AOI22xp33_ASAP7_75t_SL i1112 (.A1(n18[2]),
    .A2(n156),
    .B1(n189),
    .B2(n16[2]),
    .Y(n322));
 OAI22xp5_ASAP7_75t_SL i1113 (.A1(n12[6]),
    .A2(n103),
    .B1(n104),
    .B2(n12[7]),
    .Y(n544));
 OAI22xp5_ASAP7_75t_SL i1114 (.A1(n243),
    .A2(n28[3]),
    .B1(n35[19]),
    .B2(n182),
    .Y(n321));
 XOR2xp5_ASAP7_75t_SL i1115 (.A(n18[1]),
    .B(n35[18]),
    .Y(n320));
 OAI22xp5_ASAP7_75t_SL i1116 (.A1(n166),
    .A2(n16[2]),
    .B1(n6[1]),
    .B2(n156),
    .Y(n541));
 OAI22xp5_ASAP7_75t_SL i1117 (.A1(n10[6]),
    .A2(n108),
    .B1(n171),
    .B2(n10[7]),
    .Y(n539));
 OAI22xp5_ASAP7_75t_SL i1118 (.A1(n54),
    .A2(n20[2]),
    .B1(n36[26]),
    .B2(n168),
    .Y(n537));
 OAI22xp5_ASAP7_75t_R i1119 (.A1(n261),
    .A2(n20[6]),
    .B1(n36[23]),
    .B2(n96),
    .Y(n319));
 SDFHx4_ASAP7_75t_SL i112 (.CLK(clk),
    .D(n436),
    .QN(n23[3]),
    .SE(n1229),
    .SI(n1061));
 AOI22xp5_ASAP7_75t_SL i1120 (.A1(n30[6]),
    .A2(n199),
    .B1(n10[5]),
    .B2(n135),
    .Y(n318));
 OAI22xp5_ASAP7_75t_SL i1121 (.A1(n118),
    .A2(n26[6]),
    .B1(n4[6]),
    .B2(n91),
    .Y(n535));
 OAI22xp5_ASAP7_75t_SL i1122 (.A1(n233),
    .A2(n20[1]),
    .B1(n36[18]),
    .B2(n142),
    .Y(n317));
 OAI22xp33_ASAP7_75t_SL i1123 (.A1(n155),
    .A2(n14[6]),
    .B1(n4[5]),
    .B2(n100),
    .Y(n316));
 OAI22xp5_ASAP7_75t_SL i1124 (.A1(n242),
    .A2(n16[3]),
    .B1(n35[3]),
    .B2(n99),
    .Y(n315));
 AOI22xp5_ASAP7_75t_SL i1125 (.A1(n35[1]),
    .A2(n191),
    .B1(n285),
    .B2(n16[1]),
    .Y(n314));
 OAI22xp5_ASAP7_75t_SL i1126 (.A1(n79),
    .A2(n26[4]),
    .B1(n34[4]),
    .B2(n161),
    .Y(n313));
 XOR2xp5_ASAP7_75t_SL i1127 (.A(n28[1]),
    .B(n35[2]),
    .Y(n312));
 OAI22xp5_ASAP7_75t_SL i1128 (.A1(n55),
    .A2(n20[1]),
    .B1(n36[25]),
    .B2(n142),
    .Y(n531));
 OAI22xp5_ASAP7_75t_SL i1129 (.A1(n269),
    .A2(n20[3]),
    .B1(n36[20]),
    .B2(n1159),
    .Y(n311));
 SDFHx4_ASAP7_75t_SL i113 (.CLK(clk),
    .D(n438),
    .QN(n23[4]),
    .SE(n1229),
    .SI(n1058));
 OAI22xp5_ASAP7_75t_SL i1130 (.A1(n10[3]),
    .A2(n196),
    .B1(n10[4]),
    .B2(n1158),
    .Y(n310));
 AOI22xp5_ASAP7_75t_R i1131 (.A1(n4[2]),
    .A2(n163),
    .B1(n183),
    .B2(n26[2]),
    .Y(n309));
 OAI22xp5_ASAP7_75t_SL i1132 (.A1(n80),
    .A2(n14[3]),
    .B1(n34[3]),
    .B2(n102),
    .Y(n308));
 OAI22xp5_ASAP7_75t_SL i1133 (.A1(n164),
    .A2(n14[2]),
    .B1(n4[1]),
    .B2(n141),
    .Y(n529));
 OAI22xp5_ASAP7_75t_SL i1134 (.A1(n244),
    .A2(n30[3]),
    .B1(n36[19]),
    .B2(n165),
    .Y(n307));
 OAI22xp5_ASAP7_75t_SL i1135 (.A1(n10[2]),
    .A2(n168),
    .B1(n20[2]),
    .B2(n145),
    .Y(n306));
 OAI22xp5_ASAP7_75t_SL i1136 (.A1(n281),
    .A2(n20[0]),
    .B1(n36[24]),
    .B2(n97),
    .Y(n527));
 OAI22xp5_ASAP7_75t_SL i1137 (.A1(n10[1]),
    .A2(n198),
    .B1(n109),
    .B2(n30[2]),
    .Y(n525));
 AOI22xp5_ASAP7_75t_SL i1138 (.A1(n6[2]),
    .A2(n186),
    .B1(n148),
    .B2(n28[2]),
    .Y(n305));
 AOI22xp5_ASAP7_75t_SL i1139 (.A1(n132),
    .A2(n34[0]),
    .B1(n83),
    .B2(n14[0]),
    .Y(n523));
 SDFHx4_ASAP7_75t_SL i114 (.CLK(clk),
    .D(n380),
    .QN(n23[5]),
    .SE(n1229),
    .SI(n1052));
 OAI22xp5_ASAP7_75t_SL i1140 (.A1(n167),
    .A2(n28[6]),
    .B1(n1220),
    .B2(n6[6]),
    .Y(n521));
 OAI22xp5_ASAP7_75t_SL i1141 (.A1(n82),
    .A2(n14[1]),
    .B1(n34[1]),
    .B2(n151),
    .Y(n304));
 XOR2xp5_ASAP7_75t_SL i1142 (.A(n28[7]),
    .B(n35[7]),
    .Y(n303));
 OAI22xp5_ASAP7_75t_SL i1143 (.A1(n81),
    .A2(n26[1]),
    .B1(n34[2]),
    .B2(n174),
    .Y(n302));
 OAI22xp5_ASAP7_75t_SL i1144 (.A1(n14[1]),
    .A2(n163),
    .B1(n26[2]),
    .B2(n151),
    .Y(n519));
 OAI22xp5_ASAP7_75t_SL i1145 (.A1(n240),
    .A2(n28[5]),
    .B1(n35[6]),
    .B2(n188),
    .Y(n301));
 OAI22xp33_ASAP7_75t_SL i1146 (.A1(n170),
    .A2(n16[6]),
    .B1(n185),
    .B2(n6[5]),
    .Y(n300));
 OAI22xp5_ASAP7_75t_SL i1147 (.A1(n252),
    .A2(n30[0]),
    .B1(n36[16]),
    .B2(n88),
    .Y(n517));
 AOI22xp5_ASAP7_75t_SL i1148 (.A1(n36[17]),
    .A2(n159),
    .B1(n250),
    .B2(n30[1]),
    .Y(n299));
 OAI22xp5_ASAP7_75t_SL i1149 (.A1(n287),
    .A2(n16[5]),
    .B1(n35[5]),
    .B2(n200),
    .Y(n298));
 SDFHx4_ASAP7_75t_SL i115 (.CLK(clk),
    .D(n354),
    .QN(n23[6]),
    .SE(n1229),
    .SI(n1051));
 AOI22xp5_ASAP7_75t_SL i1150 (.A1(n20[0]),
    .A2(n180),
    .B1(n10[0]),
    .B2(n97),
    .Y(n297));
 AOI22xp5_ASAP7_75t_SL i1151 (.A1(n35[4]),
    .A2(n154),
    .B1(n279),
    .B2(n28[4]),
    .Y(n296));
 AOI22xp5_ASAP7_75t_L i1152 (.A1(n37[31]),
    .A2(n121),
    .B1(n2[7]),
    .B2(n39),
    .Y(n515));
 OAI22xp5_ASAP7_75t_SL i1153 (.A1(n138),
    .A2(n26[0]),
    .B1(n4[0]),
    .B2(n136),
    .Y(n295));
 OAI22xp5_ASAP7_75t_SL i1154 (.A1(n263),
    .A2(n28[5]),
    .B1(n188),
    .B2(n35[21]),
    .Y(n513));
 OAI22xp5_ASAP7_75t_SL i1155 (.A1(n122),
    .A2(n12[6]),
    .B1(n2[6]),
    .B2(n104),
    .Y(n512));
 AOI22x1_ASAP7_75t_SL i1156 (.A1(n186),
    .A2(n18[2]),
    .B1(n189),
    .B2(n28[2]),
    .Y(n511));
 AO22x2_ASAP7_75t_SL i1157 (.A1(n20[0]),
    .A2(n88),
    .B1(n30[0]),
    .B2(n97),
    .Y(n509));
 OAI22x1_ASAP7_75t_SL i1158 (.A1(n116),
    .A2(n16[3]),
    .B1(n99),
    .B2(n6[3]),
    .Y(n507));
 OAI22x1_ASAP7_75t_SL i1159 (.A1(n112),
    .A2(n10[3]),
    .B1(n8[3]),
    .B2(n1158),
    .Y(n504));
 SDFHx4_ASAP7_75t_SL i116 (.CLK(clk),
    .D(n444),
    .QN(n23[7]),
    .SE(n1229),
    .SI(n1135));
 OAI22xp5_ASAP7_75t_SL i1160 (.A1(n32[6]),
    .A2(n152),
    .B1(n85),
    .B2(n22[6]),
    .Y(n503));
 AO22x1_ASAP7_75t_SL i1161 (.A1(n8[5]),
    .A2(n199),
    .B1(n139),
    .B2(n10[5]),
    .Y(n501));
 OAI22x1_ASAP7_75t_SL i1162 (.A1(n148),
    .A2(n16[2]),
    .B1(n6[2]),
    .B2(n156),
    .Y(n500));
 OAI22x1_ASAP7_75t_SL i1163 (.A1(n149),
    .A2(n10[0]),
    .B1(n180),
    .B2(n8[0]),
    .Y(n498));
 AOI22xp5_ASAP7_75t_SL i1164 (.A1(n1164),
    .A2(n20[5]),
    .B1(n143),
    .B2(n30[5]),
    .Y(n495));
 OAI22xp5_ASAP7_75t_SL i1165 (.A1(n134),
    .A2(n10[6]),
    .B1(n8[6]),
    .B2(n171),
    .Y(n494));
 OAI22x1_ASAP7_75t_SL i1166 (.A1(n113),
    .A2(n10[2]),
    .B1(n8[2]),
    .B2(n145),
    .Y(n493));
 OAI22x1_ASAP7_75t_SL i1167 (.A1(n184),
    .A2(n32[4]),
    .B1(n2[4]),
    .B2(n197),
    .Y(n491));
 OAI22x1_ASAP7_75t_SL i1168 (.A1(n16[0]),
    .A2(n169),
    .B1(n6[0]),
    .B2(n173),
    .Y(n489));
 OAI22x1_ASAP7_75t_SL i1169 (.A1(n228),
    .A2(n28[1]),
    .B1(n18[1]),
    .B2(n175),
    .Y(n487));
 SDFHx4_ASAP7_75t_SL i117 (.CLK(clk),
    .D(n446),
    .QN(n21[0]),
    .SE(n1229),
    .SI(n1134));
 AOI22x1_ASAP7_75t_SL i1170 (.A1(n157),
    .A2(n22[5]),
    .B1(n94),
    .B2(n32[5]),
    .Y(n484));
 OAI22x1_ASAP7_75t_SL i1171 (.A1(n28[0]),
    .A2(n133),
    .B1(n18[0]),
    .B2(n146),
    .Y(n483));
 OAI22x1_ASAP7_75t_SL i1172 (.A1(n121),
    .A2(n12[7]),
    .B1(n2[7]),
    .B2(n103),
    .Y(n481));
 OA22x2_ASAP7_75t_SL i1173 (.A1(n28[7]),
    .A2(n1160),
    .B1(n89),
    .B2(n18[7]),
    .Y(n478));
 OA22x2_ASAP7_75t_SL i1174 (.A1(n10[7]),
    .A2(n95),
    .B1(n108),
    .B2(n20[7]),
    .Y(n476));
 OA22x2_ASAP7_75t_SL i1175 (.A1(n121),
    .A2(n32[7]),
    .B1(n84),
    .B2(n2[7]),
    .Y(n475));
 OA22x2_ASAP7_75t_SL i1176 (.A1(n12[7]),
    .A2(n93),
    .B1(n103),
    .B2(n22[7]),
    .Y(n474));
 AND2x2_ASAP7_75t_SL i1177 (.A(net129),
    .B(net130),
    .Y(n294));
 INVxp67_ASAP7_75t_SL i1178 (.A(n292),
    .Y(n293));
 NOR2xp33_ASAP7_75t_SL i1179 (.A(n1[1]),
    .B(n1[0]),
    .Y(n292));
 SDFHx4_ASAP7_75t_SL i118 (.CLK(clk),
    .D(n447),
    .QN(n21[2]),
    .SE(n1229),
    .SI(n1133));
 INVx1_ASAP7_75t_SL i1180 (.A(n35[16]),
    .Y(n291));
 INVx1_ASAP7_75t_SL i1181 (.A(n16[1]),
    .Y(n191));
 INVx1_ASAP7_75t_SL i1182 (.A(n35[29]),
    .Y(n290));
 INVx1_ASAP7_75t_SL i1183 (.A(n36[6]),
    .Y(n289));
 INVx1_ASAP7_75t_SL i1184 (.A(n1[0]),
    .Y(n172));
 INVx1_ASAP7_75t_SL i1185 (.A(n37[1]),
    .Y(n288));
 INVx1_ASAP7_75t_SL i1186 (.A(n35[5]),
    .Y(n287));
 INVx1_ASAP7_75t_SL i1187 (.A(n35[26]),
    .Y(n286));
 INVx1_ASAP7_75t_SL i1188 (.A(n35[1]),
    .Y(n285));
 INVx3_ASAP7_75t_SL i1189 (.A(n22[1]),
    .Y(n176));
 SDFHx4_ASAP7_75t_SL i119 (.CLK(clk),
    .D(n430),
    .QN(n21[3]),
    .SE(n1229),
    .SI(n1123));
 INVx1_ASAP7_75t_SL i1190 (.A(n37[0]),
    .Y(n284));
 INVx1_ASAP7_75t_SL i1191 (.A(n36[12]),
    .Y(n283));
 INVx1_ASAP7_75t_SL i1192 (.A(n36[9]),
    .Y(n282));
 INVx3_ASAP7_75t_SL i1193 (.A(n14[0]),
    .Y(n132));
 INVx1_ASAP7_75t_SL i1194 (.A(n36[24]),
    .Y(n281));
 INVx1_ASAP7_75t_SL i1195 (.A(n35[15]),
    .Y(n280));
 INVx1_ASAP7_75t_SL i1196 (.A(n6[5]),
    .Y(n170));
 INVx2_ASAP7_75t_SL i1197 (.A(n18[5]),
    .Y(n144));
 INVx3_ASAP7_75t_SL i1198 (.A(n8[6]),
    .Y(n134));
 INVx1_ASAP7_75t_SL i1199 (.A(n28[3]),
    .Y(n182));
 INVx2_ASAP7_75t_SL i12 (.A(n20[7]),
    .Y(n95));
 SDFHx4_ASAP7_75t_SL i120 (.CLK(clk),
    .D(n448),
    .QN(n21[4]),
    .SE(n1229),
    .SI(n1122));
 INVx3_ASAP7_75t_SL i1200 (.A(n18[4]),
    .Y(n178));
 INVx3_ASAP7_75t_SL i1201 (.A(n32[4]),
    .Y(n197));
 INVx3_ASAP7_75t_SL i1202 (.A(n18[2]),
    .Y(n189));
 INVx4_ASAP7_75t_SL i1203 (.A(n4[2]),
    .Y(n183));
 INVx3_ASAP7_75t_SL i1204 (.A(n8[0]),
    .Y(n149));
 INVx3_ASAP7_75t_SL i1205 (.A(n32[1]),
    .Y(n147));
 INVx3_ASAP7_75t_SL i1206 (.A(n30[6]),
    .Y(n135));
 INVx1_ASAP7_75t_SL i1207 (.A(n35[4]),
    .Y(n279));
 INVx1_ASAP7_75t_SL i1208 (.A(n36[0]),
    .Y(n278));
 INVx1_ASAP7_75t_SL i1209 (.A(n1152),
    .Y(n277));
 SDFHx4_ASAP7_75t_SL i121 (.CLK(clk),
    .D(n449),
    .QN(n21[5]),
    .SE(n1229),
    .SI(n1048));
 INVx1_ASAP7_75t_SL i1210 (.A(n36[22]),
    .Y(n276));
 INVx1_ASAP7_75t_SL i1211 (.A(n37[9]),
    .Y(n275));
 INVx1_ASAP7_75t_SL i1212 (.A(n36[13]),
    .Y(n274));
 INVx1_ASAP7_75t_SL i1213 (.A(n37[14]),
    .Y(n273));
 INVx1_ASAP7_75t_SL i1214 (.A(n37[23]),
    .Y(n272));
 INVx1_ASAP7_75t_SL i1215 (.A(n35[14]),
    .Y(n271));
 INVx1_ASAP7_75t_SL i1216 (.A(n1154),
    .Y(n270));
 INVx1_ASAP7_75t_SL i1217 (.A(n36[20]),
    .Y(n269));
 INVx3_ASAP7_75t_SL i1218 (.A(n24[0]),
    .Y(n130));
 INVx1_ASAP7_75t_SL i1219 (.A(n37[16]),
    .Y(n268));
 SDFHx4_ASAP7_75t_SL i122 (.CLK(clk),
    .D(n443),
    .QN(n21[6]),
    .SE(n1229),
    .SI(n1047));
 INVx1_ASAP7_75t_SL i1220 (.A(n37[22]),
    .Y(n267));
 INVx2_ASAP7_75t_SL i1221 (.A(n32[2]),
    .Y(n131));
 INVx1_ASAP7_75t_SL i1222 (.A(n2[2]),
    .Y(n187));
 INVx1_ASAP7_75t_SL i1223 (.A(n36[5]),
    .Y(n266));
 INVx1_ASAP7_75t_SL i1224 (.A(n37[24]),
    .Y(n265));
 INVx1_ASAP7_75t_SL i1225 (.A(n35[24]),
    .Y(n264));
 INVx1_ASAP7_75t_SL i1226 (.A(n35[21]),
    .Y(n263));
 INVx1_ASAP7_75t_SL i1227 (.A(n35[28]),
    .Y(n262));
 INVx1_ASAP7_75t_SL i1228 (.A(n12[2]),
    .Y(n153));
 INVx2_ASAP7_75t_SL i1229 (.A(n16[0]),
    .Y(n173));
 SDFHx4_ASAP7_75t_SL i123 (.CLK(clk),
    .D(n401),
    .QN(n21[7]),
    .SE(n1229),
    .SI(n1132));
 INVx4_ASAP7_75t_SL i1230 (.A(n18[0]),
    .Y(n133));
 INVx1_ASAP7_75t_SL i1231 (.A(n36[23]),
    .Y(n261));
 INVx1_ASAP7_75t_SL i1232 (.A(n35[10]),
    .Y(n260));
 INVx1_ASAP7_75t_SL i1233 (.A(n35[9]),
    .Y(n259));
 INVx1_ASAP7_75t_SL i1234 (.A(n37[17]),
    .Y(n258));
 INVx1_ASAP7_75t_SL i1235 (.A(n36[11]),
    .Y(n257));
 INVx3_ASAP7_75t_SL i1236 (.A(n26[1]),
    .Y(n174));
 INVx1_ASAP7_75t_SL i1237 (.A(n35[30]),
    .Y(n256));
 INVx1_ASAP7_75t_SL i1238 (.A(n35[23]),
    .Y(n255));
 INVx1_ASAP7_75t_SL i1239 (.A(n35[22]),
    .Y(n254));
 SDFHx4_ASAP7_75t_SL i124 (.CLK(clk),
    .D(n453),
    .QN(n19[0]),
    .SE(n1229),
    .SI(n1131));
 INVx1_ASAP7_75t_SL i1240 (.A(n37[11]),
    .Y(n253));
 INVx1_ASAP7_75t_SL i1241 (.A(n36[16]),
    .Y(n252));
 INVx1_ASAP7_75t_SL i1242 (.A(n37[8]),
    .Y(n251));
 INVx1_ASAP7_75t_SL i1243 (.A(n36[17]),
    .Y(n250));
 INVx1_ASAP7_75t_SL i1244 (.A(n36[10]),
    .Y(n249));
 INVx1_ASAP7_75t_SL i1245 (.A(n35[25]),
    .Y(n248));
 INVx1_ASAP7_75t_SL i1246 (.A(n35[11]),
    .Y(n247));
 INVx1_ASAP7_75t_SL i1247 (.A(n35[8]),
    .Y(n246));
 INVx1_ASAP7_75t_SL i1248 (.A(n36[8]),
    .Y(n245));
 INVx1_ASAP7_75t_SL i1249 (.A(n36[19]),
    .Y(n244));
 SDFHx4_ASAP7_75t_SL i125 (.CLK(clk),
    .D(n439),
    .QN(n19[2]),
    .SE(n1229),
    .SI(n1130));
 INVx1_ASAP7_75t_SL i1250 (.A(n35[19]),
    .Y(n243));
 INVx1_ASAP7_75t_SL i1251 (.A(n35[3]),
    .Y(n242));
 INVx3_ASAP7_75t_SL i1252 (.A(n28[1]),
    .Y(n175));
 INVx1_ASAP7_75t_SL i1253 (.A(n36[7]),
    .Y(n241));
 INVx2_ASAP7_75t_SL i1254 (.A(n14[1]),
    .Y(n151));
 INVxp33_ASAP7_75t_SL i1255 (.A(n35[6]),
    .Y(n240));
 INVx1_ASAP7_75t_SL i1256 (.A(n36[3]),
    .Y(n239));
 INVx1_ASAP7_75t_SL i1257 (.A(n4[1]),
    .Y(n164));
 INVx1_ASAP7_75t_SL i1258 (.A(n37[7]),
    .Y(n238));
 INVx1_ASAP7_75t_SL i1259 (.A(n36[1]),
    .Y(n237));
 SDFHx4_ASAP7_75t_SL i126 (.CLK(clk),
    .D(n416),
    .QN(n19[3]),
    .SE(n1229),
    .SI(n1121));
 INVx1_ASAP7_75t_SL i1260 (.A(n35[12]),
    .Y(n236));
 INVx1_ASAP7_75t_SL i1261 (.A(n1151),
    .Y(n235));
 INVx1_ASAP7_75t_SL i1262 (.A(n37[4]),
    .Y(n234));
 INVx1_ASAP7_75t_SL i1263 (.A(n36[18]),
    .Y(n233));
 INVx1_ASAP7_75t_SL i1264 (.A(n36[14]),
    .Y(n232));
 INVx1_ASAP7_75t_SL i1265 (.A(n37[3]),
    .Y(n231));
 INVx1_ASAP7_75t_SL i1266 (.A(n6[1]),
    .Y(n166));
 INVx3_ASAP7_75t_SL i1267 (.A(n6[6]),
    .Y(n167));
 INVx3_ASAP7_75t_SL i1268 (.A(n32[5]),
    .Y(n157));
 INVx1_ASAP7_75t_SL i1269 (.A(n4[5]),
    .Y(n155));
 SDFHx4_ASAP7_75t_SL i127 (.CLK(clk),
    .D(n454),
    .QN(n19[4]),
    .SE(n1229),
    .SI(n1120));
 INVx3_ASAP7_75t_SL i1270 (.A(n24[4]),
    .Y(n158));
 INVx3_ASAP7_75t_SL i1271 (.A(n6[2]),
    .Y(n148));
 INVx2_ASAP7_75t_L i1272 (.A(n10[5]),
    .Y(n199));
 INVx3_ASAP7_75t_SL i1273 (.A(n16[2]),
    .Y(n156));
 INVx3_ASAP7_75t_SL i1274 (.A(n14[2]),
    .Y(n141));
 INVx3_ASAP7_75t_SL i1275 (.A(n26[2]),
    .Y(n163));
 INVx3_ASAP7_75t_SL i1276 (.A(n2[4]),
    .Y(n184));
 INVx3_ASAP7_75t_SL i1277 (.A(n2[0]),
    .Y(n194));
 INVx3_ASAP7_75t_SL i1278 (.A(n26[4]),
    .Y(n161));
 INVx3_ASAP7_75t_SL i1279 (.A(n22[6]),
    .Y(n152));
 SDFHx4_ASAP7_75t_SL i128 (.CLK(clk),
    .D(n455),
    .QN(n19[5]),
    .SE(n1229),
    .SI(n1043));
 INVx3_ASAP7_75t_SL i1280 (.A(n10[2]),
    .Y(n145));
 INVx3_ASAP7_75t_SL i1281 (.A(n30[1]),
    .Y(n159));
 INVx2_ASAP7_75t_SL i1282 (.A(n24[5]),
    .Y(n195));
 INVx3_ASAP7_75t_SL i1283 (.A(n24[2]),
    .Y(n160));
 INVx3_ASAP7_75t_SL i1284 (.A(n28[4]),
    .Y(n154));
 INVx2_ASAP7_75t_SL i1285 (.A(n10[0]),
    .Y(n180));
 INVx3_ASAP7_75t_SL i1286 (.A(n28[5]),
    .Y(n188));
 INVx2_ASAP7_75t_SL i1287 (.A(n24[1]),
    .Y(n230));
 INVx2_ASAP7_75t_SL i1288 (.A(n4[0]),
    .Y(n138));
 INVx2_ASAP7_75t_SL i1289 (.A(n22[2]),
    .Y(n229));
 SDFHx4_ASAP7_75t_SL i129 (.CLK(clk),
    .D(n457),
    .QN(n19[6]),
    .SE(n1229),
    .SI(n1042));
 INVx2_ASAP7_75t_SL i1290 (.A(n14[5]),
    .Y(n190));
 INVx2_ASAP7_75t_SL i1291 (.A(n20[5]),
    .Y(n143));
 INVx3_ASAP7_75t_SL i1292 (.A(n30[2]),
    .Y(n198));
 INVx3_ASAP7_75t_SL i1293 (.A(n18[6]),
    .Y(n193));
 INVx2_ASAP7_75t_SL i1294 (.A(n18[1]),
    .Y(n228));
 INVx3_ASAP7_75t_SL i1295 (.A(n28[0]),
    .Y(n146));
 INVx2_ASAP7_75t_SL i1296 (.A(n16[5]),
    .Y(n200));
 INVx3_ASAP7_75t_SL i1297 (.A(n2[5]),
    .Y(n181));
 INVx3_ASAP7_75t_SL i1298 (.A(n26[5]),
    .Y(n140));
 INVx1_ASAP7_75t_SL i1299 (.A(n8[5]),
    .Y(n139));
 INVxp67_ASAP7_75t_R i13 (.A(n20[6]),
    .Y(n96));
 SDFHx4_ASAP7_75t_SL i130 (.CLK(clk),
    .D(n458),
    .QN(n19[7]),
    .SE(n1229),
    .SI(n1129));
 INVx4_ASAP7_75t_SL i1300 (.A(n20[2]),
    .Y(n168));
 INVx3_ASAP7_75t_SL i1301 (.A(n20[1]),
    .Y(n142));
 INVx3_ASAP7_75t_SL i1302 (.A(n12[0]),
    .Y(n137));
 INVx1_ASAP7_75t_SL i1303 (.A(n30[3]),
    .Y(n165));
 INVx3_ASAP7_75t_SL i1304 (.A(n28[2]),
    .Y(n186));
 INVx2_ASAP7_75t_SL i1305 (.A(n26[0]),
    .Y(n136));
 INVx2_ASAP7_75t_SL i1306 (.A(n6[0]),
    .Y(n169));
 INVx3_ASAP7_75t_SL i1307 (.A(n16[6]),
    .Y(n185));
 INVx3_ASAP7_75t_SL i1308 (.A(n10[6]),
    .Y(n171));
 INVx3_ASAP7_75t_SL i1309 (.A(n1153),
    .Y(n227));
 SDFHx4_ASAP7_75t_SL i131 (.CLK(clk),
    .D(n461),
    .QN(n17[0]),
    .SE(n1229),
    .SI(n1041));
 INVx3_ASAP7_75t_SL i1310 (.A(n1155),
    .Y(n226));
 XNOR2xp5_ASAP7_75t_SL i1311 (.A(n486),
    .B(n930),
    .Y(n225));
 XOR2x2_ASAP7_75t_SL i1312 (.A(n34[31]),
    .B(n4[7]),
    .Y(n224));
 XNOR2x1_ASAP7_75t_SL i1313 (.B(n18[3]),
    .Y(n223),
    .A(n28[3]));
 XNOR2xp5_ASAP7_75t_SL i1314 (.A(n34[13]),
    .B(n101),
    .Y(n222));
 XNOR2xp5_ASAP7_75t_SL i1315 (.A(n37[15]),
    .B(n93),
    .Y(n221));
 XNOR2xp5_ASAP7_75t_SL i1316 (.A(n35[13]),
    .B(n98),
    .Y(n220));
 XOR2x2_ASAP7_75t_SL i1317 (.A(n35[31]),
    .B(n6[7]),
    .Y(n219));
 XNOR2xp5_ASAP7_75t_SL i1318 (.A(n36[31]),
    .B(n8[7]),
    .Y(n218));
 XNOR2x2_ASAP7_75t_SL i1319 (.A(n35[0]),
    .B(n16[0]),
    .Y(n217));
 SDFHx4_ASAP7_75t_SL i132 (.CLK(clk),
    .D(n462),
    .QN(n17[1]),
    .SE(n1229),
    .SI(n1040));
 DFFHQNx1_ASAP7_75t_SL i1320 (.CLK(clk),
    .D(n210),
    .QN(net259));
 SDFHx4_ASAP7_75t_SL i1321 (.CLK(clk),
    .D(n209),
    .QN(n25[2]),
    .SE(n1229),
    .SI(n216));
 SDFHx4_ASAP7_75t_SL i1322 (.CLK(clk),
    .D(n207),
    .QN(n21[1]),
    .SE(n1229),
    .SI(n215));
 SDFHx4_ASAP7_75t_SL i1323 (.CLK(clk),
    .D(n208),
    .QN(n19[1]),
    .SE(n1229),
    .SI(n214));
 SDFHx1_ASAP7_75t_SL i1324 (.CLK(clk),
    .QN(net260),
    .D(n138),
    .SE(n34[0]),
    .SI(n4[0]));
 SDFHx1_ASAP7_75t_SL i1325 (.CLK(clk),
    .QN(net299),
    .D(n164),
    .SE(n34[1]),
    .SI(n4[1]));
 SDFHx1_ASAP7_75t_SL i1326 (.CLK(clk),
    .QN(net310),
    .D(n183),
    .SE(n34[2]),
    .SI(n4[2]));
 SDFHx1_ASAP7_75t_SL i1327 (.CLK(clk),
    .QN(net321),
    .D(n120),
    .SE(n34[3]),
    .SI(n4[3]));
 SDFHx1_ASAP7_75t_SL i1328 (.CLK(clk),
    .QN(net332),
    .D(n119),
    .SE(n34[4]),
    .SI(n4[4]));
 SDFHx1_ASAP7_75t_SL i1329 (.CLK(clk),
    .QN(net343),
    .D(n155),
    .SE(n34[5]),
    .SI(n4[5]));
 SDFHx4_ASAP7_75t_SL i133 (.CLK(clk),
    .D(n463),
    .QN(n17[2]),
    .SE(n1229),
    .SI(n1201));
 SDFHx1_ASAP7_75t_SL i1330 (.CLK(clk),
    .QN(net354),
    .D(n118),
    .SE(n34[6]),
    .SI(n4[6]));
 SDFHx1_ASAP7_75t_SL i1331 (.CLK(clk),
    .QN(net365),
    .D(n117),
    .SE(n34[7]),
    .SI(n4[7]));
 SDFHx1_ASAP7_75t_SL i1332 (.CLK(clk),
    .QN(net376),
    .D(n132),
    .SE(n34[8]),
    .SI(n14[0]));
 SDFHx1_ASAP7_75t_SL i1333 (.CLK(clk),
    .QN(net387),
    .D(n151),
    .SE(n34[9]),
    .SI(n14[1]));
 SDFHx1_ASAP7_75t_SL i1334 (.CLK(clk),
    .QN(net271),
    .D(n141),
    .SE(n34[10]),
    .SI(n14[2]));
 SDFHx1_ASAP7_75t_SL i1335 (.CLK(clk),
    .QN(net282),
    .D(n102),
    .SE(n34[11]),
    .SI(n14[3]));
 SDFHx1_ASAP7_75t_SL i1336 (.CLK(clk),
    .QN(net291),
    .D(n101),
    .SE(n34[12]),
    .SI(n14[4]));
 SDFHx1_ASAP7_75t_SL i1337 (.CLK(clk),
    .QN(net292),
    .D(n190),
    .SE(n34[13]),
    .SI(n14[5]));
 SDFHx1_ASAP7_75t_SL i1338 (.CLK(clk),
    .QN(net293),
    .D(n100),
    .SE(n34[14]),
    .SI(n14[6]));
 SDFHx1_ASAP7_75t_SL i1339 (.CLK(clk),
    .QN(net294),
    .D(n1157),
    .SE(n34[15]),
    .SI(n14[7]));
 SDFHx4_ASAP7_75t_SL i134 (.CLK(clk),
    .D(n466),
    .QN(n17[3]),
    .SE(n1229),
    .SI(n1127));
 SDFHx1_ASAP7_75t_SL i1340 (.CLK(clk),
    .QN(net295),
    .D(n130),
    .SE(n34[16]),
    .SI(n24[0]));
 SDFHx1_ASAP7_75t_SL i1341 (.CLK(clk),
    .QN(net296),
    .D(n68),
    .SE(n24[1]),
    .SI(n34[17]));
 SDFHx1_ASAP7_75t_SL i1342 (.CLK(clk),
    .QN(net297),
    .D(n160),
    .SE(n34[18]),
    .SI(n24[2]));
 SDFHx1_ASAP7_75t_SL i1343 (.CLK(clk),
    .QN(net298),
    .D(n1222),
    .SE(n34[19]),
    .SI(n24[3]));
 SDFHx1_ASAP7_75t_SL i1344 (.CLK(clk),
    .QN(net300),
    .D(n158),
    .SE(n34[20]),
    .SI(n24[4]));
 SDFHx1_ASAP7_75t_SL i1345 (.CLK(clk),
    .QN(net301),
    .D(n195),
    .SE(n34[21]),
    .SI(n24[5]));
 SDFHx1_ASAP7_75t_SL i1346 (.CLK(clk),
    .QN(net302),
    .D(n92),
    .SE(n34[22]),
    .SI(n24[6]));
 SDFHx1_ASAP7_75t_SL i1347 (.CLK(clk),
    .QN(net303),
    .D(n1156),
    .SE(n34[23]),
    .SI(n24[7]));
 SDFHx1_ASAP7_75t_SL i1348 (.CLK(clk),
    .QN(net304),
    .D(n136),
    .SE(n34[24]),
    .SI(n26[0]));
 SDFHx1_ASAP7_75t_SL i1349 (.CLK(clk),
    .QN(net305),
    .D(n174),
    .SE(n34[25]),
    .SI(n26[1]));
 SDFHx4_ASAP7_75t_SL i135 (.CLK(clk),
    .D(n467),
    .QN(n17[4]),
    .SE(n1229),
    .SI(n1039));
 SDFHx1_ASAP7_75t_SL i1350 (.CLK(clk),
    .QN(net306),
    .D(n163),
    .SE(n34[26]),
    .SI(n26[2]));
 SDFHx1_ASAP7_75t_SL i1351 (.CLK(clk),
    .QN(net307),
    .D(n1227),
    .SE(n34[27]),
    .SI(n26[3]));
 SDFHx1_ASAP7_75t_SL i1352 (.CLK(clk),
    .QN(net308),
    .D(n161),
    .SE(n34[28]),
    .SI(n26[4]));
 SDFHx1_ASAP7_75t_SL i1353 (.CLK(clk),
    .QN(net309),
    .D(n140),
    .SE(n34[29]),
    .SI(n26[5]));
 SDFHx1_ASAP7_75t_SL i1354 (.CLK(clk),
    .QN(net311),
    .D(n91),
    .SE(n34[30]),
    .SI(n26[6]));
 SDFHx1_ASAP7_75t_SL i1355 (.CLK(clk),
    .QN(net312),
    .D(n90),
    .SE(n34[31]),
    .SI(n26[7]));
 SDFHx1_ASAP7_75t_SL i1356 (.CLK(clk),
    .QN(net313),
    .D(n169),
    .SE(n35[0]),
    .SI(n6[0]));
 SDFHx1_ASAP7_75t_SL i1357 (.CLK(clk),
    .QN(net314),
    .D(n166),
    .SE(n35[1]),
    .SI(n6[1]));
 SDFHx1_ASAP7_75t_SL i1358 (.CLK(clk),
    .QN(net315),
    .D(n148),
    .SE(n35[2]),
    .SI(n6[2]));
 SDFHx1_ASAP7_75t_SL i1359 (.CLK(clk),
    .QN(net316),
    .D(n116),
    .SE(n35[3]),
    .SI(n6[3]));
 SDFHx4_ASAP7_75t_SL i136 (.CLK(clk),
    .D(n470),
    .QN(n17[5]),
    .SE(n1229),
    .SI(n1126));
 SDFHx1_ASAP7_75t_SL i1360 (.CLK(clk),
    .QN(net317),
    .D(n115),
    .SE(n35[4]),
    .SI(n6[4]));
 SDFHx1_ASAP7_75t_SL i1361 (.CLK(clk),
    .QN(net318),
    .D(n170),
    .SE(n35[5]),
    .SI(n6[5]));
 SDFHx1_ASAP7_75t_SL i1362 (.CLK(clk),
    .QN(net319),
    .D(n167),
    .SE(n35[6]),
    .SI(n6[6]));
 SDFHx1_ASAP7_75t_SL i1363 (.CLK(clk),
    .QN(net320),
    .D(n114),
    .SE(n35[7]),
    .SI(n6[7]));
 SDFHx1_ASAP7_75t_SL i1364 (.CLK(clk),
    .QN(net322),
    .D(n173),
    .SE(n35[8]),
    .SI(n16[0]));
 SDFHx1_ASAP7_75t_SL i1365 (.CLK(clk),
    .QN(net323),
    .D(n191),
    .SE(n35[9]),
    .SI(n16[1]));
 SDFHx1_ASAP7_75t_SL i1366 (.CLK(clk),
    .QN(net324),
    .D(n156),
    .SE(n35[10]),
    .SI(n16[2]));
 SDFHx1_ASAP7_75t_SL i1367 (.CLK(clk),
    .QN(net325),
    .D(n99),
    .SE(n35[11]),
    .SI(n16[3]));
 SDFHx1_ASAP7_75t_SL i1368 (.CLK(clk),
    .QN(net326),
    .D(n98),
    .SE(n35[12]),
    .SI(n16[4]));
 SDFHx1_ASAP7_75t_SL i1369 (.CLK(clk),
    .QN(net327),
    .D(n200),
    .SE(n35[13]),
    .SI(n16[5]));
 SDFHx4_ASAP7_75t_SL i137 (.CLK(clk),
    .D(n472),
    .QN(n17[6]),
    .SE(n1229),
    .SI(n1037));
 SDFHx1_ASAP7_75t_SL i1370 (.CLK(clk),
    .QN(net328),
    .D(n185),
    .SE(n35[14]),
    .SI(n16[6]));
 SDFHx1_ASAP7_75t_SL i1371 (.CLK(clk),
    .QN(net329),
    .D(n1161),
    .SE(n35[15]),
    .SI(n16[7]));
 SDFHx1_ASAP7_75t_SL i1372 (.CLK(clk),
    .QN(net330),
    .D(n133),
    .SE(n35[16]),
    .SI(n18[0]));
 SDFHx1_ASAP7_75t_SL i1373 (.CLK(clk),
    .QN(net331),
    .D(n129),
    .SE(n18[1]),
    .SI(n35[17]));
 SDFHx1_ASAP7_75t_SL i1374 (.CLK(clk),
    .QN(net333),
    .D(n189),
    .SE(n35[18]),
    .SI(n18[2]));
 SDFHx1_ASAP7_75t_SL i1375 (.CLK(clk),
    .QN(net334),
    .D(n179),
    .SE(n35[19]),
    .SI(n18[3]));
 SDFHx1_ASAP7_75t_SL i1376 (.CLK(clk),
    .QN(net335),
    .D(n178),
    .SE(n35[20]),
    .SI(n18[4]));
 SDFHx1_ASAP7_75t_SL i1377 (.CLK(clk),
    .QN(net336),
    .D(n144),
    .SE(n35[21]),
    .SI(n18[5]));
 SDFHx1_ASAP7_75t_SL i1378 (.CLK(clk),
    .QN(net337),
    .D(n193),
    .SE(n35[22]),
    .SI(n18[6]));
 SDFHx1_ASAP7_75t_SL i1379 (.CLK(clk),
    .QN(net338),
    .D(n1160),
    .SE(n35[23]),
    .SI(n18[7]));
 SDFHx4_ASAP7_75t_SL i138 (.CLK(clk),
    .D(n364),
    .QN(n17[7]),
    .SE(n1229),
    .SI(n1114));
 SDFHx1_ASAP7_75t_SL i1380 (.CLK(clk),
    .QN(net339),
    .D(n146),
    .SE(n35[24]),
    .SI(n28[0]));
 SDFHx1_ASAP7_75t_SL i1381 (.CLK(clk),
    .QN(net340),
    .D(n175),
    .SE(n35[25]),
    .SI(n28[1]));
 SDFHx1_ASAP7_75t_SL i1382 (.CLK(clk),
    .QN(net341),
    .D(n186),
    .SE(n35[26]),
    .SI(n28[2]));
 SDFHx1_ASAP7_75t_SL i1383 (.CLK(clk),
    .QN(net342),
    .D(n182),
    .SE(n35[27]),
    .SI(n28[3]));
 SDFHx1_ASAP7_75t_SL i1384 (.CLK(clk),
    .QN(net344),
    .D(n154),
    .SE(n35[28]),
    .SI(n28[4]));
 SDFHx1_ASAP7_75t_SL i1385 (.CLK(clk),
    .QN(net345),
    .D(n188),
    .SE(n35[29]),
    .SI(n28[5]));
 SDFHx1_ASAP7_75t_SL i1386 (.CLK(clk),
    .QN(net346),
    .D(n1220),
    .SE(n35[30]),
    .SI(n28[6]));
 SDFHx1_ASAP7_75t_SL i1387 (.CLK(clk),
    .QN(net347),
    .D(n89),
    .SE(n35[31]),
    .SI(n28[7]));
 SDFHx1_ASAP7_75t_SL i1388 (.CLK(clk),
    .QN(net348),
    .D(n149),
    .SE(n36[0]),
    .SI(n8[0]));
 SDFHx1_ASAP7_75t_SL i1389 (.CLK(clk),
    .QN(net349),
    .D(n150),
    .SE(n36[1]),
    .SI(n8[1]));
 SDFHx4_ASAP7_75t_SL i139 (.CLK(clk),
    .D(n362),
    .QN(n15[0]),
    .SE(n1229),
    .SI(n1112));
 SDFHx1_ASAP7_75t_SL i1390 (.CLK(clk),
    .QN(net350),
    .D(n113),
    .SE(n36[2]),
    .SI(n8[2]));
 SDFHx1_ASAP7_75t_SL i1391 (.CLK(clk),
    .QN(net351),
    .D(n112),
    .SE(n36[3]),
    .SI(n8[3]));
 SDFHx1_ASAP7_75t_SL i1392 (.CLK(clk),
    .QN(net352),
    .D(n111),
    .SE(n36[4]),
    .SI(n8[4]));
 SDFHx1_ASAP7_75t_SL i1393 (.CLK(clk),
    .QN(net353),
    .D(n139),
    .SE(n36[5]),
    .SI(n8[5]));
 SDFHx1_ASAP7_75t_SL i1394 (.CLK(clk),
    .QN(net355),
    .D(n134),
    .SE(n36[6]),
    .SI(n8[6]));
 SDFHx1_ASAP7_75t_SL i1395 (.CLK(clk),
    .QN(net356),
    .D(n110),
    .SE(n36[7]),
    .SI(n8[7]));
 SDFHx1_ASAP7_75t_SL i1396 (.CLK(clk),
    .QN(net357),
    .D(n180),
    .SE(n36[8]),
    .SI(n10[0]));
 SDFHx1_ASAP7_75t_SL i1397 (.CLK(clk),
    .QN(net358),
    .D(n109),
    .SE(n36[9]),
    .SI(n10[1]));
 SDFHx1_ASAP7_75t_SL i1398 (.CLK(clk),
    .QN(net359),
    .D(n145),
    .SE(n36[10]),
    .SI(n10[2]));
 SDFHx1_ASAP7_75t_SL i1399 (.CLK(clk),
    .QN(net360),
    .D(n1158),
    .SE(n36[11]),
    .SI(n10[3]));
 INVx2_ASAP7_75t_SL i14 (.A(n20[0]),
    .Y(n97));
 SDFHx4_ASAP7_75t_SL i140 (.CLK(clk),
    .D(n361),
    .QN(n15[1]),
    .SE(n1229),
    .SI(n1111));
 SDFHx1_ASAP7_75t_SL i1400 (.CLK(clk),
    .QN(net361),
    .D(n196),
    .SE(n36[12]),
    .SI(n10[4]));
 SDFHx1_ASAP7_75t_SL i1401 (.CLK(clk),
    .QN(net362),
    .D(n199),
    .SE(n36[13]),
    .SI(n10[5]));
 SDFHx1_ASAP7_75t_SL i1402 (.CLK(clk),
    .QN(net363),
    .D(n171),
    .SE(n36[14]),
    .SI(n10[6]));
 SDFHx1_ASAP7_75t_SL i1403 (.CLK(clk),
    .QN(net364),
    .D(n108),
    .SE(n36[15]),
    .SI(n10[7]));
 SDFHx1_ASAP7_75t_SL i1404 (.CLK(clk),
    .QN(net366),
    .D(n97),
    .SE(n36[16]),
    .SI(n20[0]));
 SDFHx1_ASAP7_75t_SL i1405 (.CLK(clk),
    .QN(net367),
    .D(n142),
    .SE(n36[17]),
    .SI(n20[1]));
 SDFHx1_ASAP7_75t_SL i1406 (.CLK(clk),
    .QN(net368),
    .D(n168),
    .SE(n36[18]),
    .SI(n20[2]));
 SDFHx1_ASAP7_75t_SL i1407 (.CLK(clk),
    .QN(net369),
    .D(n1159),
    .SE(n36[19]),
    .SI(n20[3]));
 SDFHx1_ASAP7_75t_SL i1408 (.CLK(clk),
    .QN(net370),
    .D(n162),
    .SE(n36[20]),
    .SI(n20[4]));
 SDFHx1_ASAP7_75t_SL i1409 (.CLK(clk),
    .QN(net371),
    .D(n143),
    .SE(n36[21]),
    .SI(n20[5]));
 SDFHx4_ASAP7_75t_SL i141 (.CLK(clk),
    .D(n359),
    .QN(n15[2]),
    .SE(n1229),
    .SI(n1216));
 SDFHx1_ASAP7_75t_SL i1410 (.CLK(clk),
    .QN(net372),
    .D(n96),
    .SE(n36[22]),
    .SI(n20[6]));
 SDFHx1_ASAP7_75t_SL i1411 (.CLK(clk),
    .QN(net373),
    .D(n95),
    .SE(n36[23]),
    .SI(n20[7]));
 SDFHx1_ASAP7_75t_SL i1412 (.CLK(clk),
    .QN(net374),
    .D(n88),
    .SE(n36[24]),
    .SI(n30[0]));
 SDFHx1_ASAP7_75t_SL i1413 (.CLK(clk),
    .QN(net375),
    .D(n159),
    .SE(n36[25]),
    .SI(n30[1]));
 SDFHx1_ASAP7_75t_SL i1414 (.CLK(clk),
    .QN(net377),
    .D(n198),
    .SE(n36[26]),
    .SI(n30[2]));
 SDFHx1_ASAP7_75t_SL i1415 (.CLK(clk),
    .QN(net378),
    .D(n165),
    .SE(n36[27]),
    .SI(n30[3]));
 SDFHx1_ASAP7_75t_SL i1416 (.CLK(clk),
    .QN(net379),
    .D(n87),
    .SE(n36[28]),
    .SI(n30[4]));
 SDFHx1_ASAP7_75t_SL i1417 (.CLK(clk),
    .QN(net380),
    .D(n1164),
    .SE(n36[29]),
    .SI(n30[5]));
 SDFHx1_ASAP7_75t_SL i1418 (.CLK(clk),
    .QN(net381),
    .D(n135),
    .SE(n36[30]),
    .SI(n30[6]));
 SDFHx1_ASAP7_75t_SL i1419 (.CLK(clk),
    .QN(net382),
    .D(n86),
    .SE(n36[31]),
    .SI(n30[7]));
 SDFHx4_ASAP7_75t_SL i142 (.CLK(clk),
    .D(n358),
    .QN(n15[3]),
    .SE(n1229),
    .SI(n1109));
 SDFHx1_ASAP7_75t_SL i1420 (.CLK(clk),
    .QN(net383),
    .D(n194),
    .SE(n37[0]),
    .SI(n2[0]));
 SDFHx1_ASAP7_75t_SL i1421 (.CLK(clk),
    .QN(net384),
    .D(n192),
    .SE(n37[1]),
    .SI(n2[1]));
 SDFHx1_ASAP7_75t_SL i1422 (.CLK(clk),
    .QN(net385),
    .D(n187),
    .SE(n37[2]),
    .SI(n2[2]));
 SDFHx1_ASAP7_75t_SL i1423 (.CLK(clk),
    .QN(net386),
    .D(n123),
    .SE(n37[3]),
    .SI(n2[3]));
 SDFHx1_ASAP7_75t_SL i1424 (.CLK(clk),
    .QN(net261),
    .D(n184),
    .SE(n37[4]),
    .SI(n2[4]));
 SDFHx1_ASAP7_75t_SL i1425 (.CLK(clk),
    .QN(net262),
    .D(n181),
    .SE(n37[5]),
    .SI(n2[5]));
 SDFHx1_ASAP7_75t_SL i1426 (.CLK(clk),
    .QN(net263),
    .D(n122),
    .SE(n37[6]),
    .SI(n2[6]));
 SDFHx1_ASAP7_75t_SL i1427 (.CLK(clk),
    .QN(net264),
    .D(n121),
    .SE(n37[7]),
    .SI(n2[7]));
 SDFHx1_ASAP7_75t_SL i1428 (.CLK(clk),
    .QN(net265),
    .D(n137),
    .SE(n37[8]),
    .SI(n12[0]));
 SDFHx1_ASAP7_75t_SL i1429 (.CLK(clk),
    .QN(net266),
    .D(n177),
    .SE(n37[9]),
    .SI(n12[1]));
 SDFHx4_ASAP7_75t_SL i143 (.CLK(clk),
    .D(n357),
    .QN(n15[4]),
    .SE(n1229),
    .SI(n1108));
 SDFHx1_ASAP7_75t_SL i1430 (.CLK(clk),
    .QN(net267),
    .D(n153),
    .SE(n37[10]),
    .SI(n12[2]));
 SDFHx1_ASAP7_75t_SL i1431 (.CLK(clk),
    .QN(net268),
    .D(n107),
    .SE(n37[11]),
    .SI(n12[3]));
 SDFHx1_ASAP7_75t_SL i1432 (.CLK(clk),
    .QN(net269),
    .D(n106),
    .SE(n37[12]),
    .SI(n12[4]));
 SDFHx1_ASAP7_75t_SL i1433 (.CLK(clk),
    .QN(net270),
    .D(n105),
    .SE(n37[13]),
    .SI(n12[5]));
 SDFHx1_ASAP7_75t_SL i1434 (.CLK(clk),
    .QN(net272),
    .D(n104),
    .SE(n37[14]),
    .SI(n12[6]));
 SDFHx1_ASAP7_75t_SL i1435 (.CLK(clk),
    .QN(net273),
    .D(n103),
    .SE(n37[15]),
    .SI(n12[7]));
 SDFHx1_ASAP7_75t_SL i1436 (.CLK(clk),
    .QN(net274),
    .D(n1225),
    .SE(n37[16]),
    .SI(n22[0]));
 SDFHx1_ASAP7_75t_SL i1437 (.CLK(clk),
    .QN(net275),
    .D(n176),
    .SE(n37[17]),
    .SI(n22[1]));
 SDFHx1_ASAP7_75t_SL i1438 (.CLK(clk),
    .QN(net276),
    .D(n47),
    .SE(n22[2]),
    .SI(n37[18]));
 SDFHx1_ASAP7_75t_SL i1439 (.CLK(clk),
    .QN(net277),
    .D(n1166),
    .SE(n37[19]),
    .SI(n22[3]));
 SDFHx4_ASAP7_75t_SL i144 (.CLK(clk),
    .D(n355),
    .QN(n15[5]),
    .SE(n1229),
    .SI(n1148));
 SDFHx1_ASAP7_75t_SL i1440 (.CLK(clk),
    .QN(net278),
    .D(n1221),
    .SE(n37[20]),
    .SI(n22[4]));
 SDFHx1_ASAP7_75t_SL i1441 (.CLK(clk),
    .QN(net279),
    .D(n94),
    .SE(n37[21]),
    .SI(n22[5]));
 SDFHx1_ASAP7_75t_SL i1442 (.CLK(clk),
    .QN(net280),
    .D(n152),
    .SE(n37[22]),
    .SI(n22[6]));
 SDFHx1_ASAP7_75t_SL i1443 (.CLK(clk),
    .QN(net281),
    .D(n93),
    .SE(n37[23]),
    .SI(n22[7]));
 SDFHx1_ASAP7_75t_SL i1444 (.CLK(clk),
    .QN(net283),
    .D(n1165),
    .SE(n37[24]),
    .SI(n32[0]));
 SDFHx1_ASAP7_75t_SL i1445 (.CLK(clk),
    .QN(net284),
    .D(n147),
    .SE(n37[25]),
    .SI(n32[1]));
 SDFHx1_ASAP7_75t_SL i1446 (.CLK(clk),
    .QN(net285),
    .D(n131),
    .SE(n37[26]),
    .SI(n32[2]));
 SDFHx1_ASAP7_75t_SL i1447 (.CLK(clk),
    .QN(net286),
    .D(n1162),
    .SE(n37[27]),
    .SI(n32[3]));
 SDFHx1_ASAP7_75t_SL i1448 (.CLK(clk),
    .QN(net287),
    .D(n197),
    .SE(n37[28]),
    .SI(n32[4]));
 SDFHx1_ASAP7_75t_SL i1449 (.CLK(clk),
    .QN(net288),
    .D(n157),
    .SE(n37[29]),
    .SI(n32[5]));
 SDFHx4_ASAP7_75t_SL i145 (.CLK(clk),
    .D(n353),
    .QN(n15[6]),
    .SE(n1229),
    .SI(n1106));
 SDFHx1_ASAP7_75t_SL i1450 (.CLK(clk),
    .QN(net289),
    .D(n85),
    .SE(n37[30]),
    .SI(n32[6]));
 SDFHx1_ASAP7_75t_SL i1451 (.CLK(clk),
    .QN(net290),
    .D(n84),
    .SE(n37[31]),
    .SI(n32[7]));
 XNOR2xp5_ASAP7_75t_SL i1452 (.A(n205),
    .B(n213),
    .Y(n216));
 XOR2xp5_ASAP7_75t_SL i1453 (.A(n127),
    .B(n212),
    .Y(n215));
 XOR2xp5_ASAP7_75t_SL i1454 (.A(n128),
    .B(n211),
    .Y(n214));
 XOR2xp5_ASAP7_75t_SL i1455 (.A(n1151),
    .B(n203),
    .Y(n213));
 XOR2xp5_ASAP7_75t_SL i1456 (.A(n202),
    .B(n206),
    .Y(n212));
 XOR2xp5_ASAP7_75t_SL i1457 (.A(n201),
    .B(n204),
    .Y(n211));
 OR3x1_ASAP7_75t_SL i1458 (.A(n1150),
    .B(n172),
    .C(net129),
    .Y(n210));
 XNOR2xp5_ASAP7_75t_SL i1459 (.A(n0[114]),
    .B(n37[18]),
    .Y(n209));
 SDFHx4_ASAP7_75t_SL i146 (.CLK(clk),
    .D(n350),
    .QN(n15[7]),
    .SE(n1229),
    .SI(n1105));
 XNOR2xp5_ASAP7_75t_SL i1460 (.A(n34[17]),
    .B(n0[17]),
    .Y(n208));
 XNOR2xp5_ASAP7_75t_SL i1461 (.A(n0[49]),
    .B(n35[17]),
    .Y(n207));
 AOI22xp5_ASAP7_75t_SL i1462 (.A1(n35[17]),
    .A2(n175),
    .B1(n129),
    .B2(n28[1]),
    .Y(n206));
 AOI22xp5_ASAP7_75t_SL i1463 (.A1(n37[18]),
    .A2(n176),
    .B1(n47),
    .B2(n22[1]),
    .Y(n205));
 AOI22xp5_ASAP7_75t_SL i1464 (.A1(n34[17]),
    .A2(n174),
    .B1(n68),
    .B2(n26[1]),
    .Y(n204));
 AOI22xp5_ASAP7_75t_R i1465 (.A1(n32[2]),
    .A2(n177),
    .B1(n12[1]),
    .B2(n131),
    .Y(n203));
 OAI22xp5_ASAP7_75t_SL i1466 (.A1(n16[0]),
    .A2(n133),
    .B1(n18[0]),
    .B2(n173),
    .Y(n202));
 OAI22xp5_ASAP7_75t_SL i1467 (.A1(n14[0]),
    .A2(n130),
    .B1(n24[0]),
    .B2(n132),
    .Y(n201));
 INVxp67_ASAP7_75t_R i1468 (.A(n18[3]),
    .Y(n179));
 INVx4_ASAP7_75t_SL i1469 (.A(n12[1]),
    .Y(n177));
 SDFHx4_ASAP7_75t_SL i147 (.CLK(clk),
    .D(n349),
    .QN(n13[0]),
    .SE(n1229),
    .SI(n1118));
 INVxp67_ASAP7_75t_SL i1470 (.A(n35[17]),
    .Y(n129));
 XOR2xp5_ASAP7_75t_SL i1471 (.A(n1154),
    .B(n1155),
    .Y(n128));
 XOR2xp5_ASAP7_75t_SL i1472 (.A(n1152),
    .B(n1153),
    .Y(n127));
 INVx2_ASAP7_75t_SL i1473 (.A(n24[7]),
    .Y(n1156));
 INVx2_ASAP7_75t_SL i1474 (.A(n14[7]),
    .Y(n1157));
 INVx3_ASAP7_75t_SL i1475 (.A(n10[3]),
    .Y(n1158));
 INVxp67_ASAP7_75t_SL i1476 (.A(n20[3]),
    .Y(n1159));
 INVx2_ASAP7_75t_SL i1477 (.A(n18[7]),
    .Y(n1160));
 INVx2_ASAP7_75t_SL i1478 (.A(n16[7]),
    .Y(n1161));
 INVx1_ASAP7_75t_SL i1479 (.A(n32[3]),
    .Y(n1162));
 SDFHx4_ASAP7_75t_SL i148 (.CLK(clk),
    .D(n365),
    .QN(n13[1]),
    .SE(n1229),
    .SI(n1104));
 INVx4_ASAP7_75t_SL i1480 (.A(n476),
    .Y(n1163));
 INVx2_ASAP7_75t_SL i1481 (.A(n30[5]),
    .Y(n1164));
 INVx1_ASAP7_75t_SL i1482 (.A(n32[0]),
    .Y(n1165));
 INVx1_ASAP7_75t_SL i1483 (.A(n22[3]),
    .Y(n1166));
 OAI22xp5_ASAP7_75t_SL i1484 (.A1(n119),
    .A2(n26[4]),
    .B1(n4[4]),
    .B2(n161),
    .Y(n1167));
 OAI22xp5_ASAP7_75t_SL i1485 (.A1(n119),
    .A2(n26[4]),
    .B1(n4[4]),
    .B2(n161),
    .Y(n1168));
 XOR2xp5_ASAP7_75t_SL i1486 (.A(n857),
    .B(n495),
    .Y(n1169));
 XOR2xp5_ASAP7_75t_SL i1487 (.A(n841),
    .B(n773),
    .Y(n1170));
 XOR2xp5_ASAP7_75t_SL i1488 (.A(n823),
    .B(n816),
    .Y(n1171));
 XOR2xp5_ASAP7_75t_SL i1489 (.A(n578),
    .B(n484),
    .Y(n1172));
 SDFHx4_ASAP7_75t_SL i149 (.CLK(clk),
    .D(n366),
    .QN(n13[2]),
    .SE(n1229),
    .SI(n1147));
 XOR2xp5_ASAP7_75t_SL i1490 (.A(n37[19]),
    .B(n32[3]),
    .Y(n1173));
 XNOR2xp5_ASAP7_75t_SL i1491 (.A(n22[3]),
    .B(n37[27]),
    .Y(n1174));
 XOR2x2_ASAP7_75t_SL i1492 (.A(n22[0]),
    .B(n32[0]),
    .Y(n1175));
 XNOR2x1_ASAP7_75t_SL i1493 (.B(n22[3]),
    .Y(n1176),
    .A(n32[3]));
 XNOR2x1_ASAP7_75t_SL i1494 (.B(n20[3]),
    .Y(n1177),
    .A(n30[3]));
 XNOR2xp5_ASAP7_75t_SL i1495 (.A(n36[4]),
    .B(n30[4]),
    .Y(n1178));
 XNOR2xp5_ASAP7_75t_SL i1496 (.A(n30[4]),
    .B(n36[29]),
    .Y(n1179));
 XNOR2xp5_ASAP7_75t_SL i1497 (.A(n20[3]),
    .B(n36[27]),
    .Y(n1180));
 XOR2xp5_ASAP7_75t_SL i1498 (.A(n36[21]),
    .B(n30[5]),
    .Y(n1181));
 OAI22xp5_ASAP7_75t_SL i1499 (.A1(n570),
    .A2(n1183),
    .B1(n1182),
    .B2(n569),
    .Y(n1184));
 INVx1_ASAP7_75t_SL i15 (.A(n16[4]),
    .Y(n98));
 SDFHx4_ASAP7_75t_SL i150 (.CLK(clk),
    .D(n368),
    .QN(n13[3]),
    .SE(n1229),
    .SI(n1102));
 INVx3_ASAP7_75t_SL i1500 (.A(n1182),
    .Y(n1183));
 OA22x2_ASAP7_75t_SL i1501 (.A1(n114),
    .A2(n28[7]),
    .B1(n89),
    .B2(n6[7]),
    .Y(n1182));
 AOI22xp5_ASAP7_75t_SL i1502 (.A1(n1183),
    .A2(n863),
    .B1(n862),
    .B2(n1182),
    .Y(n1185));
 XNOR2xp5_ASAP7_75t_SL i1503 (.A(n1182),
    .B(n919),
    .Y(n1186));
 AOI22xp5_ASAP7_75t_SL i1504 (.A1(n486),
    .A2(n1183),
    .B1(n487),
    .B2(n1182),
    .Y(n1187));
 AOI22xp5_ASAP7_75t_SL i1505 (.A1(n1183),
    .A2(n223),
    .B1(n1182),
    .B2(n778),
    .Y(n1188));
 AOI22xp5_ASAP7_75t_SL i1506 (.A1(n796),
    .A2(n1183),
    .B1(n797),
    .B2(n1182),
    .Y(n1189));
 OAI22xp5_ASAP7_75t_SL i1507 (.A1(n554),
    .A2(n1191),
    .B1(n1190),
    .B2(n553),
    .Y(n1192));
 INVx3_ASAP7_75t_SL i1508 (.A(n1190),
    .Y(n1191));
 OA22x2_ASAP7_75t_SL i1509 (.A1(n117),
    .A2(n26[7]),
    .B1(n90),
    .B2(n4[7]),
    .Y(n1190));
 SDFHx4_ASAP7_75t_SL i151 (.CLK(clk),
    .D(n371),
    .QN(n13[4]),
    .SE(n1229),
    .SI(n1101));
 AOI22xp5_ASAP7_75t_SL i1510 (.A1(n558),
    .A2(n1191),
    .B1(n557),
    .B2(n1190),
    .Y(n1193));
 XNOR2xp5_ASAP7_75t_SL i1511 (.A(n1190),
    .B(n918),
    .Y(n1194));
 AOI22xp5_ASAP7_75t_SL i1512 (.A1(n790),
    .A2(n1191),
    .B1(n791),
    .B2(n1190),
    .Y(n1195));
 AOI22xp5_ASAP7_75t_SL i1513 (.A1(n1191),
    .A2(n1232),
    .B1(n1190),
    .B2(n777),
    .Y(n1196));
 AOI22xp5_ASAP7_75t_SL i1514 (.A1(n812),
    .A2(n1191),
    .B1(n813),
    .B2(n1190),
    .Y(n1197));
 INVx3_ASAP7_75t_SL i1515 (.A(n2[1]),
    .Y(n192));
 OAI22xp5_ASAP7_75t_SL i1516 (.A1(n1198),
    .A2(n761),
    .B1(n1199),
    .B2(n760),
    .Y(n1200));
 AO22x2_ASAP7_75t_SL i1517 (.A1(n2[1]),
    .A2(n177),
    .B1(n192),
    .B2(n12[1]),
    .Y(n1198));
 INVx2_ASAP7_75t_SL i1518 (.A(n1198),
    .Y(n1199));
 XNOR2xp5_ASAP7_75t_SL i1519 (.A(n1198),
    .B(n916),
    .Y(n1201));
 SDFHx4_ASAP7_75t_SL i152 (.CLK(clk),
    .D(n372),
    .QN(n13[5]),
    .SE(n1229),
    .SI(n1145));
 OAI22xp5_ASAP7_75t_SL i1520 (.A1(n1198),
    .A2(n474),
    .B1(n124),
    .B2(n1199),
    .Y(n1202));
 AOI22xp5_ASAP7_75t_SL i1521 (.A1(n1204),
    .A2(n1177),
    .B1(n769),
    .B2(n1203),
    .Y(n1205));
 INVx3_ASAP7_75t_SL i1522 (.A(n1203),
    .Y(n1204));
 OA22x2_ASAP7_75t_SL i1523 (.A1(n110),
    .A2(n30[7]),
    .B1(n86),
    .B2(n8[7]),
    .Y(n1203));
 XNOR2xp5_ASAP7_75t_SL i1524 (.A(n1203),
    .B(n985),
    .Y(n1206));
 AOI22xp5_ASAP7_75t_SL i1525 (.A1(n787),
    .A2(n1204),
    .B1(n788),
    .B2(n1203),
    .Y(n1207));
 AOI22xp5_ASAP7_75t_SL i1526 (.A1(n1210),
    .A2(n1204),
    .B1(n502),
    .B2(n1203),
    .Y(n1208));
 AOI22xp5_ASAP7_75t_SL i1527 (.A1(n1204),
    .A2(n540),
    .B1(n539),
    .B2(n1203),
    .Y(n1209));
 XNOR2x1_ASAP7_75t_SL i1528 (.B(n20[4]),
    .Y(n1210),
    .A(n10[4]));
 INVx2_ASAP7_75t_SL i1529 (.A(n10[4]),
    .Y(n196));
 SDFHx4_ASAP7_75t_SL i153 (.CLK(clk),
    .D(n374),
    .QN(n13[6]),
    .SE(n1229),
    .SI(n1100));
 INVx1_ASAP7_75t_SL i1530 (.A(n20[4]),
    .Y(n162));
 XNOR2x1_ASAP7_75t_SL i1531 (.B(n20[7]),
    .Y(n1211),
    .A(n30[7]));
 XOR2xp5_ASAP7_75t_SL i1532 (.A(n35[20]),
    .B(n18[3]),
    .Y(n1212));
 INVx2_ASAP7_75t_SL i1533 (.A(n26[3]),
    .Y(n1227));
 INVx3_ASAP7_75t_SL i1534 (.A(n8[1]),
    .Y(n150));
 OAI22xp5_ASAP7_75t_SL i1535 (.A1(n1213),
    .A2(n1211),
    .B1(n1214),
    .B2(n479),
    .Y(n1215));
 AO22x2_ASAP7_75t_SL i1536 (.A1(n8[1]),
    .A2(n109),
    .B1(n150),
    .B2(n10[1]),
    .Y(n1213));
 INVx1_ASAP7_75t_SL i1537 (.A(n1213),
    .Y(n1214));
 XNOR2xp5_ASAP7_75t_SL i1538 (.A(n1213),
    .B(n1023),
    .Y(n1216));
 OAI22xp5_ASAP7_75t_SL i1539 (.A1(n1213),
    .A2(n476),
    .B1(n1163),
    .B2(n1214),
    .Y(n1217));
 SDFHx4_ASAP7_75t_SL i154 (.CLK(clk),
    .D(n375),
    .QN(n13[7]),
    .SE(n1229),
    .SI(n1099));
 OAI22xp5_ASAP7_75t_SL i1540 (.A1(n1218),
    .A2(n1204),
    .B1(n1203),
    .B2(n1226),
    .Y(n1219));
 INVx1_ASAP7_75t_SL i1541 (.A(n1226),
    .Y(n1218));
 INVx2_ASAP7_75t_SL i1542 (.A(n28[6]),
    .Y(n1220));
 INVx1_ASAP7_75t_SL i1543 (.A(n22[4]),
    .Y(n1221));
 INVx2_ASAP7_75t_SL i1544 (.A(n24[3]),
    .Y(n1222));
 OAI22xp5_ASAP7_75t_SL i1545 (.A1(n48),
    .A2(n12[4]),
    .B1(n37[13]),
    .B2(n106),
    .Y(n1223));
 OAI22xp5_ASAP7_75t_SL i1546 (.A1(n12[3]),
    .A2(n106),
    .B1(n12[4]),
    .B2(n107),
    .Y(n1224));
 INVx1_ASAP7_75t_SL i1547 (.A(n22[0]),
    .Y(n1225));
 XNOR2xp5_ASAP7_75t_SL i1548 (.A(n36[15]),
    .B(n95),
    .Y(n1226));
 INVx4_ASAP7_75t_SL i1549 (.A(n1228),
    .Y(n1229));
 SDFHx4_ASAP7_75t_SL i155 (.CLK(clk),
    .D(n376),
    .QN(n11[0]),
    .SE(n1229),
    .SI(n1116));
 DFFHQNx1_ASAP7_75t_SL i1550 (.CLK(clk),
    .D(n38),
    .QN(n1228));
 XOR2xp5_ASAP7_75t_SL i1551 (.A(n37[12]),
    .B(n22[4]),
    .Y(n1230));
 XNOR2xp5_ASAP7_75t_SL i1552 (.A(n18[3]),
    .B(n35[27]),
    .Y(n1231));
 XNOR2x1_ASAP7_75t_SL i1553 (.B(n24[3]),
    .Y(n1232),
    .A(n26[3]));
 HAxp5_ASAP7_75t_R i1554 (.A(n0[95]),
    .B(n36[31]),
    .CON(n126),
    .SN(n389));
 SDFHx4_ASAP7_75t_SL i156 (.CLK(clk),
    .D(n379),
    .QN(n11[1]),
    .SE(n1229),
    .SI(n1097));
 SDFHx4_ASAP7_75t_SL i157 (.CLK(clk),
    .D(n381),
    .QN(n11[2]),
    .SE(n1229),
    .SI(n1144));
 SDFHx4_ASAP7_75t_SL i158 (.CLK(clk),
    .D(n382),
    .QN(n11[3]),
    .SE(n1229),
    .SI(n1095));
 SDFHx4_ASAP7_75t_SL i159 (.CLK(clk),
    .D(n384),
    .QN(n11[4]),
    .SE(n1229),
    .SI(n1093));
 INVx1_ASAP7_75t_SL i16 (.A(n16[3]),
    .Y(n99));
 SDFHx4_ASAP7_75t_SL i160 (.CLK(clk),
    .D(n385),
    .QN(n11[5]),
    .SE(n1229),
    .SI(n1142));
 SDFHx4_ASAP7_75t_SL i161 (.CLK(clk),
    .D(n388),
    .QN(n11[6]),
    .SE(n1229),
    .SI(n1149));
 SDFHx4_ASAP7_75t_SL i162 (.CLK(clk),
    .D(n390),
    .QN(n11[7]),
    .SE(n1229),
    .SI(n1031));
 SDFHx4_ASAP7_75t_SL i163 (.CLK(clk),
    .D(n391),
    .QN(n9[0]),
    .SE(n1229),
    .SI(n1036));
 SDFHx4_ASAP7_75t_SL i164 (.CLK(clk),
    .D(n393),
    .QN(n9[1]),
    .SE(n1229),
    .SI(n1089));
 SDFHx4_ASAP7_75t_SL i165 (.CLK(clk),
    .D(n394),
    .QN(n9[2]),
    .SE(n1229),
    .SI(n1141));
 SDFHx4_ASAP7_75t_SL i166 (.CLK(clk),
    .D(n397),
    .QN(n9[3]),
    .SE(n1229),
    .SI(n1087));
 SDFHx4_ASAP7_75t_SL i167 (.CLK(clk),
    .D(n398),
    .QN(n9[4]),
    .SE(n1229),
    .SI(n1086));
 SDFHx4_ASAP7_75t_SL i168 (.CLK(clk),
    .D(n402),
    .QN(n9[5]),
    .SE(n1229),
    .SI(n1085));
 SDFHx4_ASAP7_75t_SL i169 (.CLK(clk),
    .D(n403),
    .QN(n9[6]),
    .SE(n1229),
    .SI(n1084));
 INVxp33_ASAP7_75t_SL i17 (.A(n14[6]),
    .Y(n100));
 SDFHx4_ASAP7_75t_SL i170 (.CLK(clk),
    .D(n405),
    .QN(n9[7]),
    .SE(n1229),
    .SI(n1034));
 SDFHx4_ASAP7_75t_SL i171 (.CLK(clk),
    .D(n407),
    .QN(n7[0]),
    .SE(n1229),
    .SI(n1206));
 SDFHx4_ASAP7_75t_SL i172 (.CLK(clk),
    .D(n409),
    .QN(n7[1]),
    .SE(n1229),
    .SI(n1080));
 SDFHx4_ASAP7_75t_SL i173 (.CLK(clk),
    .D(n410),
    .QN(n7[2]),
    .SE(n1229),
    .SI(n1140));
 SDFHx4_ASAP7_75t_SL i174 (.CLK(clk),
    .D(n412),
    .QN(n7[3]),
    .SE(n1229),
    .SI(n1078));
 SDFHx4_ASAP7_75t_SL i175 (.CLK(clk),
    .D(n414),
    .QN(n7[4]),
    .SE(n1229),
    .SI(n1077));
 SDFHx4_ASAP7_75t_SL i176 (.CLK(clk),
    .D(n418),
    .QN(n7[5]),
    .SE(n1229),
    .SI(n1075));
 SDFHx4_ASAP7_75t_SL i177 (.CLK(clk),
    .D(n419),
    .QN(n7[6]),
    .SE(n1229),
    .SI(n1073));
 SDFHx4_ASAP7_75t_SL i178 (.CLK(clk),
    .D(n420),
    .QN(n7[7]),
    .SE(n1229),
    .SI(n1033));
 SDFHx4_ASAP7_75t_SL i179 (.CLK(clk),
    .D(n421),
    .QN(n5[0]),
    .SE(n1229),
    .SI(n1186));
 INVxp67_ASAP7_75t_SL i18 (.A(n14[4]),
    .Y(n101));
 SDFHx4_ASAP7_75t_SL i180 (.CLK(clk),
    .D(n434),
    .QN(n5[1]),
    .SE(n1229),
    .SI(n1071));
 SDFHx4_ASAP7_75t_SL i181 (.CLK(clk),
    .D(n452),
    .QN(n5[2]),
    .SE(n1229),
    .SI(n1070));
 SDFHx4_ASAP7_75t_SL i182 (.CLK(clk),
    .D(n425),
    .QN(n5[3]),
    .SE(n1229),
    .SI(n1069));
 SDFHx4_ASAP7_75t_SL i183 (.CLK(clk),
    .D(n427),
    .QN(n5[4]),
    .SE(n1229),
    .SI(n1067));
 SDFHx4_ASAP7_75t_SL i184 (.CLK(clk),
    .D(n428),
    .QN(n5[5]),
    .SE(n1229),
    .SI(n1064));
 SDFHx4_ASAP7_75t_SL i185 (.CLK(clk),
    .D(n429),
    .QN(n5[6]),
    .SE(n1229),
    .SI(n1063));
 SDFHx4_ASAP7_75t_SL i186 (.CLK(clk),
    .D(n432),
    .QN(n5[7]),
    .SE(n1229),
    .SI(n1137));
 SDFHx4_ASAP7_75t_SL i187 (.CLK(clk),
    .D(n435),
    .QN(n3[0]),
    .SE(n1229),
    .SI(n1194));
 SDFHx4_ASAP7_75t_SL i188 (.CLK(clk),
    .D(n433),
    .QN(n3[1]),
    .SE(n1229),
    .SI(n1062));
 SDFHx4_ASAP7_75t_SL i189 (.CLK(clk),
    .D(n437),
    .QN(n3[2]),
    .SE(n1229),
    .SI(n1060));
 INVx2_ASAP7_75t_SL i19 (.A(n14[3]),
    .Y(n102));
 SDFHx4_ASAP7_75t_SL i190 (.CLK(clk),
    .D(n413),
    .QN(n3[3]),
    .SE(n1229),
    .SI(n1057));
 SDFHx4_ASAP7_75t_SL i191 (.CLK(clk),
    .D(n400),
    .QN(n3[4]),
    .SE(n1229),
    .SI(n1056));
 SDFHx4_ASAP7_75t_SL i192 (.CLK(clk),
    .D(n440),
    .QN(n3[5]),
    .SE(n1229),
    .SI(n1055));
 SDFHx4_ASAP7_75t_SL i193 (.CLK(clk),
    .D(n441),
    .QN(n3[6]),
    .SE(n1229),
    .SI(n1053));
 SDFHx4_ASAP7_75t_SL i194 (.CLK(clk),
    .D(n442),
    .QN(n3[7]),
    .SE(n1229),
    .SI(n1136));
 DFFHQNx1_ASAP7_75t_SL i195 (.CLK(clk),
    .D(n727),
    .QN(n0[0]));
 DFFHQNx1_ASAP7_75t_SL i196 (.CLK(clk),
    .D(n753),
    .QN(n0[1]));
 DFFHQNx1_ASAP7_75t_SL i197 (.CLK(clk),
    .D(n726),
    .QN(n0[2]));
 DFFHQNx1_ASAP7_75t_SL i198 (.CLK(clk),
    .D(n725),
    .QN(n0[3]));
 DFFHQNx1_ASAP7_75t_SL i199 (.CLK(clk),
    .D(n724),
    .QN(n0[4]));
 INVxp33_ASAP7_75t_SL i2 (.A(n32[6]),
    .Y(n85));
 INVx2_ASAP7_75t_SL i20 (.A(n12[7]),
    .Y(n103));
 DFFHQNx1_ASAP7_75t_SL i200 (.CLK(clk),
    .D(n723),
    .QN(n0[5]));
 DFFHQNx1_ASAP7_75t_SL i201 (.CLK(clk),
    .D(n722),
    .QN(n0[6]));
 DFFHQNx1_ASAP7_75t_SL i202 (.CLK(clk),
    .D(n721),
    .QN(n0[7]));
 DFFHQNx1_ASAP7_75t_SL i203 (.CLK(clk),
    .D(n720),
    .QN(n0[8]));
 DFFHQNx1_ASAP7_75t_SL i204 (.CLK(clk),
    .D(n719),
    .QN(n0[9]));
 DFFHQNx1_ASAP7_75t_SL i205 (.CLK(clk),
    .D(n718),
    .QN(n0[10]));
 DFFHQNx1_ASAP7_75t_SL i206 (.CLK(clk),
    .D(n737),
    .QN(n0[11]));
 DFFHQNx1_ASAP7_75t_SL i207 (.CLK(clk),
    .D(n717),
    .QN(n0[12]));
 DFFHQNx1_ASAP7_75t_SL i208 (.CLK(clk),
    .D(n716),
    .QN(n0[13]));
 DFFHQNx1_ASAP7_75t_SL i209 (.CLK(clk),
    .D(n715),
    .QN(n0[14]));
 INVxp33_ASAP7_75t_SL i21 (.A(n12[6]),
    .Y(n104));
 DFFHQNx1_ASAP7_75t_SL i210 (.CLK(clk),
    .D(n714),
    .QN(n0[15]));
 DFFHQNx1_ASAP7_75t_SL i211 (.CLK(clk),
    .D(n713),
    .QN(n0[16]));
 DFFHQNx1_ASAP7_75t_SL i212 (.CLK(clk),
    .D(n712),
    .QN(n0[17]));
 DFFHQNx1_ASAP7_75t_SL i213 (.CLK(clk),
    .D(n711),
    .QN(n0[18]));
 DFFHQNx1_ASAP7_75t_SL i214 (.CLK(clk),
    .D(n743),
    .QN(n0[19]));
 DFFHQNx1_ASAP7_75t_SL i215 (.CLK(clk),
    .D(n710),
    .QN(n0[20]));
 DFFHQNx1_ASAP7_75t_SL i216 (.CLK(clk),
    .D(n709),
    .QN(n0[21]));
 DFFHQNx1_ASAP7_75t_SL i217 (.CLK(clk),
    .D(n708),
    .QN(n0[22]));
 DFFHQNx1_ASAP7_75t_SL i218 (.CLK(clk),
    .D(n749),
    .QN(n0[23]));
 DFFHQNx1_ASAP7_75t_SL i219 (.CLK(clk),
    .D(n707),
    .QN(n0[24]));
 INVxp67_ASAP7_75t_R i22 (.A(n12[5]),
    .Y(n105));
 DFFHQNx1_ASAP7_75t_SL i220 (.CLK(clk),
    .D(n706),
    .QN(n0[25]));
 DFFHQNx1_ASAP7_75t_SL i221 (.CLK(clk),
    .D(n705),
    .QN(n0[26]));
 DFFHQNx1_ASAP7_75t_SL i222 (.CLK(clk),
    .D(n704),
    .QN(n0[27]));
 DFFHQNx1_ASAP7_75t_SL i223 (.CLK(clk),
    .D(n703),
    .QN(n0[28]));
 DFFHQNx1_ASAP7_75t_SL i224 (.CLK(clk),
    .D(n702),
    .QN(n0[29]));
 DFFHQNx1_ASAP7_75t_SL i225 (.CLK(clk),
    .D(n701),
    .QN(n0[30]));
 DFFHQNx1_ASAP7_75t_SL i226 (.CLK(clk),
    .D(n700),
    .QN(n0[31]));
 DFFHQNx1_ASAP7_75t_SL i227 (.CLK(clk),
    .D(n699),
    .QN(n0[32]));
 DFFHQNx1_ASAP7_75t_SL i228 (.CLK(clk),
    .D(n698),
    .QN(n0[33]));
 DFFHQNx1_ASAP7_75t_SL i229 (.CLK(clk),
    .D(n697),
    .QN(n0[34]));
 INVx1_ASAP7_75t_SL i23 (.A(n12[4]),
    .Y(n106));
 DFFHQNx1_ASAP7_75t_SL i230 (.CLK(clk),
    .D(n696),
    .QN(n0[35]));
 DFFHQNx1_ASAP7_75t_SL i231 (.CLK(clk),
    .D(n695),
    .QN(n0[36]));
 DFFHQNx1_ASAP7_75t_SL i232 (.CLK(clk),
    .D(n694),
    .QN(n0[37]));
 DFFHQNx1_ASAP7_75t_SL i233 (.CLK(clk),
    .D(n693),
    .QN(n0[38]));
 DFFHQNx1_ASAP7_75t_SL i234 (.CLK(clk),
    .D(n692),
    .QN(n0[39]));
 DFFHQNx1_ASAP7_75t_SL i235 (.CLK(clk),
    .D(n691),
    .QN(n0[40]));
 DFFHQNx1_ASAP7_75t_SL i236 (.CLK(clk),
    .D(n690),
    .QN(n0[41]));
 DFFHQNx1_ASAP7_75t_SL i237 (.CLK(clk),
    .D(n689),
    .QN(n0[42]));
 DFFHQNx1_ASAP7_75t_SL i238 (.CLK(clk),
    .D(n746),
    .QN(n0[43]));
 DFFHQNx1_ASAP7_75t_SL i239 (.CLK(clk),
    .D(n688),
    .QN(n0[44]));
 INVx2_ASAP7_75t_SL i24 (.A(n12[3]),
    .Y(n107));
 DFFHQNx1_ASAP7_75t_SL i240 (.CLK(clk),
    .D(n687),
    .QN(n0[45]));
 DFFHQNx1_ASAP7_75t_SL i241 (.CLK(clk),
    .D(n686),
    .QN(n0[46]));
 DFFHQNx1_ASAP7_75t_SL i242 (.CLK(clk),
    .D(n685),
    .QN(n0[47]));
 DFFHQNx1_ASAP7_75t_SL i243 (.CLK(clk),
    .D(n684),
    .QN(n0[48]));
 DFFHQNx1_ASAP7_75t_SL i244 (.CLK(clk),
    .D(n748),
    .QN(n0[49]));
 DFFHQNx1_ASAP7_75t_SL i245 (.CLK(clk),
    .D(n683),
    .QN(n0[50]));
 DFFHQNx1_ASAP7_75t_SL i246 (.CLK(clk),
    .D(n732),
    .QN(n0[51]));
 DFFHQNx1_ASAP7_75t_SL i247 (.CLK(clk),
    .D(n735),
    .QN(n0[52]));
 DFFHQNx1_ASAP7_75t_SL i248 (.CLK(clk),
    .D(n742),
    .QN(n0[53]));
 DFFHQNx1_ASAP7_75t_SL i249 (.CLK(clk),
    .D(n682),
    .QN(n0[54]));
 INVx1_ASAP7_75t_SL i25 (.A(n10[7]),
    .Y(n108));
 DFFHQNx1_ASAP7_75t_SL i250 (.CLK(clk),
    .D(n681),
    .QN(n0[55]));
 DFFHQNx1_ASAP7_75t_SL i251 (.CLK(clk),
    .D(n680),
    .QN(n0[56]));
 DFFHQNx1_ASAP7_75t_SL i252 (.CLK(clk),
    .D(n679),
    .QN(n0[57]));
 DFFHQNx1_ASAP7_75t_SL i253 (.CLK(clk),
    .D(n678),
    .QN(n0[58]));
 DFFHQNx1_ASAP7_75t_SL i254 (.CLK(clk),
    .D(n677),
    .QN(n0[59]));
 DFFHQNx1_ASAP7_75t_SL i255 (.CLK(clk),
    .D(n676),
    .QN(n0[60]));
 DFFHQNx1_ASAP7_75t_SL i256 (.CLK(clk),
    .D(n675),
    .QN(n0[61]));
 DFFHQNx1_ASAP7_75t_SL i257 (.CLK(clk),
    .D(n674),
    .QN(n0[62]));
 DFFHQNx1_ASAP7_75t_SL i258 (.CLK(clk),
    .D(n673),
    .QN(n0[63]));
 DFFHQNx1_ASAP7_75t_SL i259 (.CLK(clk),
    .D(n672),
    .QN(n0[64]));
 INVx2_ASAP7_75t_SL i26 (.A(n10[1]),
    .Y(n109));
 DFFHQNx1_ASAP7_75t_SL i260 (.CLK(clk),
    .D(n671),
    .QN(n0[65]));
 DFFHQNx1_ASAP7_75t_SL i261 (.CLK(clk),
    .D(n670),
    .QN(n0[66]));
 DFFHQNx1_ASAP7_75t_SL i262 (.CLK(clk),
    .D(n669),
    .QN(n0[67]));
 DFFHQNx1_ASAP7_75t_SL i263 (.CLK(clk),
    .D(n755),
    .QN(n0[68]));
 DFFHQNx1_ASAP7_75t_SL i264 (.CLK(clk),
    .D(n668),
    .QN(n0[69]));
 DFFHQNx1_ASAP7_75t_SL i265 (.CLK(clk),
    .D(n667),
    .QN(n0[70]));
 DFFHQNx1_ASAP7_75t_SL i266 (.CLK(clk),
    .D(n666),
    .QN(n0[71]));
 DFFHQNx1_ASAP7_75t_SL i267 (.CLK(clk),
    .D(n665),
    .QN(n0[72]));
 DFFHQNx1_ASAP7_75t_SL i268 (.CLK(clk),
    .D(n664),
    .QN(n0[73]));
 DFFHQNx1_ASAP7_75t_SL i269 (.CLK(clk),
    .D(n730),
    .QN(n0[74]));
 INVxp67_ASAP7_75t_SL i27 (.A(n8[7]),
    .Y(n110));
 DFFHQNx1_ASAP7_75t_SL i270 (.CLK(clk),
    .D(n731),
    .QN(n0[75]));
 DFFHQNx1_ASAP7_75t_SL i271 (.CLK(clk),
    .D(n663),
    .QN(n0[76]));
 DFFHQNx1_ASAP7_75t_SL i272 (.CLK(clk),
    .D(n662),
    .QN(n0[77]));
 DFFHQNx1_ASAP7_75t_SL i273 (.CLK(clk),
    .D(n661),
    .QN(n0[78]));
 DFFHQNx1_ASAP7_75t_SL i274 (.CLK(clk),
    .D(n738),
    .QN(n0[79]));
 DFFHQNx1_ASAP7_75t_SL i275 (.CLK(clk),
    .D(n740),
    .QN(n0[80]));
 DFFHQNx1_ASAP7_75t_SL i276 (.CLK(clk),
    .D(n660),
    .QN(n0[81]));
 DFFHQNx1_ASAP7_75t_SL i277 (.CLK(clk),
    .D(n659),
    .QN(n0[82]));
 DFFHQNx1_ASAP7_75t_SL i278 (.CLK(clk),
    .D(n658),
    .QN(n0[83]));
 DFFHQNx1_ASAP7_75t_SL i279 (.CLK(clk),
    .D(n657),
    .QN(n0[84]));
 INVxp67_ASAP7_75t_R i28 (.A(n8[4]),
    .Y(n111));
 DFFHQNx1_ASAP7_75t_SL i280 (.CLK(clk),
    .D(n656),
    .QN(n0[85]));
 DFFHQNx1_ASAP7_75t_SL i281 (.CLK(clk),
    .D(n750),
    .QN(n0[86]));
 DFFHQNx1_ASAP7_75t_SL i282 (.CLK(clk),
    .D(n655),
    .QN(n0[87]));
 DFFHQNx1_ASAP7_75t_SL i283 (.CLK(clk),
    .D(n654),
    .QN(n0[88]));
 DFFHQNx1_ASAP7_75t_SL i284 (.CLK(clk),
    .D(n653),
    .QN(n0[89]));
 DFFHQNx1_ASAP7_75t_SL i285 (.CLK(clk),
    .D(n628),
    .QN(n0[90]));
 DFFHQNx1_ASAP7_75t_SL i286 (.CLK(clk),
    .D(n652),
    .QN(n0[91]));
 DFFHQNx1_ASAP7_75t_SL i287 (.CLK(clk),
    .D(n651),
    .QN(n0[92]));
 DFFHQNx1_ASAP7_75t_SL i288 (.CLK(clk),
    .D(n650),
    .QN(n0[93]));
 DFFHQNx1_ASAP7_75t_SL i289 (.CLK(clk),
    .D(n649),
    .QN(n0[94]));
 INVx2_ASAP7_75t_SL i29 (.A(n8[3]),
    .Y(n112));
 DFFHQNx1_ASAP7_75t_SL i290 (.CLK(clk),
    .D(n733),
    .QN(n0[95]));
 DFFHQNx1_ASAP7_75t_SL i291 (.CLK(clk),
    .D(n744),
    .QN(n0[96]));
 DFFHQNx1_ASAP7_75t_SL i292 (.CLK(clk),
    .D(n648),
    .QN(n0[97]));
 DFFHQNx1_ASAP7_75t_SL i293 (.CLK(clk),
    .D(n754),
    .QN(n0[98]));
 DFFHQNx1_ASAP7_75t_SL i294 (.CLK(clk),
    .D(n630),
    .QN(n0[99]));
 DFFHQNx1_ASAP7_75t_SL i295 (.CLK(clk),
    .D(n629),
    .QN(n0[100]));
 DFFHQNx1_ASAP7_75t_SL i296 (.CLK(clk),
    .D(n647),
    .QN(n0[101]));
 DFFHQNx1_ASAP7_75t_SL i297 (.CLK(clk),
    .D(n646),
    .QN(n0[102]));
 DFFHQNx1_ASAP7_75t_SL i298 (.CLK(clk),
    .D(n728),
    .QN(n0[103]));
 DFFHQNx1_ASAP7_75t_SL i299 (.CLK(clk),
    .D(n645),
    .QN(n0[104]));
 INVx2_ASAP7_75t_SL i3 (.A(n30[7]),
    .Y(n86));
 INVxp67_ASAP7_75t_R i30 (.A(n8[2]),
    .Y(n113));
 DFFHQNx1_ASAP7_75t_SL i300 (.CLK(clk),
    .D(n644),
    .QN(n0[105]));
 DFFHQNx1_ASAP7_75t_SL i301 (.CLK(clk),
    .D(n643),
    .QN(n0[106]));
 DFFHQNx1_ASAP7_75t_SL i302 (.CLK(clk),
    .D(n642),
    .QN(n0[107]));
 DFFHQNx1_ASAP7_75t_SL i303 (.CLK(clk),
    .D(n641),
    .QN(n0[108]));
 DFFHQNx1_ASAP7_75t_SL i304 (.CLK(clk),
    .D(n747),
    .QN(n0[109]));
 DFFHQNx1_ASAP7_75t_SL i305 (.CLK(clk),
    .D(n736),
    .QN(n0[110]));
 DFFHQNx1_ASAP7_75t_SL i306 (.CLK(clk),
    .D(n640),
    .QN(n0[111]));
 DFFHQNx1_ASAP7_75t_SL i307 (.CLK(clk),
    .D(n639),
    .QN(n0[112]));
 DFFHQNx1_ASAP7_75t_SL i308 (.CLK(clk),
    .D(n739),
    .QN(n0[113]));
 DFFHQNx1_ASAP7_75t_SL i309 (.CLK(clk),
    .D(n741),
    .QN(n0[114]));
 INVxp67_ASAP7_75t_SL i31 (.A(n6[7]),
    .Y(n114));
 DFFHQNx1_ASAP7_75t_SL i310 (.CLK(clk),
    .D(n745),
    .QN(n0[115]));
 DFFHQNx1_ASAP7_75t_SL i311 (.CLK(clk),
    .D(n638),
    .QN(n0[116]));
 DFFHQNx1_ASAP7_75t_SL i312 (.CLK(clk),
    .D(n637),
    .QN(n0[117]));
 DFFHQNx1_ASAP7_75t_SL i313 (.CLK(clk),
    .D(n636),
    .QN(n0[118]));
 DFFHQNx1_ASAP7_75t_SL i314 (.CLK(clk),
    .D(n635),
    .QN(n0[119]));
 DFFHQNx1_ASAP7_75t_SL i315 (.CLK(clk),
    .D(n751),
    .QN(n0[120]));
 DFFHQNx1_ASAP7_75t_SL i316 (.CLK(clk),
    .D(n752),
    .QN(n0[121]));
 DFFHQNx1_ASAP7_75t_SL i317 (.CLK(clk),
    .D(n634),
    .QN(n0[122]));
 DFFHQNx1_ASAP7_75t_SL i318 (.CLK(clk),
    .D(n633),
    .QN(n0[123]));
 DFFHQNx1_ASAP7_75t_SL i319 (.CLK(clk),
    .D(n632),
    .QN(n0[124]));
 INVx2_ASAP7_75t_SL i32 (.A(n6[4]),
    .Y(n115));
 DFFHQNx1_ASAP7_75t_SL i320 (.CLK(clk),
    .D(n729),
    .QN(n0[125]));
 DFFHQNx1_ASAP7_75t_SL i321 (.CLK(clk),
    .D(n734),
    .QN(n0[126]));
 DFFHQNx1_ASAP7_75t_SL i322 (.CLK(clk),
    .D(n631),
    .QN(n0[127]));
 XOR2xp5_ASAP7_75t_SL i323 (.A(n818),
    .B(n1000),
    .Y(n1149));
 XNOR2xp5_ASAP7_75t_SL i324 (.A(n616),
    .B(n1169),
    .Y(n1148));
 XNOR2xp5_ASAP7_75t_SL i325 (.A(n1014),
    .B(n1152),
    .Y(n1147));
 XNOR2xp5_ASAP7_75t_SL i326 (.A(n1012),
    .B(n1011),
    .Y(n1146));
 XNOR2xp5_ASAP7_75t_SL i327 (.A(n220),
    .B(n1170),
    .Y(n1145));
 XNOR2xp5_ASAP7_75t_SL i328 (.A(n1154),
    .B(n1005),
    .Y(n1144));
 XNOR2xp5_ASAP7_75t_SL i329 (.A(n808),
    .B(n1004),
    .Y(n1143));
 INVx2_ASAP7_75t_SL i33 (.A(n6[3]),
    .Y(n116));
 XNOR2xp5_ASAP7_75t_SL i330 (.A(n222),
    .B(n1171),
    .Y(n1142));
 XNOR2xp5_ASAP7_75t_SL i331 (.A(n592),
    .B(n995),
    .Y(n1141));
 XOR2xp5_ASAP7_75t_SL i332 (.A(n623),
    .B(n899),
    .Y(n1140));
 XOR2xp5_ASAP7_75t_SL i333 (.A(n326),
    .B(n881),
    .Y(n1139));
 XOR2xp5_ASAP7_75t_SL i334 (.A(n317),
    .B(n896),
    .Y(n1138));
 XOR2xp5_ASAP7_75t_SL i335 (.A(n303),
    .B(n897),
    .Y(n1137));
 XOR2xp5_ASAP7_75t_SL i336 (.A(n612),
    .B(n894),
    .Y(n1136));
 XOR2xp5_ASAP7_75t_SL i337 (.A(n319),
    .B(n1209),
    .Y(n1135));
 XOR2xp5_ASAP7_75t_SL i338 (.A(n489),
    .B(n952),
    .Y(n1134));
 XOR2xp5_ASAP7_75t_SL i339 (.A(n320),
    .B(n950),
    .Y(n1133));
 INVxp67_ASAP7_75t_SL i34 (.A(n4[7]),
    .Y(n117));
 XOR2xp5_ASAP7_75t_SL i340 (.A(n594),
    .B(n1185),
    .Y(n1132));
 XOR2xp5_ASAP7_75t_SL i341 (.A(n784),
    .B(n942),
    .Y(n1131));
 XOR2xp5_ASAP7_75t_SL i342 (.A(n611),
    .B(n940),
    .Y(n1130));
 XOR2xp5_ASAP7_75t_SL i343 (.A(n340),
    .B(n1193),
    .Y(n1129));
 XNOR2xp5_ASAP7_75t_SL i344 (.A(n931),
    .B(n932),
    .Y(n1128));
 XNOR2xp5_ASAP7_75t_SL i345 (.A(n929),
    .B(n928),
    .Y(n1127));
 XNOR2xp5_ASAP7_75t_SL i346 (.A(n1223),
    .B(n1172),
    .Y(n1126));
 XOR2xp5_ASAP7_75t_SL i347 (.A(n1017),
    .B(n776),
    .Y(n1125));
 XOR2xp5_ASAP7_75t_SL i348 (.A(n804),
    .B(n994),
    .Y(n1124));
 XOR2xp5_ASAP7_75t_SL i349 (.A(n949),
    .B(n892),
    .Y(n1123));
 INVxp33_ASAP7_75t_SL i35 (.A(n4[6]),
    .Y(n118));
 XOR2xp5_ASAP7_75t_SL i350 (.A(n947),
    .B(n891),
    .Y(n1122));
 XOR2xp5_ASAP7_75t_SL i351 (.A(n939),
    .B(n889),
    .Y(n1121));
 XOR2xp5_ASAP7_75t_SL i352 (.A(n937),
    .B(n888),
    .Y(n1120));
 XOR2xp5_ASAP7_75t_SL i353 (.A(n791),
    .B(n1008),
    .Y(n1119));
 XNOR2xp5_ASAP7_75t_SL i354 (.A(n765),
    .B(n1016),
    .Y(n1118));
 XOR2xp5_ASAP7_75t_SL i355 (.A(n921),
    .B(n758),
    .Y(n1117));
 XNOR2xp5_ASAP7_75t_SL i356 (.A(n757),
    .B(n1007),
    .Y(n1116));
 XOR2xp5_ASAP7_75t_SL i357 (.A(n917),
    .B(n477),
    .Y(n1115));
 XNOR2xp5_ASAP7_75t_SL i358 (.A(n512),
    .B(n1026),
    .Y(n1114));
 XNOR2xp5_ASAP7_75t_SL i359 (.A(n944),
    .B(n914),
    .Y(n1113));
 INVx2_ASAP7_75t_SL i36 (.A(n4[4]),
    .Y(n119));
 XNOR2xp5_ASAP7_75t_SL i360 (.A(n763),
    .B(n1025),
    .Y(n1112));
 XOR2xp5_ASAP7_75t_SL i361 (.A(n906),
    .B(n1024),
    .Y(n1111));
 XNOR2xp5_ASAP7_75t_SL i362 (.A(n766),
    .B(n1022),
    .Y(n1110));
 XOR2xp5_ASAP7_75t_SL i363 (.A(n905),
    .B(n1021),
    .Y(n1109));
 XOR2xp5_ASAP7_75t_SL i364 (.A(n904),
    .B(n1020),
    .Y(n1108));
 XOR2xp5_ASAP7_75t_SL i365 (.A(n1019),
    .B(n774),
    .Y(n1107));
 XOR2xp5_ASAP7_75t_SL i366 (.A(n501),
    .B(n1018),
    .Y(n1106));
 XNOR2xp5_ASAP7_75t_SL i367 (.A(n494),
    .B(n1219),
    .Y(n1105));
 XOR2xp5_ASAP7_75t_SL i368 (.A(n924),
    .B(n922),
    .Y(n1104));
 XNOR2xp5_ASAP7_75t_SL i369 (.A(n760),
    .B(n1015),
    .Y(n1103));
 INVx2_ASAP7_75t_SL i37 (.A(n4[3]),
    .Y(n120));
 XOR2xp5_ASAP7_75t_SL i370 (.A(n913),
    .B(n1013),
    .Y(n1102));
 XOR2xp5_ASAP7_75t_SL i371 (.A(n912),
    .B(n1010),
    .Y(n1101));
 XOR2xp5_ASAP7_75t_SL i372 (.A(n766),
    .B(n1009),
    .Y(n1100));
 XNOR2xp5_ASAP7_75t_SL i373 (.A(n775),
    .B(n1184),
    .Y(n1099));
 XNOR2xp5_ASAP7_75t_SL i374 (.A(n1006),
    .B(n911),
    .Y(n1098));
 XOR2xp5_ASAP7_75t_SL i375 (.A(n923),
    .B(n920),
    .Y(n1097));
 XNOR2xp5_ASAP7_75t_SL i376 (.A(n903),
    .B(n1200),
    .Y(n1096));
 XOR2xp5_ASAP7_75t_SL i377 (.A(n910),
    .B(n1003),
    .Y(n1095));
 XNOR2xp5_ASAP7_75t_SL i378 (.A(n1002),
    .B(n909),
    .Y(n1094));
 XOR2xp5_ASAP7_75t_SL i379 (.A(n908),
    .B(n1001),
    .Y(n1093));
 INVxp67_ASAP7_75t_SL i38 (.A(n2[7]),
    .Y(n121));
 XNOR2xp5_ASAP7_75t_SL i380 (.A(n997),
    .B(n902),
    .Y(n1092));
 XNOR2xp5_ASAP7_75t_SL i381 (.A(n818),
    .B(n999),
    .Y(n1091));
 XOR2xp5_ASAP7_75t_SL i382 (.A(n996),
    .B(n817),
    .Y(n1090));
 XOR2xp5_ASAP7_75t_SL i383 (.A(n901),
    .B(n915),
    .Y(n1089));
 XNOR2xp5_ASAP7_75t_SL i384 (.A(n992),
    .B(n900),
    .Y(n1088));
 XOR2xp5_ASAP7_75t_SL i385 (.A(n993),
    .B(n885),
    .Y(n1087));
 XOR2xp5_ASAP7_75t_SL i386 (.A(n991),
    .B(n884),
    .Y(n1086));
 XNOR2xp5_ASAP7_75t_SL i387 (.A(n485),
    .B(n990),
    .Y(n1085));
 XNOR2xp5_ASAP7_75t_SL i388 (.A(n503),
    .B(n988),
    .Y(n1084));
 XNOR2xp5_ASAP7_75t_SL i389 (.A(n987),
    .B(n1202),
    .Y(n1083));
 INVxp33_ASAP7_75t_SL i39 (.A(n2[6]),
    .Y(n122));
 XNOR2xp5_ASAP7_75t_SL i390 (.A(n983),
    .B(n883),
    .Y(n1082));
 XNOR2xp5_ASAP7_75t_SL i391 (.A(n772),
    .B(n984),
    .Y(n1081));
 XOR2xp5_ASAP7_75t_SL i392 (.A(n982),
    .B(n1207),
    .Y(n1080));
 XNOR2xp5_ASAP7_75t_SL i393 (.A(n980),
    .B(n882),
    .Y(n1079));
 XOR2xp5_ASAP7_75t_SL i394 (.A(n981),
    .B(n1205),
    .Y(n1078));
 XOR2xp5_ASAP7_75t_SL i395 (.A(n979),
    .B(n1208),
    .Y(n1077));
 XOR2xp5_ASAP7_75t_SL i396 (.A(n485),
    .B(n976),
    .Y(n1076));
 XNOR2xp5_ASAP7_75t_SL i397 (.A(n496),
    .B(n978),
    .Y(n1075));
 XNOR2xp5_ASAP7_75t_SL i398 (.A(n771),
    .B(n977),
    .Y(n1074));
 XNOR2xp5_ASAP7_75t_SL i399 (.A(n770),
    .B(n975),
    .Y(n1073));
 INVxp67_ASAP7_75t_R i4 (.A(n30[4]),
    .Y(n87));
 INVx2_ASAP7_75t_SL i40 (.A(n2[3]),
    .Y(n123));
 XNOR2xp5_ASAP7_75t_SL i400 (.A(n512),
    .B(n973),
    .Y(n1072));
 XOR2xp5_ASAP7_75t_SL i401 (.A(n1187),
    .B(n898),
    .Y(n1071));
 XOR2xp5_ASAP7_75t_SL i402 (.A(n312),
    .B(n972),
    .Y(n1070));
 XOR2xp5_ASAP7_75t_SL i403 (.A(n970),
    .B(n1188),
    .Y(n1069));
 XNOR2xp5_ASAP7_75t_SL i404 (.A(n503),
    .B(n971),
    .Y(n1068));
 XOR2xp5_ASAP7_75t_SL i405 (.A(n968),
    .B(n1189),
    .Y(n1067));
 XNOR2xp5_ASAP7_75t_SL i406 (.A(n479),
    .B(n964),
    .Y(n1066));
 XNOR2xp5_ASAP7_75t_SL i407 (.A(n967),
    .B(n1217),
    .Y(n1065));
 XNOR2xp5_ASAP7_75t_SL i408 (.A(n774),
    .B(n966),
    .Y(n1064));
 XNOR2xp5_ASAP7_75t_SL i409 (.A(n776),
    .B(n965),
    .Y(n1063));
 INVxp67_ASAP7_75t_SL i41 (.A(n474),
    .Y(n124));
 XOR2xp5_ASAP7_75t_SL i410 (.A(n895),
    .B(n1195),
    .Y(n1062));
 XNOR2xp5_ASAP7_75t_SL i411 (.A(n963),
    .B(n880),
    .Y(n1061));
 XOR2xp5_ASAP7_75t_SL i412 (.A(n302),
    .B(n962),
    .Y(n1060));
 XNOR2xp5_ASAP7_75t_SL i413 (.A(n955),
    .B(n1215),
    .Y(n1059));
 XNOR2xp5_ASAP7_75t_SL i414 (.A(n960),
    .B(n879),
    .Y(n1058));
 XOR2xp5_ASAP7_75t_SL i415 (.A(n961),
    .B(n1196),
    .Y(n1057));
 XOR2xp5_ASAP7_75t_SL i416 (.A(n959),
    .B(n1197),
    .Y(n1056));
 XNOR2xp5_ASAP7_75t_SL i417 (.A(n817),
    .B(n958),
    .Y(n1055));
 XOR2xp5_ASAP7_75t_SL i418 (.A(n788),
    .B(n953),
    .Y(n1054));
 XNOR2xp5_ASAP7_75t_SL i419 (.A(n804),
    .B(n956),
    .Y(n1053));
 INVx2_ASAP7_75t_SL i42 (.A(n475),
    .Y(n125));
 XOR2xp5_ASAP7_75t_SL i420 (.A(n957),
    .B(n501),
    .Y(n1052));
 XNOR2xp5_ASAP7_75t_SL i421 (.A(n494),
    .B(n954),
    .Y(n1051));
 XNOR2xp5_ASAP7_75t_SL i422 (.A(n951),
    .B(n893),
    .Y(n1050));
 XNOR2xp5_ASAP7_75t_SL i423 (.A(n948),
    .B(n890),
    .Y(n1049));
 XOR2xp5_ASAP7_75t_SL i424 (.A(n946),
    .B(n766),
    .Y(n1048));
 XNOR2xp5_ASAP7_75t_SL i425 (.A(n775),
    .B(n945),
    .Y(n1047));
 XNOR2xp5_ASAP7_75t_SL i426 (.A(n501),
    .B(n943),
    .Y(n1046));
 XOR2xp5_ASAP7_75t_SL i427 (.A(n496),
    .B(n941),
    .Y(n1045));
 XNOR2xp5_ASAP7_75t_SL i428 (.A(n770),
    .B(n938),
    .Y(n1044));
 XOR2xp5_ASAP7_75t_SL i429 (.A(n936),
    .B(n818),
    .Y(n1043));
 INVx1_ASAP7_75t_SL \i43/i0  (.A(n37[31]),
    .Y(n39));
 INVx1_ASAP7_75t_SL \i43/i1  (.A(n37[30]),
    .Y(n40));
 INVx1_ASAP7_75t_SL \i43/i10  (.A(n37[10]),
    .Y(n49));
 DFFHQNx1_ASAP7_75t_L \i43/i100  (.CLK(clk),
    .D(\i43/n429 ),
    .QN(n36[18]));
 SDFHx1_ASAP7_75t_SL \i43/i101  (.CLK(clk),
    .QN(n36[19]),
    .D(\i43/n95 ),
    .SE(n38),
    .SI(\i43/n331 ));
 SDFHx1_ASAP7_75t_SL \i43/i102  (.CLK(clk),
    .QN(n36[20]),
    .D(\i43/n174 ),
    .SE(n38),
    .SI(\i43/n330 ));
 SDFHx1_ASAP7_75t_SL \i43/i103  (.CLK(clk),
    .QN(n36[21]),
    .D(\i43/n115 ),
    .SE(n38),
    .SI(\i43/n328 ));
 SDFHx1_ASAP7_75t_SL \i43/i104  (.CLK(clk),
    .QN(n36[22]),
    .D(\i43/n106 ),
    .SE(n38),
    .SI(\i43/n310 ));
 SDFHx1_ASAP7_75t_SL \i43/i105  (.CLK(clk),
    .QN(n36[23]),
    .D(\i43/n136 ),
    .SE(n38),
    .SI(\i43/n326 ));
 DFFHQNx1_ASAP7_75t_SL \i43/i106  (.CLK(clk),
    .D(\i43/n428 ),
    .QN(n36[24]));
 SDFHx1_ASAP7_75t_SL \i43/i107  (.CLK(clk),
    .QN(n36[25]),
    .D(\i43/n164 ),
    .SE(n38),
    .SI(\i43/n324 ));
 SDFHx1_ASAP7_75t_SL \i43/i108  (.CLK(clk),
    .QN(n36[26]),
    .D(\i43/n112 ),
    .SE(n38),
    .SI(\i43/n61 ));
 SDFHx1_ASAP7_75t_SL \i43/i109  (.CLK(clk),
    .QN(n36[27]),
    .D(\i43/n109 ),
    .SE(n38),
    .SI(\i43/n450 ));
 INVxp33_ASAP7_75t_SL \i43/i11  (.A(n37[6]),
    .Y(n50));
 SDFHx1_ASAP7_75t_SL \i43/i110  (.CLK(clk),
    .QN(n36[28]),
    .D(\i43/n143 ),
    .SE(n38),
    .SI(\i43/n323 ));
 SDFHx1_ASAP7_75t_SL \i43/i111  (.CLK(clk),
    .QN(n36[29]),
    .D(\i43/n154 ),
    .SE(n38),
    .SI(\i43/n325 ));
 SDFHx1_ASAP7_75t_SL \i43/i112  (.CLK(clk),
    .QN(n36[30]),
    .D(\i43/n126 ),
    .SE(n38),
    .SI(\i43/n327 ));
 SDFHx1_ASAP7_75t_SL \i43/i113  (.CLK(clk),
    .QN(n36[31]),
    .D(\i43/n119 ),
    .SE(n38),
    .SI(\i43/n62 ));
 DFFHQNx1_ASAP7_75t_L \i43/i114  (.CLK(clk),
    .D(\i43/n424 ),
    .QN(n35[0]));
 SDFHx1_ASAP7_75t_SL \i43/i115  (.CLK(clk),
    .QN(n35[1]),
    .D(\i43/n142 ),
    .SE(n38),
    .SI(\i43/n316 ));
 SDFHx1_ASAP7_75t_SL \i43/i116  (.CLK(clk),
    .QN(n35[2]),
    .D(\i43/n102 ),
    .SE(n38),
    .SI(\i43/n315 ));
 SDFHx1_ASAP7_75t_SL \i43/i117  (.CLK(clk),
    .QN(n35[3]),
    .D(\i43/n149 ),
    .SE(n38),
    .SI(\i43/n314 ));
 SDFHx1_ASAP7_75t_SL \i43/i118  (.CLK(clk),
    .QN(n35[4]),
    .D(\i43/n100 ),
    .SE(n38),
    .SI(\i43/n313 ));
 SDFHx1_ASAP7_75t_SL \i43/i119  (.CLK(clk),
    .QN(n35[5]),
    .D(\i43/n116 ),
    .SE(n38),
    .SI(\i43/n59 ));
 INVx1_ASAP7_75t_SL \i43/i12  (.A(n37[5]),
    .Y(n51));
 SDFHx1_ASAP7_75t_SL \i43/i120  (.CLK(clk),
    .QN(n35[6]),
    .D(\i43/n101 ),
    .SE(n38),
    .SI(\i43/n312 ));
 SDFHx1_ASAP7_75t_SL \i43/i121  (.CLK(clk),
    .QN(n35[7]),
    .D(\i43/n93 ),
    .SE(n38),
    .SI(\i43/n311 ));
 DFFHQNx1_ASAP7_75t_L \i43/i122  (.CLK(clk),
    .D(\i43/n423 ),
    .QN(n35[8]));
 SDFHx1_ASAP7_75t_SL \i43/i123  (.CLK(clk),
    .QN(n35[9]),
    .D(\i43/n175 ),
    .SE(n38),
    .SI(\i43/n333 ));
 SDFHx1_ASAP7_75t_SL \i43/i124  (.CLK(clk),
    .QN(n35[10]),
    .D(\i43/n130 ),
    .SE(n38),
    .SI(\i43/n307 ));
 SDFHx1_ASAP7_75t_SL \i43/i125  (.CLK(clk),
    .QN(n35[11]),
    .D(\i43/n117 ),
    .SE(n38),
    .SI(\i43/n306 ));
 SDFHx1_ASAP7_75t_SL \i43/i126  (.CLK(clk),
    .QN(n35[12]),
    .D(\i43/n124 ),
    .SE(n38),
    .SI(\i43/n305 ));
 SDFHx1_ASAP7_75t_SL \i43/i127  (.CLK(clk),
    .QN(n35[13]),
    .D(\i43/n155 ),
    .SE(n38),
    .SI(\i43/n55 ));
 SDFHx1_ASAP7_75t_SL \i43/i128  (.CLK(clk),
    .QN(n35[14]),
    .D(\i43/n122 ),
    .SE(n38),
    .SI(\i43/n304 ));
 SDFHx1_ASAP7_75t_SL \i43/i129  (.CLK(clk),
    .QN(n35[15]),
    .D(\i43/n137 ),
    .SE(n38),
    .SI(\i43/n302 ));
 INVx1_ASAP7_75t_SL \i43/i13  (.A(n36[30]),
    .Y(n52));
 DFFHQNx1_ASAP7_75t_L \i43/i130  (.CLK(clk),
    .D(\i43/n422 ),
    .QN(n35[16]));
 SDFHx1_ASAP7_75t_SL \i43/i131  (.CLK(clk),
    .QN(n35[17]),
    .D(\i43/n180 ),
    .SE(n38),
    .SI(\i43/n301 ));
 SDFHx1_ASAP7_75t_SL \i43/i132  (.CLK(clk),
    .QN(n35[18]),
    .D(\i43/n110 ),
    .SE(n38),
    .SI(\i43/n299 ));
 SDFHx1_ASAP7_75t_SL \i43/i133  (.CLK(clk),
    .QN(n35[19]),
    .D(\i43/n153 ),
    .SE(n38),
    .SI(\i43/n298 ));
 SDFHx1_ASAP7_75t_SL \i43/i134  (.CLK(clk),
    .QN(n35[20]),
    .D(\i43/n132 ),
    .SE(n38),
    .SI(\i43/n300 ));
 SDFHx1_ASAP7_75t_SL \i43/i135  (.CLK(clk),
    .QN(n35[21]),
    .D(\i43/n96 ),
    .SE(n38),
    .SI(\i43/n56 ));
 SDFHx1_ASAP7_75t_SL \i43/i136  (.CLK(clk),
    .QN(n35[22]),
    .D(\i43/n157 ),
    .SE(n38),
    .SI(\i43/n303 ));
 SDFHx1_ASAP7_75t_SL \i43/i137  (.CLK(clk),
    .QN(n35[23]),
    .D(\i43/n177 ),
    .SE(n38),
    .SI(\i43/n364 ));
 SDFHx1_ASAP7_75t_SL \i43/i138  (.CLK(clk),
    .QN(n35[24]),
    .D(\i43/n141 ),
    .SE(n38),
    .SI(\i43/n420 ));
 DFFHQNx1_ASAP7_75t_L \i43/i139  (.CLK(clk),
    .D(\i43/n449 ),
    .QN(n35[25]));
 INVx1_ASAP7_75t_SL \i43/i14  (.A(n36[28]),
    .Y(n53));
 DFFHQNx1_ASAP7_75t_SL \i43/i140  (.CLK(clk),
    .D(\i43/n448 ),
    .QN(n35[26]));
 SDFHx1_ASAP7_75t_SL \i43/i141  (.CLK(clk),
    .QN(n35[27]),
    .D(\i43/n162 ),
    .SE(n38),
    .SI(\i43/n417 ));
 DFFHQNx1_ASAP7_75t_L \i43/i142  (.CLK(clk),
    .D(\i43/n447 ),
    .QN(n35[28]));
 SDFHx1_ASAP7_75t_SL \i43/i143  (.CLK(clk),
    .QN(n35[29]),
    .D(\i43/n138 ),
    .SE(n38),
    .SI(\i43/n451 ));
 DFFHQNx1_ASAP7_75t_L \i43/i144  (.CLK(clk),
    .D(\i43/n446 ),
    .QN(n35[30]));
 SDFHx1_ASAP7_75t_SL \i43/i145  (.CLK(clk),
    .QN(n35[31]),
    .D(\i43/n178 ),
    .SE(n38),
    .SI(\i43/n452 ));
 SDFHx4_ASAP7_75t_SL \i43/i146  (.CLK(clk),
    .D(\i43/n118 ),
    .QN(n34[0]),
    .SE(n38),
    .SI(\i43/n414 ));
 SDFHx4_ASAP7_75t_SL \i43/i147  (.CLK(clk),
    .D(\i43/n99 ),
    .QN(n34[1]),
    .SE(n38),
    .SI(\i43/n453 ));
 SDFHx4_ASAP7_75t_SL \i43/i148  (.CLK(clk),
    .D(\i43/n121 ),
    .QN(n34[2]),
    .SE(n38),
    .SI(\i43/n437 ));
 SDFHx4_ASAP7_75t_SL \i43/i149  (.CLK(clk),
    .D(\i43/n127 ),
    .QN(n34[3]),
    .SE(n38),
    .SI(\i43/n454 ));
 INVx1_ASAP7_75t_SL \i43/i15  (.A(n36[26]),
    .Y(n54));
 SDFHx4_ASAP7_75t_SL \i43/i150  (.CLK(clk),
    .D(\i43/n152 ),
    .QN(n34[4]),
    .SE(n38),
    .SI(\i43/n455 ));
 SDFHx4_ASAP7_75t_SL \i43/i151  (.CLK(clk),
    .D(\i43/n151 ),
    .QN(n34[5]),
    .SE(n38),
    .SI(\i43/n397 ));
 SDFHx4_ASAP7_75t_SL \i43/i152  (.CLK(clk),
    .D(\i43/n120 ),
    .QN(n34[6]),
    .SE(n38),
    .SI(\i43/n396 ));
 SDFHx4_ASAP7_75t_SL \i43/i153  (.CLK(clk),
    .D(\i43/n114 ),
    .QN(n34[7]),
    .SE(n38),
    .SI(\i43/n395 ));
 SDFHx4_ASAP7_75t_SL \i43/i154  (.CLK(clk),
    .D(\i43/n160 ),
    .QN(n34[8]),
    .SE(n38),
    .SI(\i43/n394 ));
 SDFHx4_ASAP7_75t_SL \i43/i155  (.CLK(clk),
    .D(\i43/n181 ),
    .QN(n34[9]),
    .SE(n38),
    .SI(\i43/n456 ));
 SDFHx4_ASAP7_75t_SL \i43/i156  (.CLK(clk),
    .D(\i43/n179 ),
    .QN(n34[10]),
    .SE(n38),
    .SI(\i43/n393 ));
 SDFHx4_ASAP7_75t_SL \i43/i157  (.CLK(clk),
    .D(\i43/n91 ),
    .QN(n34[11]),
    .SE(n38),
    .SI(\i43/n457 ));
 SDFHx4_ASAP7_75t_SL \i43/i158  (.CLK(clk),
    .D(\i43/n134 ),
    .QN(n34[12]),
    .SE(n38),
    .SI(\i43/n458 ));
 SDFHx4_ASAP7_75t_SL \i43/i159  (.CLK(clk),
    .D(\i43/n104 ),
    .QN(n34[13]),
    .SE(n38),
    .SI(\i43/n392 ));
 INVx1_ASAP7_75t_SL \i43/i16  (.A(n36[25]),
    .Y(n55));
 SDFHx4_ASAP7_75t_SL \i43/i160  (.CLK(clk),
    .D(\i43/n159 ),
    .QN(n34[14]),
    .SE(n38),
    .SI(\i43/n391 ));
 SDFHx4_ASAP7_75t_SL \i43/i161  (.CLK(clk),
    .D(\i43/n163 ),
    .QN(n34[15]),
    .SE(n38),
    .SI(\i43/n390 ));
 SDFHx4_ASAP7_75t_SL \i43/i162  (.CLK(clk),
    .D(\i43/n103 ),
    .QN(n34[16]),
    .SE(n38),
    .SI(\i43/n398 ));
 SDFHx4_ASAP7_75t_SL \i43/i163  (.CLK(clk),
    .D(\i43/n108 ),
    .QN(n34[17]),
    .SE(n38),
    .SI(\i43/n459 ));
 SDFHx4_ASAP7_75t_SL \i43/i164  (.CLK(clk),
    .D(\i43/n145 ),
    .QN(n34[18]),
    .SE(n38),
    .SI(\i43/n388 ));
 SDFHx4_ASAP7_75t_SL \i43/i165  (.CLK(clk),
    .D(\i43/n182 ),
    .QN(n34[19]),
    .SE(n38),
    .SI(\i43/n460 ));
 SDFHx4_ASAP7_75t_SL \i43/i166  (.CLK(clk),
    .D(\i43/n172 ),
    .QN(n34[20]),
    .SE(n38),
    .SI(\i43/n461 ));
 SDFHx4_ASAP7_75t_SL \i43/i167  (.CLK(clk),
    .D(\i43/n92 ),
    .QN(n34[21]),
    .SE(n38),
    .SI(\i43/n387 ));
 SDFHx4_ASAP7_75t_SL \i43/i168  (.CLK(clk),
    .D(\i43/n176 ),
    .QN(n34[22]),
    .SE(n38),
    .SI(\i43/n386 ));
 SDFHx4_ASAP7_75t_SL \i43/i169  (.CLK(clk),
    .D(\i43/n140 ),
    .QN(n34[23]),
    .SE(n38),
    .SI(\i43/n389 ));
 INVx1_ASAP7_75t_SL \i43/i17  (.A(n34[30]),
    .Y(n56));
 SDFHx4_ASAP7_75t_SL \i43/i170  (.CLK(clk),
    .D(\i43/n139 ),
    .QN(n34[24]),
    .SE(n38),
    .SI(\i43/n445 ));
 SDFHx4_ASAP7_75t_SL \i43/i171  (.CLK(clk),
    .D(\i43/n156 ),
    .QN(n34[25]),
    .SE(n38),
    .SI(\i43/n444 ));
 SDFHx4_ASAP7_75t_SL \i43/i172  (.CLK(clk),
    .D(\i43/n183 ),
    .QN(n34[26]),
    .SE(n38),
    .SI(\i43/n443 ));
 SDFHx4_ASAP7_75t_SL \i43/i173  (.CLK(clk),
    .D(\i43/n135 ),
    .QN(n34[27]),
    .SE(n38),
    .SI(\i43/n442 ));
 SDFHx4_ASAP7_75t_SL \i43/i174  (.CLK(clk),
    .D(\i43/n111 ),
    .QN(n34[28]),
    .SE(n38),
    .SI(\i43/n441 ));
 SDFHx4_ASAP7_75t_SL \i43/i175  (.CLK(clk),
    .D(\i43/n129 ),
    .QN(n34[29]),
    .SE(n38),
    .SI(\i43/n440 ));
 SDFHx4_ASAP7_75t_SL \i43/i176  (.CLK(clk),
    .D(\i43/n131 ),
    .QN(n34[30]),
    .SE(n38),
    .SI(\i43/n439 ));
 SDFHx4_ASAP7_75t_SL \i43/i177  (.CLK(clk),
    .D(\i43/n147 ),
    .QN(n34[31]),
    .SE(n38),
    .SI(\i43/n438 ));
 AOI22xp5_ASAP7_75t_SL \i43/i178  (.A1(n38),
    .A2(\i43/n419 ),
    .B1(net81),
    .B2(net129),
    .Y(\i43/n449 ));
 AOI22xp5_ASAP7_75t_SL \i43/i179  (.A1(n38),
    .A2(\i43/n418 ),
    .B1(net82),
    .B2(net129),
    .Y(\i43/n448 ));
 INVx1_ASAP7_75t_SL \i43/i18  (.A(n34[29]),
    .Y(n57));
 AOI22xp5_ASAP7_75t_SL \i43/i180  (.A1(n38),
    .A2(\i43/n416 ),
    .B1(net85),
    .B2(net129),
    .Y(\i43/n447 ));
 AOI22xp5_ASAP7_75t_SL \i43/i181  (.A1(n38),
    .A2(\i43/n415 ),
    .B1(net87),
    .B2(net129),
    .Y(\i43/n446 ));
 XOR2xp5_ASAP7_75t_SL \i43/i182  (.A(\i43/n69 ),
    .B(\i43/n385 ),
    .Y(\i43/n445 ));
 AOI22xp33_ASAP7_75t_SL \i43/i183  (.A1(\i43/n409 ),
    .A2(\i43/n196 ),
    .B1(\i43/n410 ),
    .B2(\i43/n195 ),
    .Y(\i43/n444 ));
 AOI22xp33_ASAP7_75t_SL \i43/i184  (.A1(\i43/n407 ),
    .A2(\i43/n194 ),
    .B1(\i43/n408 ),
    .B2(\i43/n193 ),
    .Y(\i43/n443 ));
 AOI22xp5_ASAP7_75t_SL \i43/i185  (.A1(\i43/n405 ),
    .A2(\i43/n189 ),
    .B1(\i43/n406 ),
    .B2(\i43/n188 ),
    .Y(\i43/n442 ));
 AOI22xp33_ASAP7_75t_SL \i43/i186  (.A1(\i43/n411 ),
    .A2(\i43/n185 ),
    .B1(\i43/n412 ),
    .B2(\i43/n184 ),
    .Y(\i43/n441 ));
 AOI22xp33_ASAP7_75t_SL \i43/i187  (.A1(\i43/n403 ),
    .A2(\i43/n187 ),
    .B1(\i43/n404 ),
    .B2(\i43/n186 ),
    .Y(\i43/n440 ));
 AOI22xp33_ASAP7_75t_SL \i43/i188  (.A1(\i43/n399 ),
    .A2(\i43/n191 ),
    .B1(\i43/n400 ),
    .B2(\i43/n190 ),
    .Y(\i43/n439 ));
 AOI22xp5_ASAP7_75t_SL \i43/i189  (.A1(\i43/n401 ),
    .A2(\i43/n41 ),
    .B1(\i43/n402 ),
    .B2(\i43/n192 ),
    .Y(\i43/n438 ));
 INVx1_ASAP7_75t_SL \i43/i19  (.A(n34[28]),
    .Y(n58));
 XOR2xp5_ASAP7_75t_SL \i43/i190  (.A(\i43/n348 ),
    .B(\i43/n222 ),
    .Y(\i43/n437 ));
 AOI22xp5_ASAP7_75t_SL \i43/i191  (.A1(n38),
    .A2(\i43/n317 ),
    .B1(net30),
    .B2(net129),
    .Y(\i43/n436 ));
 AOI22xp5_ASAP7_75t_L \i43/i192  (.A1(\i43/n318 ),
    .A2(n38),
    .B1(net129),
    .B2(net31),
    .Y(\i43/n435 ));
 AOI22xp5_ASAP7_75t_SL \i43/i193  (.A1(n38),
    .A2(\i43/n363 ),
    .B1(net89),
    .B2(net129),
    .Y(\i43/n434 ));
 AOI22xp5_ASAP7_75t_SL \i43/i194  (.A1(n38),
    .A2(\i43/n58 ),
    .B1(net91),
    .B2(net129),
    .Y(\i43/n433 ));
 AOI22xp5_ASAP7_75t_SL \i43/i195  (.A1(n38),
    .A2(\i43/n352 ),
    .B1(net98),
    .B2(net129),
    .Y(\i43/n432 ));
 AOI22xp5_ASAP7_75t_SL \i43/i196  (.A1(n38),
    .A2(\i43/n60 ),
    .B1(net100),
    .B2(net129),
    .Y(\i43/n431 ));
 AOI22xp5_ASAP7_75t_SL \i43/i197  (.A1(n38),
    .A2(\i43/n329 ),
    .B1(net107),
    .B2(net129),
    .Y(\i43/n430 ));
 AOI22xp5_ASAP7_75t_SL \i43/i198  (.A1(n38),
    .A2(\i43/n54 ),
    .B1(net109),
    .B2(net129),
    .Y(\i43/n429 ));
 AOI22xp5_ASAP7_75t_SL \i43/i199  (.A1(n38),
    .A2(\i43/n332 ),
    .B1(net115),
    .B2(net129),
    .Y(\i43/n428 ));
 INVx1_ASAP7_75t_SL \i43/i2  (.A(n37[29]),
    .Y(n41));
 INVxp67_ASAP7_75t_SL \i43/i20  (.A(n34[27]),
    .Y(n59));
 AOI22xp5_ASAP7_75t_SL \i43/i200  (.A1(\i43/n321 ),
    .A2(n38),
    .B1(net129),
    .B2(net27),
    .Y(\i43/n427 ));
 AOI22xp5_ASAP7_75t_SL \i43/i201  (.A1(n38),
    .A2(\i43/n319 ),
    .B1(net25),
    .B2(net129),
    .Y(\i43/n426 ));
 AOI22xp5_ASAP7_75t_SL \i43/i202  (.A1(n38),
    .A2(\i43/n322 ),
    .B1(net28),
    .B2(net129),
    .Y(\i43/n425 ));
 AOI22xp33_ASAP7_75t_SL \i43/i203  (.A1(n38),
    .A2(\i43/n337 ),
    .B1(net54),
    .B2(net129),
    .Y(\i43/n424 ));
 AOI22xp33_ASAP7_75t_SL \i43/i204  (.A1(n38),
    .A2(\i43/n339 ),
    .B1(net63),
    .B2(net129),
    .Y(\i43/n423 ));
 AOI22xp33_ASAP7_75t_SL \i43/i205  (.A1(n38),
    .A2(\i43/n335 ),
    .B1(net71),
    .B2(net129),
    .Y(\i43/n422 ));
 AOI22xp5_ASAP7_75t_SL \i43/i206  (.A1(n38),
    .A2(\i43/n340 ),
    .B1(net24),
    .B2(net129),
    .Y(\i43/n421 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i207  (.A(\i43/n243 ),
    .B(\i43/n340 ),
    .Y(\i43/n420 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i208  (.A(\i43/n346 ),
    .B(\i43/n242 ),
    .Y(\i43/n419 ));
 XOR2xp5_ASAP7_75t_SL \i43/i209  (.A(\i43/n241 ),
    .B(\i43/n462 ),
    .Y(\i43/n418 ));
 INVx1_ASAP7_75t_SL \i43/i21  (.A(n34[26]),
    .Y(n60));
 XNOR2xp5_ASAP7_75t_SL \i43/i210  (.A(\i43/n463 ),
    .B(\i43/n240 ),
    .Y(\i43/n417 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i211  (.A(\i43/n464 ),
    .B(\i43/n239 ),
    .Y(\i43/n416 ));
 XOR2xp5_ASAP7_75t_SL \i43/i212  (.A(\i43/n237 ),
    .B(\i43/n343 ),
    .Y(\i43/n415 ));
 AOI22xp5_ASAP7_75t_SL \i43/i213  (.A1(n34[0]),
    .A2(\i43/n336 ),
    .B1(n83),
    .B2(\i43/n337 ),
    .Y(\i43/n414 ));
 AOI22xp5_ASAP7_75t_SL \i43/i214  (.A1(n38),
    .A2(\i43/n309 ),
    .B1(net29),
    .B2(net129),
    .Y(\i43/n413 ));
 INVxp67_ASAP7_75t_SL \i43/i215  (.A(\i43/n411 ),
    .Y(\i43/n412 ));
 INVxp67_ASAP7_75t_SL \i43/i216  (.A(\i43/n409 ),
    .Y(\i43/n410 ));
 INVxp67_ASAP7_75t_SL \i43/i217  (.A(\i43/n407 ),
    .Y(\i43/n408 ));
 INVx1_ASAP7_75t_SL \i43/i218  (.A(\i43/n405 ),
    .Y(\i43/n406 ));
 INVxp67_ASAP7_75t_SL \i43/i219  (.A(\i43/n403 ),
    .Y(\i43/n404 ));
 INVx1_ASAP7_75t_SL \i43/i22  (.A(n34[25]),
    .Y(n61));
 INVx1_ASAP7_75t_SL \i43/i220  (.A(\i43/n401 ),
    .Y(\i43/n402 ));
 INVxp67_ASAP7_75t_SL \i43/i221  (.A(\i43/n399 ),
    .Y(\i43/n400 ));
 AOI22xp5_ASAP7_75t_SL \i43/i222  (.A1(n34[16]),
    .A2(\i43/n334 ),
    .B1(n69),
    .B2(\i43/n335 ),
    .Y(\i43/n398 ));
 XOR2xp5_ASAP7_75t_SL \i43/i223  (.A(\i43/n345 ),
    .B(\i43/n217 ),
    .Y(\i43/n397 ));
 XOR2xp5_ASAP7_75t_SL \i43/i224  (.A(\i43/n57 ),
    .B(\i43/n214 ),
    .Y(\i43/n396 ));
 XOR2xp5_ASAP7_75t_SL \i43/i225  (.A(\i43/n63 ),
    .B(\i43/n213 ),
    .Y(\i43/n395 ));
 AOI22xp5_ASAP7_75t_SL \i43/i226  (.A1(n34[8]),
    .A2(\i43/n338 ),
    .B1(n76),
    .B2(\i43/n339 ),
    .Y(\i43/n394 ));
 XOR2xp5_ASAP7_75t_SL \i43/i227  (.A(\i43/n342 ),
    .B(\i43/n207 ),
    .Y(\i43/n393 ));
 XOR2xp5_ASAP7_75t_SL \i43/i228  (.A(\i43/n341 ),
    .B(\i43/n208 ),
    .Y(\i43/n392 ));
 XOR2xp5_ASAP7_75t_SL \i43/i229  (.A(\i43/n65 ),
    .B(\i43/n215 ),
    .Y(\i43/n391 ));
 INVx1_ASAP7_75t_SL \i43/i23  (.A(n34[24]),
    .Y(n62));
 XOR2xp5_ASAP7_75t_SL \i43/i230  (.A(\i43/n64 ),
    .B(\i43/n219 ),
    .Y(\i43/n390 ));
 XOR2xp5_ASAP7_75t_SL \i43/i231  (.A(\i43/n67 ),
    .B(\i43/n265 ),
    .Y(\i43/n389 ));
 XOR2xp5_ASAP7_75t_SL \i43/i232  (.A(\i43/n347 ),
    .B(\i43/n212 ),
    .Y(\i43/n388 ));
 XOR2xp5_ASAP7_75t_SL \i43/i233  (.A(\i43/n296 ),
    .B(\i43/n211 ),
    .Y(\i43/n387 ));
 XOR2xp5_ASAP7_75t_SL \i43/i234  (.A(\i43/n66 ),
    .B(\i43/n268 ),
    .Y(\i43/n386 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i235  (.A(n34[28]),
    .B(\i43/n290 ),
    .Y(\i43/n411 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i236  (.A(n34[25]),
    .B(\i43/n291 ),
    .Y(\i43/n409 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i237  (.A(n34[26]),
    .B(\i43/n297 ),
    .Y(\i43/n407 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i238  (.A(n34[27]),
    .B(\i43/n292 ),
    .Y(\i43/n405 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i239  (.A(n34[24]),
    .B(\i43/n344 ),
    .Y(\i43/n385 ));
 INVx1_ASAP7_75t_SL \i43/i24  (.A(n34[23]),
    .Y(n63));
 XNOR2xp5_ASAP7_75t_SL \i43/i240  (.A(n34[29]),
    .B(\i43/n293 ),
    .Y(\i43/n403 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i241  (.A(n34[31]),
    .B(\i43/n295 ),
    .Y(\i43/n401 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i242  (.A(n34[30]),
    .B(\i43/n294 ),
    .Y(\i43/n399 ));
 AOI22xp33_ASAP7_75t_SL \i43/i243  (.A1(n38),
    .A2(\i43/n42 ),
    .B1(net125),
    .B2(net129),
    .Y(\i43/n384 ));
 AOI22xp33_ASAP7_75t_SL \i43/i244  (.A1(n38),
    .A2(\i43/n251 ),
    .B1(net126),
    .B2(net129),
    .Y(\i43/n383 ));
 AOI22xp33_ASAP7_75t_SL \i43/i245  (.A1(n38),
    .A2(\i43/n50 ),
    .B1(net2),
    .B2(net129),
    .Y(\i43/n382 ));
 AOI22xp33_ASAP7_75t_SL \i43/i246  (.A1(n38),
    .A2(\i43/n253 ),
    .B1(net3),
    .B2(net129),
    .Y(\i43/n381 ));
 AOI22xp33_ASAP7_75t_SL \i43/i247  (.A1(n38),
    .A2(\i43/n249 ),
    .B1(net4),
    .B2(net129),
    .Y(\i43/n380 ));
 AOI22xp33_ASAP7_75t_SL \i43/i248  (.A1(n38),
    .A2(\i43/n49 ),
    .B1(net5),
    .B2(net129),
    .Y(\i43/n379 ));
 AOI22xp5_ASAP7_75t_SL \i43/i249  (.A1(n38),
    .A2(\i43/n72 ),
    .B1(net6),
    .B2(net129),
    .Y(\i43/n378 ));
 INVx1_ASAP7_75t_SL \i43/i25  (.A(n34[22]),
    .Y(n64));
 AOI22xp33_ASAP7_75t_SL \i43/i250  (.A1(n38),
    .A2(\i43/n45 ),
    .B1(net7),
    .B2(net129),
    .Y(\i43/n377 ));
 AOI22xp33_ASAP7_75t_SL \i43/i251  (.A1(n38),
    .A2(\i43/n254 ),
    .B1(net8),
    .B2(net129),
    .Y(\i43/n376 ));
 AOI22xp33_ASAP7_75t_SL \i43/i252  (.A1(n38),
    .A2(\i43/n201 ),
    .B1(net11),
    .B2(net129),
    .Y(\i43/n375 ));
 AOI22xp33_ASAP7_75t_SL \i43/i253  (.A1(n38),
    .A2(\i43/n47 ),
    .B1(net13),
    .B2(net129),
    .Y(\i43/n374 ));
 AOI22xp33_ASAP7_75t_SL \i43/i254  (.A1(n38),
    .A2(\i43/n51 ),
    .B1(net14),
    .B2(net129),
    .Y(\i43/n373 ));
 AOI22xp33_ASAP7_75t_SL \i43/i255  (.A1(n38),
    .A2(\i43/n250 ),
    .B1(net10),
    .B2(net129),
    .Y(\i43/n372 ));
 AOI22xp5_ASAP7_75t_SL \i43/i256  (.A1(n38),
    .A2(\i43/n70 ),
    .B1(net15),
    .B2(net129),
    .Y(\i43/n371 ));
 AOI22xp33_ASAP7_75t_SL \i43/i257  (.A1(n38),
    .A2(\i43/n202 ),
    .B1(net17),
    .B2(net129),
    .Y(\i43/n370 ));
 AOI22xp33_ASAP7_75t_SL \i43/i258  (.A1(n38),
    .A2(\i43/n53 ),
    .B1(net16),
    .B2(net129),
    .Y(\i43/n369 ));
 AOI22xp33_ASAP7_75t_SL \i43/i259  (.A1(n38),
    .A2(\i43/n248 ),
    .B1(net19),
    .B2(net129),
    .Y(\i43/n368 ));
 INVxp33_ASAP7_75t_SL \i43/i26  (.A(n34[21]),
    .Y(n65));
 AOI22xp33_ASAP7_75t_SL \i43/i260  (.A1(n38),
    .A2(\i43/n204 ),
    .B1(net20),
    .B2(net129),
    .Y(\i43/n367 ));
 AOI22xp33_ASAP7_75t_SL \i43/i261  (.A1(n38),
    .A2(\i43/n43 ),
    .B1(net21),
    .B2(net129),
    .Y(\i43/n366 ));
 AOI22xp33_ASAP7_75t_SL \i43/i262  (.A1(n38),
    .A2(\i43/n52 ),
    .B1(net22),
    .B2(net129),
    .Y(\i43/n365 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i263  (.A(\i43/n265 ),
    .B(\i43/n52 ),
    .Y(\i43/n364 ));
 XOR2xp5_ASAP7_75t_SL \i43/i264  (.A(\i43/n71 ),
    .B(n36[0]),
    .Y(\i43/n363 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i265  (.A(n36[1]),
    .B(\i43/n42 ),
    .Y(\i43/n362 ));
 AOI22xp5_ASAP7_75t_SL \i43/i266  (.A1(n38),
    .A2(\i43/n71 ),
    .B1(net124),
    .B2(net129),
    .Y(\i43/n361 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i267  (.A(n36[3]),
    .B(\i43/n44 ),
    .Y(\i43/n360 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i268  (.A(n36[4]),
    .B(\i43/n50 ),
    .Y(\i43/n359 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i269  (.A(n36[5]),
    .B(\i43/n253 ),
    .Y(\i43/n358 ));
 INVx1_ASAP7_75t_SL \i43/i27  (.A(n34[20]),
    .Y(n66));
 XNOR2xp5_ASAP7_75t_SL \i43/i270  (.A(n36[6]),
    .B(\i43/n249 ),
    .Y(\i43/n357 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i271  (.A(n36[7]),
    .B(\i43/n49 ),
    .Y(\i43/n356 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i272  (.A(n36[9]),
    .B(\i43/n45 ),
    .Y(\i43/n355 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i273  (.A(n36[11]),
    .B(\i43/n48 ),
    .Y(\i43/n354 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i274  (.A(n36[12]),
    .B(\i43/n250 ),
    .Y(\i43/n353 ));
 XOR2xp5_ASAP7_75t_SL \i43/i275  (.A(\i43/n72 ),
    .B(n36[8]),
    .Y(\i43/n352 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i276  (.A(n36[13]),
    .B(\i43/n201 ),
    .Y(\i43/n351 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i277  (.A(n36[14]),
    .B(\i43/n47 ),
    .Y(\i43/n350 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i278  (.A(n36[15]),
    .B(\i43/n51 ),
    .Y(\i43/n349 ));
 AOI22xp5_ASAP7_75t_SL \i43/i279  (.A1(\i43/n274 ),
    .A2(\i43/n0 [2]),
    .B1(\i43/n273 ),
    .B2(\i43/n74 ),
    .Y(\i43/n348 ));
 INVx1_ASAP7_75t_SL \i43/i28  (.A(n34[19]),
    .Y(n67));
 AOI22xp5_ASAP7_75t_SL \i43/i280  (.A1(\i43/n230 ),
    .A2(\i43/n0 [18]),
    .B1(\i43/n229 ),
    .B2(\i43/n83 ),
    .Y(\i43/n347 ));
 XOR2xp5_ASAP7_75t_SL \i43/i281  (.A(\i43/n247 ),
    .B(\i43/n2 [25]),
    .Y(\i43/n346 ));
 OAI22xp5_ASAP7_75t_SL \i43/i282  (.A1(\i43/n270 ),
    .A2(\i43/n169 ),
    .B1(\i43/n269 ),
    .B2(\i43/n0 [5]),
    .Y(\i43/n345 ));
 XOR2xp5_ASAP7_75t_SL \i43/i283  (.A(\i43/n257 ),
    .B(n35[24]),
    .Y(\i43/n344 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i284  (.A(\i43/n2 [30]),
    .B(\i43/n245 ),
    .Y(\i43/n343 ));
 AOI22xp5_ASAP7_75t_SL \i43/i285  (.A1(\i43/n280 ),
    .A2(\i43/n0 [10]),
    .B1(\i43/n279 ),
    .B2(\i43/n87 ),
    .Y(\i43/n342 ));
 OAI22xp5_ASAP7_75t_SL \i43/i286  (.A1(\i43/n278 ),
    .A2(\i43/n171 ),
    .B1(\i43/n277 ),
    .B2(\i43/n0 [13]),
    .Y(\i43/n341 ));
 INVx1_ASAP7_75t_SL \i43/i287  (.A(\i43/n338 ),
    .Y(\i43/n339 ));
 INVx1_ASAP7_75t_SL \i43/i288  (.A(\i43/n336 ),
    .Y(\i43/n337 ));
 INVx1_ASAP7_75t_SL \i43/i289  (.A(\i43/n334 ),
    .Y(\i43/n335 ));
 INVxp67_ASAP7_75t_SL \i43/i29  (.A(n34[17]),
    .Y(n68));
 XNOR2xp5_ASAP7_75t_SL \i43/i290  (.A(\i43/n209 ),
    .B(\i43/n45 ),
    .Y(\i43/n333 ));
 XOR2xp5_ASAP7_75t_SL \i43/i291  (.A(\i43/n69 ),
    .B(\i43/n257 ),
    .Y(\i43/n332 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i292  (.A(n36[19]),
    .B(\i43/n46 ),
    .Y(\i43/n331 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i293  (.A(n36[20]),
    .B(\i43/n248 ),
    .Y(\i43/n330 ));
 XOR2xp5_ASAP7_75t_SL \i43/i294  (.A(\i43/n70 ),
    .B(n36[16]),
    .Y(\i43/n329 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i295  (.A(n36[21]),
    .B(\i43/n204 ),
    .Y(\i43/n328 ));
 AOI22xp5_ASAP7_75t_SL \i43/i296  (.A1(\i43/n260 ),
    .A2(\i43/n190 ),
    .B1(\i43/n261 ),
    .B2(\i43/n191 ),
    .Y(\i43/n327 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i297  (.A(n36[23]),
    .B(\i43/n52 ),
    .Y(\i43/n326 ));
 AOI22xp5_ASAP7_75t_SL \i43/i298  (.A1(\i43/n258 ),
    .A2(\i43/n186 ),
    .B1(\i43/n259 ),
    .B2(\i43/n187 ),
    .Y(\i43/n325 ));
 AOI22xp5_ASAP7_75t_SL \i43/i299  (.A1(\i43/n266 ),
    .A2(\i43/n195 ),
    .B1(\i43/n267 ),
    .B2(\i43/n196 ),
    .Y(\i43/n324 ));
 INVx1_ASAP7_75t_SL \i43/i3  (.A(n37[28]),
    .Y(n42));
 INVx1_ASAP7_75t_SL \i43/i30  (.A(n34[16]),
    .Y(n69));
 AOI22xp5_ASAP7_75t_SL \i43/i300  (.A1(\i43/n263 ),
    .A2(\i43/n184 ),
    .B1(\i43/n264 ),
    .B2(\i43/n185 ),
    .Y(\i43/n323 ));
 OAI22xp5_ASAP7_75t_SL \i43/i301  (.A1(n42),
    .A2(\i43/n185 ),
    .B1(n37[28]),
    .B2(\i43/n184 ),
    .Y(\i43/n322 ));
 OAI22xp5_ASAP7_75t_SL \i43/i302  (.A1(\i43/n165 ),
    .A2(\i43/n189 ),
    .B1(\i43/n188 ),
    .B2(n37[27]),
    .Y(\i43/n321 ));
 AOI22xp5_ASAP7_75t_SL \i43/i303  (.A1(n37[26]),
    .A2(\i43/n193 ),
    .B1(n43),
    .B2(\i43/n194 ),
    .Y(\i43/n320 ));
 OAI22xp5_ASAP7_75t_SL \i43/i304  (.A1(n44),
    .A2(\i43/n196 ),
    .B1(n37[25]),
    .B2(\i43/n195 ),
    .Y(\i43/n319 ));
 OAI22xp5_ASAP7_75t_SL \i43/i305  (.A1(n39),
    .A2(\i43/n41 ),
    .B1(n37[31]),
    .B2(\i43/n192 ),
    .Y(\i43/n318 ));
 OAI22xp33_ASAP7_75t_SL \i43/i306  (.A1(\i43/n191 ),
    .A2(n40),
    .B1(\i43/n190 ),
    .B2(n37[30]),
    .Y(\i43/n317 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i307  (.A(\i43/n206 ),
    .B(\i43/n42 ),
    .Y(\i43/n316 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i308  (.A(\i43/n222 ),
    .B(\i43/n251 ),
    .Y(\i43/n315 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i309  (.A(\i43/n220 ),
    .B(\i43/n44 ),
    .Y(\i43/n314 ));
 INVx1_ASAP7_75t_SL \i43/i31  (.A(n34[15]),
    .Y(n70));
 XNOR2xp5_ASAP7_75t_SL \i43/i310  (.A(\i43/n218 ),
    .B(\i43/n50 ),
    .Y(\i43/n313 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i311  (.A(\i43/n214 ),
    .B(\i43/n249 ),
    .Y(\i43/n312 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i312  (.A(\i43/n213 ),
    .B(\i43/n49 ),
    .Y(\i43/n311 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i313  (.A(n36[22]),
    .B(\i43/n43 ),
    .Y(\i43/n310 ));
 OAI22xp5_ASAP7_75t_SL \i43/i314  (.A1(n41),
    .A2(\i43/n187 ),
    .B1(n37[29]),
    .B2(\i43/n186 ),
    .Y(\i43/n309 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i315  (.A(n36[17]),
    .B(\i43/n53 ),
    .Y(\i43/n308 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i316  (.A(\i43/n207 ),
    .B(\i43/n254 ),
    .Y(\i43/n307 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i317  (.A(\i43/n223 ),
    .B(\i43/n48 ),
    .Y(\i43/n306 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i318  (.A(\i43/n205 ),
    .B(\i43/n250 ),
    .Y(\i43/n305 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i319  (.A(\i43/n215 ),
    .B(\i43/n47 ),
    .Y(\i43/n304 ));
 INVx1_ASAP7_75t_SL \i43/i32  (.A(n34[14]),
    .Y(n71));
 XNOR2xp5_ASAP7_75t_SL \i43/i320  (.A(\i43/n268 ),
    .B(\i43/n43 ),
    .Y(\i43/n303 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i321  (.A(\i43/n219 ),
    .B(\i43/n51 ),
    .Y(\i43/n302 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i322  (.A(\i43/n210 ),
    .B(\i43/n53 ),
    .Y(\i43/n301 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i323  (.A(\i43/n221 ),
    .B(\i43/n248 ),
    .Y(\i43/n300 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i324  (.A(\i43/n212 ),
    .B(\i43/n202 ),
    .Y(\i43/n299 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i325  (.A(\i43/n216 ),
    .B(\i43/n46 ),
    .Y(\i43/n298 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i326  (.A(n35[26]),
    .B(\i43/n256 ),
    .Y(\i43/n297 ));
 OAI22xp5_ASAP7_75t_SL \i43/i327  (.A1(\i43/n286 ),
    .A2(\i43/n75 ),
    .B1(\i43/n285 ),
    .B2(\i43/n0 [21]),
    .Y(\i43/n296 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i328  (.A(n35[31]),
    .B(\i43/n262 ),
    .Y(\i43/n295 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i329  (.A(n35[30]),
    .B(\i43/n261 ),
    .Y(\i43/n294 ));
 INVx1_ASAP7_75t_SL \i43/i33  (.A(n34[12]),
    .Y(n72));
 XNOR2xp5_ASAP7_75t_SL \i43/i330  (.A(n35[29]),
    .B(\i43/n259 ),
    .Y(\i43/n293 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i331  (.A(n35[27]),
    .B(\i43/n255 ),
    .Y(\i43/n292 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i332  (.A(n35[25]),
    .B(\i43/n267 ),
    .Y(\i43/n291 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i333  (.A(n35[28]),
    .B(\i43/n264 ),
    .Y(\i43/n290 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i334  (.A(n37[24]),
    .B(\i43/n69 ),
    .Y(\i43/n340 ));
 AOI22xp5_ASAP7_75t_SL \i43/i335  (.A1(\i43/n226 ),
    .A2(\i43/n199 ),
    .B1(\i43/n227 ),
    .B2(\i43/n72 ),
    .Y(\i43/n338 ));
 AOI22xp5_ASAP7_75t_SL \i43/i336  (.A1(\i43/n233 ),
    .A2(\i43/n198 ),
    .B1(\i43/n234 ),
    .B2(\i43/n71 ),
    .Y(\i43/n336 ));
 AOI22xp5_ASAP7_75t_SL \i43/i337  (.A1(\i43/n231 ),
    .A2(\i43/n197 ),
    .B1(\i43/n232 ),
    .B2(\i43/n70 ),
    .Y(\i43/n334 ));
 INVx1_ASAP7_75t_SL \i43/i338  (.A(\i43/n285 ),
    .Y(\i43/n286 ));
 INVx1_ASAP7_75t_SL \i43/i339  (.A(\i43/n279 ),
    .Y(\i43/n280 ));
 INVx1_ASAP7_75t_SL \i43/i34  (.A(n34[11]),
    .Y(n73));
 INVx1_ASAP7_75t_SL \i43/i340  (.A(\i43/n277 ),
    .Y(\i43/n278 ));
 INVx1_ASAP7_75t_SL \i43/i341  (.A(\i43/n273 ),
    .Y(\i43/n274 ));
 INVx1_ASAP7_75t_SL \i43/i342  (.A(\i43/n269 ),
    .Y(\i43/n270 ));
 INVxp67_ASAP7_75t_SL \i43/i343  (.A(\i43/n267 ),
    .Y(\i43/n266 ));
 INVxp67_ASAP7_75t_SL \i43/i344  (.A(\i43/n264 ),
    .Y(\i43/n263 ));
 INVxp67_ASAP7_75t_SL \i43/i345  (.A(\i43/n261 ),
    .Y(\i43/n260 ));
 INVxp67_ASAP7_75t_SL \i43/i346  (.A(\i43/n259 ),
    .Y(\i43/n258 ));
 INVxp67_ASAP7_75t_SL \i43/i347  (.A(\i43/n44 ),
    .Y(\i43/n252 ));
 XOR2xp5_ASAP7_75t_SL \i43/i348  (.A(n37[1]),
    .B(n34[1]),
    .Y(\i43/n289 ));
 XOR2xp5_ASAP7_75t_SL \i43/i349  (.A(n37[23]),
    .B(n34[23]),
    .Y(\i43/n288 ));
 INVx1_ASAP7_75t_SL \i43/i35  (.A(n34[10]),
    .Y(n74));
 XNOR2xp5_ASAP7_75t_SL \i43/i350  (.A(n37[25]),
    .B(n35[25]),
    .Y(\i43/n247 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i351  (.A(n41),
    .B(n35[29]),
    .Y(\i43/n246 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i352  (.A(n40),
    .B(n35[30]),
    .Y(\i43/n245 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i353  (.A(n39),
    .B(n35[31]),
    .Y(\i43/n244 ));
 XOR2xp5_ASAP7_75t_SL \i43/i354  (.A(n37[22]),
    .B(n34[22]),
    .Y(\i43/n287 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i355  (.A(n34[21]),
    .B(n37[21]),
    .Y(\i43/n285 ));
 XOR2xp5_ASAP7_75t_SL \i43/i356  (.A(n37[19]),
    .B(n34[19]),
    .Y(\i43/n284 ));
 XOR2xp5_ASAP7_75t_SL \i43/i357  (.A(n37[14]),
    .B(n34[14]),
    .Y(\i43/n283 ));
 XOR2xp5_ASAP7_75t_SL \i43/i358  (.A(n37[17]),
    .B(n34[17]),
    .Y(\i43/n282 ));
 XOR2xp5_ASAP7_75t_SL \i43/i359  (.A(n37[15]),
    .B(n34[15]),
    .Y(\i43/n281 ));
 INVx1_ASAP7_75t_SL \i43/i36  (.A(n34[9]),
    .Y(n75));
 XOR2xp5_ASAP7_75t_SL \i43/i360  (.A(n35[24]),
    .B(n36[24]),
    .Y(\i43/n243 ));
 OAI22xp5_ASAP7_75t_SL \i43/i361  (.A1(n55),
    .A2(\i43/n0 [25]),
    .B1(n36[25]),
    .B2(\i43/n73 ),
    .Y(\i43/n242 ));
 OAI22xp5_ASAP7_75t_SL \i43/i362  (.A1(n54),
    .A2(\i43/n0 [26]),
    .B1(n36[26]),
    .B2(\i43/n76 ),
    .Y(\i43/n241 ));
 OAI22xp5_ASAP7_75t_SL \i43/i363  (.A1(\i43/n168 ),
    .A2(\i43/n0 [27]),
    .B1(n36[27]),
    .B2(\i43/n86 ),
    .Y(\i43/n240 ));
 XOR2xp5_ASAP7_75t_SL \i43/i364  (.A(n37[10]),
    .B(n34[10]),
    .Y(\i43/n279 ));
 OAI22xp5_ASAP7_75t_SL \i43/i365  (.A1(n53),
    .A2(\i43/n0 [28]),
    .B1(n36[28]),
    .B2(\i43/n81 ),
    .Y(\i43/n239 ));
 OAI22xp5_ASAP7_75t_SL \i43/i366  (.A1(\i43/n166 ),
    .A2(\i43/n0 [29]),
    .B1(n36[29]),
    .B2(\i43/n90 ),
    .Y(\i43/n238 ));
 AOI22xp5_ASAP7_75t_SL \i43/i367  (.A1(n36[30]),
    .A2(\i43/n77 ),
    .B1(n52),
    .B2(\i43/n0 [30]),
    .Y(\i43/n237 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i368  (.A(n34[13]),
    .B(n37[13]),
    .Y(\i43/n277 ));
 XOR2xp5_ASAP7_75t_SL \i43/i369  (.A(\i43/n0 [31]),
    .B(n36[31]),
    .Y(\i43/n236 ));
 INVx1_ASAP7_75t_SL \i43/i37  (.A(n34[8]),
    .Y(n76));
 XOR2xp5_ASAP7_75t_SL \i43/i370  (.A(n37[11]),
    .B(n34[11]),
    .Y(\i43/n276 ));
 XOR2xp5_ASAP7_75t_SL \i43/i371  (.A(n37[9]),
    .B(n34[9]),
    .Y(\i43/n275 ));
 XOR2xp5_ASAP7_75t_SL \i43/i372  (.A(n37[2]),
    .B(n34[2]),
    .Y(\i43/n273 ));
 XOR2xp5_ASAP7_75t_SL \i43/i373  (.A(n37[3]),
    .B(n34[3]),
    .Y(\i43/n272 ));
 XOR2xp5_ASAP7_75t_SL \i43/i374  (.A(n37[7]),
    .B(n34[7]),
    .Y(\i43/n271 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i375  (.A(n34[5]),
    .B(n37[5]),
    .Y(\i43/n269 ));
 XOR2xp5_ASAP7_75t_SL \i43/i376  (.A(n35[22]),
    .B(n36[22]),
    .Y(\i43/n268 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i377  (.A(n37[25]),
    .B(n36[25]),
    .Y(\i43/n267 ));
 XOR2xp5_ASAP7_75t_SL \i43/i378  (.A(n35[23]),
    .B(n36[23]),
    .Y(\i43/n265 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i379  (.A(n37[28]),
    .B(n36[28]),
    .Y(\i43/n264 ));
 INVxp67_ASAP7_75t_R \i43/i38  (.A(n34[6]),
    .Y(n77));
 XNOR2xp5_ASAP7_75t_SL \i43/i380  (.A(n37[31]),
    .B(n36[31]),
    .Y(\i43/n262 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i381  (.A(n37[30]),
    .B(n36[30]),
    .Y(\i43/n261 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i382  (.A(n37[29]),
    .B(n36[29]),
    .Y(\i43/n259 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i383  (.A(n37[24]),
    .B(n36[24]),
    .Y(\i43/n257 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i384  (.A(n37[26]),
    .B(n36[26]),
    .Y(\i43/n256 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i385  (.A(n37[27]),
    .B(n36[27]),
    .Y(\i43/n255 ));
 OAI22xp5_ASAP7_75t_SL \i43/i386  (.A1(n49),
    .A2(\i43/n0 [10]),
    .B1(n37[10]),
    .B2(\i43/n87 ),
    .Y(\i43/n254 ));
 OAI22xp5_ASAP7_75t_SL \i43/i387  (.A1(n51),
    .A2(\i43/n0 [5]),
    .B1(n37[5]),
    .B2(\i43/n169 ),
    .Y(\i43/n253 ));
 OAI22xp5_ASAP7_75t_SL \i43/i388  (.A1(\i43/n68 ),
    .A2(\i43/n0 [2]),
    .B1(n37[2]),
    .B2(\i43/n74 ),
    .Y(\i43/n251 ));
 OAI22xp5_ASAP7_75t_SL \i43/i389  (.A1(\i43/n167 ),
    .A2(\i43/n0 [12]),
    .B1(n37[12]),
    .B2(\i43/n84 ),
    .Y(\i43/n250 ));
 INVx1_ASAP7_75t_SL \i43/i39  (.A(n34[5]),
    .Y(n78));
 OAI22xp5_ASAP7_75t_SL \i43/i390  (.A1(n50),
    .A2(\i43/n0 [6]),
    .B1(n37[6]),
    .B2(\i43/n170 ),
    .Y(\i43/n249 ));
 OAI22xp5_ASAP7_75t_SL \i43/i391  (.A1(n46),
    .A2(\i43/n0 [20]),
    .B1(n37[20]),
    .B2(\i43/n78 ),
    .Y(\i43/n248 ));
 INVx1_ASAP7_75t_SL \i43/i392  (.A(\i43/n233 ),
    .Y(\i43/n234 ));
 INVx1_ASAP7_75t_SL \i43/i393  (.A(\i43/n231 ),
    .Y(\i43/n232 ));
 INVx1_ASAP7_75t_SL \i43/i394  (.A(\i43/n229 ),
    .Y(\i43/n230 ));
 INVx1_ASAP7_75t_SL \i43/i395  (.A(\i43/n226 ),
    .Y(\i43/n227 ));
 INVxp67_ASAP7_75t_SL \i43/i396  (.A(\i43/n46 ),
    .Y(\i43/n203 ));
 INVxp67_ASAP7_75t_SL \i43/i397  (.A(\i43/n48 ),
    .Y(\i43/n200 ));
 INVx1_ASAP7_75t_SL \i43/i398  (.A(\i43/n199 ),
    .Y(\i43/n72 ));
 INVx1_ASAP7_75t_SL \i43/i399  (.A(\i43/n198 ),
    .Y(\i43/n71 ));
 INVx1_ASAP7_75t_SL \i43/i4  (.A(n37[26]),
    .Y(n43));
 INVx1_ASAP7_75t_SL \i43/i40  (.A(n34[4]),
    .Y(n79));
 INVx1_ASAP7_75t_SL \i43/i400  (.A(\i43/n197 ),
    .Y(\i43/n70 ));
 INVx2_ASAP7_75t_SL \i43/i401  (.A(\i43/n196 ),
    .Y(\i43/n195 ));
 INVx2_ASAP7_75t_SL \i43/i402  (.A(\i43/n194 ),
    .Y(\i43/n193 ));
 INVx1_ASAP7_75t_SL \i43/i403  (.A(\i43/n41 ),
    .Y(\i43/n192 ));
 INVx2_ASAP7_75t_SL \i43/i404  (.A(\i43/n191 ),
    .Y(\i43/n190 ));
 INVx1_ASAP7_75t_SL \i43/i405  (.A(\i43/n189 ),
    .Y(\i43/n188 ));
 INVx1_ASAP7_75t_SL \i43/i406  (.A(\i43/n187 ),
    .Y(\i43/n186 ));
 INVx1_ASAP7_75t_SL \i43/i407  (.A(\i43/n185 ),
    .Y(\i43/n184 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i408  (.A(n34[20]),
    .B(n46),
    .Y(\i43/n235 ));
 XOR2xp5_ASAP7_75t_SL \i43/i409  (.A(n35[0]),
    .B(n36[0]),
    .Y(\i43/n233 ));
 INVx1_ASAP7_75t_SL \i43/i41  (.A(n34[3]),
    .Y(n80));
 XOR2xp5_ASAP7_75t_SL \i43/i410  (.A(n35[16]),
    .B(n36[16]),
    .Y(\i43/n231 ));
 XOR2xp5_ASAP7_75t_SL \i43/i411  (.A(n37[18]),
    .B(n34[18]),
    .Y(\i43/n229 ));
 XOR2xp5_ASAP7_75t_SL \i43/i412  (.A(n37[4]),
    .B(n34[4]),
    .Y(\i43/n228 ));
 XOR2xp5_ASAP7_75t_SL \i43/i413  (.A(n35[8]),
    .B(n36[8]),
    .Y(\i43/n226 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i414  (.A(n34[12]),
    .B(\i43/n167 ),
    .Y(\i43/n225 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i415  (.A(n34[6]),
    .B(n50),
    .Y(\i43/n224 ));
 XOR2xp5_ASAP7_75t_SL \i43/i416  (.A(n35[11]),
    .B(n36[11]),
    .Y(\i43/n223 ));
 XOR2xp5_ASAP7_75t_SL \i43/i417  (.A(n35[2]),
    .B(n36[2]),
    .Y(\i43/n222 ));
 XOR2xp5_ASAP7_75t_SL \i43/i418  (.A(n35[20]),
    .B(n36[20]),
    .Y(\i43/n221 ));
 XOR2xp5_ASAP7_75t_SL \i43/i419  (.A(n35[3]),
    .B(n36[3]),
    .Y(\i43/n220 ));
 INVx1_ASAP7_75t_SL \i43/i42  (.A(n34[2]),
    .Y(n81));
 XOR2xp5_ASAP7_75t_SL \i43/i420  (.A(n35[15]),
    .B(n36[15]),
    .Y(\i43/n219 ));
 XOR2xp5_ASAP7_75t_SL \i43/i421  (.A(n35[4]),
    .B(n36[4]),
    .Y(\i43/n218 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i422  (.A(n36[5]),
    .B(n35[5]),
    .Y(\i43/n217 ));
 XOR2xp5_ASAP7_75t_SL \i43/i423  (.A(n35[19]),
    .B(n36[19]),
    .Y(\i43/n216 ));
 XOR2xp5_ASAP7_75t_SL \i43/i424  (.A(n35[14]),
    .B(n36[14]),
    .Y(\i43/n215 ));
 XOR2xp5_ASAP7_75t_SL \i43/i425  (.A(n35[6]),
    .B(n36[6]),
    .Y(\i43/n214 ));
 XOR2xp5_ASAP7_75t_SL \i43/i426  (.A(n35[7]),
    .B(n36[7]),
    .Y(\i43/n213 ));
 XOR2xp5_ASAP7_75t_SL \i43/i427  (.A(n35[18]),
    .B(n36[18]),
    .Y(\i43/n212 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i428  (.A(n36[21]),
    .B(n35[21]),
    .Y(\i43/n211 ));
 XOR2xp5_ASAP7_75t_SL \i43/i429  (.A(n35[17]),
    .B(n36[17]),
    .Y(\i43/n210 ));
 INVx1_ASAP7_75t_SL \i43/i43  (.A(n34[1]),
    .Y(n82));
 XOR2xp5_ASAP7_75t_SL \i43/i430  (.A(n35[9]),
    .B(n36[9]),
    .Y(\i43/n209 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i431  (.A(n36[13]),
    .B(n35[13]),
    .Y(\i43/n208 ));
 XOR2xp5_ASAP7_75t_SL \i43/i432  (.A(n35[10]),
    .B(n36[10]),
    .Y(\i43/n207 ));
 XOR2xp5_ASAP7_75t_SL \i43/i433  (.A(n35[1]),
    .B(n36[1]),
    .Y(\i43/n206 ));
 XOR2xp5_ASAP7_75t_SL \i43/i434  (.A(n35[12]),
    .B(n36[12]),
    .Y(\i43/n205 ));
 OAI22xp5_ASAP7_75t_SL \i43/i435  (.A1(n45),
    .A2(\i43/n0 [21]),
    .B1(n37[21]),
    .B2(\i43/n75 ),
    .Y(\i43/n204 ));
 OAI22xp5_ASAP7_75t_SL \i43/i436  (.A1(n47),
    .A2(\i43/n0 [18]),
    .B1(n37[18]),
    .B2(\i43/n83 ),
    .Y(\i43/n202 ));
 OAI22xp5_ASAP7_75t_SL \i43/i437  (.A1(n48),
    .A2(\i43/n0 [13]),
    .B1(n37[13]),
    .B2(\i43/n171 ),
    .Y(\i43/n201 ));
 XNOR2x1_ASAP7_75t_SL \i43/i438  (.B(n37[8]),
    .Y(\i43/n199 ),
    .A(\i43/n0 [8]));
 XNOR2x1_ASAP7_75t_SL \i43/i439  (.B(n37[0]),
    .Y(\i43/n198 ),
    .A(\i43/n0 [0]));
 INVx1_ASAP7_75t_SL \i43/i44  (.A(n34[0]),
    .Y(n83));
 XNOR2x1_ASAP7_75t_SL \i43/i440  (.B(n37[16]),
    .Y(\i43/n197 ),
    .A(\i43/n0 [16]));
 OAI22x1_ASAP7_75t_SL \i43/i441  (.A1(\i43/n85 ),
    .A2(\i43/n0 [25]),
    .B1(\i43/n2 [25]),
    .B2(\i43/n73 ),
    .Y(\i43/n196 ));
 OAI22x1_ASAP7_75t_SL \i43/i442  (.A1(\i43/n79 ),
    .A2(\i43/n0 [26]),
    .B1(\i43/n2 [26]),
    .B2(\i43/n76 ),
    .Y(\i43/n194 ));
 XNOR2x2_ASAP7_75t_SL \i43/i443  (.A(\i43/n2 [24]),
    .B(\i43/n0 [24]),
    .Y(\i43/n69 ));
 OAI22xp5_ASAP7_75t_SL \i43/i444  (.A1(\i43/n80 ),
    .A2(\i43/n0 [30]),
    .B1(\i43/n2 [30]),
    .B2(\i43/n77 ),
    .Y(\i43/n191 ));
 OAI22x1_ASAP7_75t_SL \i43/i445  (.A1(\i43/n89 ),
    .A2(\i43/n0 [27]),
    .B1(\i43/n86 ),
    .B2(\i43/n2 [27]),
    .Y(\i43/n189 ));
 OAI22x1_ASAP7_75t_SL \i43/i446  (.A1(\i43/n82 ),
    .A2(\i43/n0 [29]),
    .B1(\i43/n2 [29]),
    .B2(\i43/n90 ),
    .Y(\i43/n187 ));
 OAI22x1_ASAP7_75t_SL \i43/i447  (.A1(\i43/n88 ),
    .A2(\i43/n0 [28]),
    .B1(\i43/n2 [28]),
    .B2(\i43/n81 ),
    .Y(\i43/n185 ));
 INVxp67_ASAP7_75t_SL \i43/i448  (.A(net47),
    .Y(\i43/n183 ));
 INVxp67_ASAP7_75t_SL \i43/i449  (.A(net39),
    .Y(\i43/n182 ));
 DFFHQNx1_ASAP7_75t_SL \i43/i45/i0  (.CLK(clk),
    .D(\i43/i45/n25 ),
    .QN(\i43/n2 [29]));
 DFFHQNx1_ASAP7_75t_SL \i43/i45/i1  (.CLK(clk),
    .D(\i43/i45/n22 ),
    .QN(\i43/n2 [28]));
 A2O1A1Ixp33_ASAP7_75t_SL \i43/i45/i10  (.A1(\i43/i45/n8 ),
    .A2(\i43/i45/n14 ),
    .B(\i43/i45/n16 ),
    .C(n38),
    .Y(\i43/i45/n22 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i43/i45/i11  (.A1(\i43/i45/n6 ),
    .A2(\i43/i45/n13 ),
    .B(\i43/i45/n16 ),
    .C(n38),
    .Y(\i43/i45/n21 ));
 NAND4xp25_ASAP7_75t_SL \i43/i45/i12  (.A(\i43/i45/n14 ),
    .B(\i43/i45/n6 ),
    .C(\i43/i45/n1 [1]),
    .D(n38),
    .Y(\i43/i45/n20 ));
 AOI21xp5_ASAP7_75t_SL \i43/i45/i13  (.A1(\i43/i45/n14 ),
    .A2(\i43/i45/n9 ),
    .B(\i43/i45/n16 ),
    .Y(\i43/i45/n19 ));
 NAND4xp25_ASAP7_75t_SL \i43/i45/i14  (.A(\i43/i45/n14 ),
    .B(\i43/i45/n7 ),
    .C(\i43/i45/n1 [0]),
    .D(n38),
    .Y(\i43/i45/n18 ));
 AND2x2_ASAP7_75t_SL \i43/i45/i15  (.A(\i43/i45/n6 ),
    .B(\i43/i45/n16 ),
    .Y(\i43/i45/n17 ));
 AND2x2_ASAP7_75t_SL \i43/i45/i16  (.A(\i43/i45/n0 [3]),
    .B(\i43/i45/n13 ),
    .Y(\i43/i45/n16 ));
 NOR3xp33_ASAP7_75t_SL \i43/i45/i17  (.A(\i43/i45/n0 [3]),
    .B(\i43/i45/n26 ),
    .C(\i43/i45/n9 ),
    .Y(\i43/i45/n15 ));
 NOR2xp33_ASAP7_75t_SL \i43/i45/i18  (.A(\i43/i45/n11 ),
    .B(\i43/i45/n0 [3]),
    .Y(\i43/i45/n14 ));
 DFFHQNx1_ASAP7_75t_SL \i43/i45/i19  (.CLK(clk),
    .D(\i43/i45/n10 ),
    .QN(\i43/n2 [24]));
 DFFHQNx1_ASAP7_75t_SL \i43/i45/i2  (.CLK(clk),
    .D(\i43/i45/n24 ),
    .QN(\i43/n2 [27]));
 NOR2xp33_ASAP7_75t_SL \i43/i45/i20  (.A(\i43/i45/n0 [1]),
    .B(\i43/i45/n26 ),
    .Y(\i43/i45/n13 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i45/i21  (.A(\i43/i45/n1 [3]),
    .B(\i43/i45/n27 ),
    .Y(\i43/i45/n0 [3]));
 NOR2xp33_ASAP7_75t_SL \i43/i45/i22  (.A(\i43/i45/n1 [3]),
    .B(\i43/i45/n27 ),
    .Y(\i43/i45/n12 ));
 AND2x2_ASAP7_75t_SL \i43/i45/i23  (.A(n38),
    .B(\i43/i45/n27 ),
    .Y(\i43/i45/n10 ));
 INVxp67_ASAP7_75t_SL \i43/i45/i24  (.A(\i43/i45/n0 [1]),
    .Y(\i43/i45/n9 ));
 AOI21xp5_ASAP7_75t_SL \i43/i45/i25  (.A1(\i43/i45/n7 ),
    .A2(\i43/i45/n6 ),
    .B(\i43/i45/n8 ),
    .Y(\i43/i45/n0 [1]));
 AND2x2_ASAP7_75t_SL \i43/i45/i26  (.A(\i43/i45/n1 [0]),
    .B(\i43/i45/n1 [1]),
    .Y(\i43/i45/n8 ));
 INVxp67_ASAP7_75t_SL \i43/i45/i27  (.A(\i43/i45/n1 [1]),
    .Y(\i43/i45/n7 ));
 INVx1_ASAP7_75t_SL \i43/i45/i28  (.A(\i43/i45/n1 [0]),
    .Y(\i43/i45/n6 ));
 DFFHQNx1_ASAP7_75t_SL \i43/i45/i29  (.CLK(clk),
    .D(\i43/i45/n3 ),
    .QN(\i43/i45/n1 [2]));
 DFFHQNx1_ASAP7_75t_SL \i43/i45/i3  (.CLK(clk),
    .D(\i43/i45/n23 ),
    .QN(\i43/n2 [26]));
 DFFHQNx1_ASAP7_75t_L \i43/i45/i30  (.CLK(clk),
    .D(\i43/i45/n2 ),
    .QN(\i43/i45/n1 [0]));
 DFFHQNx1_ASAP7_75t_SL \i43/i45/i31  (.CLK(clk),
    .D(\i43/i45/n5 ),
    .QN(\i43/i45/n1 [3]));
 DFFHQNx1_ASAP7_75t_SL \i43/i45/i32  (.CLK(clk),
    .D(\i43/i45/n4 ),
    .QN(\i43/i45/n1 [1]));
 NAND2xp5_ASAP7_75t_SL \i43/i45/i33  (.A(n38),
    .B(\i43/i45/n0 [3]),
    .Y(\i43/i45/n5 ));
 NAND2xp5_ASAP7_75t_SL \i43/i45/i34  (.A(n38),
    .B(\i43/i45/n0 [1]),
    .Y(\i43/i45/n4 ));
 NAND2xp5_ASAP7_75t_SL \i43/i45/i35  (.A(n38),
    .B(\i43/i45/n26 ),
    .Y(\i43/i45/n3 ));
 OR2x2_ASAP7_75t_SL \i43/i45/i36  (.A(net129),
    .B(\i43/i45/n1 [0]),
    .Y(\i43/i45/n2 ));
 INVxp33_ASAP7_75t_SL \i43/i45/i37  (.A(\i43/i45/n11 ),
    .Y(\i43/i45/n26 ));
 HAxp5_ASAP7_75t_SL \i43/i45/i38  (.A(\i43/i45/n8 ),
    .B(\i43/i45/n1 [2]),
    .CON(\i43/i45/n27 ),
    .SN(\i43/i45/n11 ));
 OR3x1_ASAP7_75t_SL \i43/i45/i4  (.A(\i43/i45/n19 ),
    .B(\i43/i45/n1 [0]),
    .C(net129),
    .Y(\i43/i45/n25 ));
 DFFHQNx1_ASAP7_75t_SL \i43/i45/i5  (.CLK(clk),
    .D(\i43/i45/n21 ),
    .QN(\i43/n2 [25]));
 DFFHQNx1_ASAP7_75t_SL \i43/i45/i6  (.CLK(clk),
    .D(\i43/i45/n18 ),
    .QN(\i43/n2 [30]));
 DFFHQNx1_ASAP7_75t_SL \i43/i45/i7  (.CLK(clk),
    .D(\i43/i45/n20 ),
    .QN(\i43/n2 [31]));
 A2O1A1Ixp33_ASAP7_75t_SL \i43/i45/i8  (.A1(\i43/i45/n6 ),
    .A2(\i43/i45/n15 ),
    .B(\i43/i45/n12 ),
    .C(n38),
    .Y(\i43/i45/n24 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i43/i45/i9  (.A1(\i43/i45/n1 [0]),
    .A2(\i43/i45/n15 ),
    .B(\i43/i45/n17 ),
    .C(n38),
    .Y(\i43/i45/n23 ));
 INVxp67_ASAP7_75t_SL \i43/i450  (.A(net128),
    .Y(\i43/n181 ));
 INVxp67_ASAP7_75t_SL \i43/i451  (.A(net72),
    .Y(\i43/n180 ));
 INVxp67_ASAP7_75t_SL \i43/i452  (.A(net12),
    .Y(\i43/n179 ));
 INVxp67_ASAP7_75t_SL \i43/i453  (.A(net88),
    .Y(\i43/n178 ));
 INVxp67_ASAP7_75t_SL \i43/i454  (.A(net79),
    .Y(\i43/n177 ));
 INVxp67_ASAP7_75t_SL \i43/i455  (.A(net43),
    .Y(\i43/n176 ));
 INVxp67_ASAP7_75t_SL \i43/i456  (.A(net64),
    .Y(\i43/n175 ));
 INVxp67_ASAP7_75t_SL \i43/i457  (.A(net111),
    .Y(\i43/n174 ));
 INVxp67_ASAP7_75t_SL \i43/i458  (.A(net99),
    .Y(\i43/n173 ));
 INVxp67_ASAP7_75t_SL \i43/i459  (.A(net41),
    .Y(\i43/n172 ));
 NOR2x1_ASAP7_75t_SL \i43/i46/i0  (.A(\i43/i46/n488 ),
    .B(\i43/i46/n514 ),
    .Y(\i43/n0 [25]));
 AND3x2_ASAP7_75t_SL \i43/i46/i1  (.A(\i43/i46/n510 ),
    .B(\i43/i46/n512 ),
    .C(\i43/i46/n492 ),
    .Y(\i43/n0 [29]));
 NOR4xp75_ASAP7_75t_SL \i43/i46/i10  (.A(\i43/i46/n500 ),
    .B(\i43/i46/n504 ),
    .C(\i43/i46/n482 ),
    .D(\i43/i46/n497 ),
    .Y(\i43/n0 [26]));
 INVx1_ASAP7_75t_SL \i43/i46/i100  (.A(\i43/i46/n420 ),
    .Y(\i43/i46/n421 ));
 INVx1_ASAP7_75t_SL \i43/i46/i101  (.A(\i43/i46/n418 ),
    .Y(\i43/i46/n419 ));
 INVx1_ASAP7_75t_SL \i43/i46/i102  (.A(\i43/i46/n415 ),
    .Y(\i43/i46/n416 ));
 INVx1_ASAP7_75t_SL \i43/i46/i103  (.A(\i43/i46/n413 ),
    .Y(\i43/i46/n414 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i104  (.A(\i43/i46/n359 ),
    .B(\i43/i46/n354 ),
    .Y(\i43/i46/n412 ));
 NOR3xp33_ASAP7_75t_SL \i43/i46/i105  (.A(\i43/i46/n280 ),
    .B(\i43/i46/n249 ),
    .C(\i43/i46/n227 ),
    .Y(\i43/i46/n411 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i106  (.A(\i43/i46/n327 ),
    .B(\i43/i46/n323 ),
    .Y(\i43/i46/n410 ));
 NAND2xp5_ASAP7_75t_L \i43/i46/i107  (.A(\i43/i46/n372 ),
    .B(\i43/i46/n326 ),
    .Y(\i43/i46/n409 ));
 NAND3xp33_ASAP7_75t_L \i43/i46/i108  (.A(\i43/i46/n269 ),
    .B(\i43/i46/n275 ),
    .C(\i43/i46/n357 ),
    .Y(\i43/i46/n408 ));
 NAND2xp5_ASAP7_75t_L \i43/i46/i109  (.A(\i43/i46/n339 ),
    .B(\i43/i46/n214 ),
    .Y(\i43/i46/n407 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i11  (.A(\i43/i46/n483 ),
    .B(\i43/i46/n499 ),
    .Y(\i43/i46/n512 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i110  (.A(\i43/i46/n360 ),
    .B(\i43/i46/n333 ),
    .Y(\i43/i46/n406 ));
 NAND5xp2_ASAP7_75t_SL \i43/i46/i111  (.A(\i43/i46/n298 ),
    .B(\i43/i46/n120 ),
    .C(\i43/i46/n182 ),
    .D(\i43/i46/n123 ),
    .E(\i43/i46/n117 ),
    .Y(\i43/i46/n405 ));
 NOR4xp25_ASAP7_75t_SL \i43/i46/i112  (.A(\i43/i46/n281 ),
    .B(\i43/i46/n197 ),
    .C(\i43/i46/n132 ),
    .D(\i43/i46/n226 ),
    .Y(\i43/i46/n404 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i113  (.A(\i43/i46/n350 ),
    .B(\i43/i46/n362 ),
    .Y(\i43/i46/n403 ));
 NAND2xp33_ASAP7_75t_SL \i43/i46/i114  (.A(\i43/i46/n322 ),
    .B(\i43/i46/n305 ),
    .Y(\i43/i46/n402 ));
 AOI221xp5_ASAP7_75t_SL \i43/i46/i115  (.A1(\i43/i46/n109 ),
    .A2(\i43/i46/n95 ),
    .B1(\i43/i46/n115 ),
    .B2(\i43/i46/n47 ),
    .C(\i43/i46/n216 ),
    .Y(\i43/i46/n423 ));
 NAND5xp2_ASAP7_75t_SL \i43/i46/i116  (.A(\i43/i46/n279 ),
    .B(\i43/i46/n206 ),
    .C(\i43/i46/n211 ),
    .D(\i43/i46/n182 ),
    .E(\i43/i46/n122 ),
    .Y(\i43/i46/n401 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i117  (.A(\i43/i46/n295 ),
    .B(\i43/i46/n372 ),
    .Y(\i43/i46/n400 ));
 OAI221xp5_ASAP7_75t_SL \i43/i46/i118  (.A1(\i43/i46/n157 ),
    .A2(\i43/i46/n54 ),
    .B1(\i43/i46/n158 ),
    .B2(\i43/i46/n39 ),
    .C(\i43/i46/n338 ),
    .Y(\i43/i46/n399 ));
 NOR2xp33_ASAP7_75t_L \i43/i46/i119  (.A(\i43/i46/n292 ),
    .B(\i43/i46/n359 ),
    .Y(\i43/i46/n422 ));
 NAND3xp33_ASAP7_75t_SL \i43/i46/i12  (.A(\i43/i46/n486 ),
    .B(\i43/i46/n423 ),
    .C(\i43/i46/n491 ),
    .Y(\i43/i46/n511 ));
 AND2x2_ASAP7_75t_SL \i43/i46/i120  (.A(\i43/i46/n289 ),
    .B(\i43/i46/n321 ),
    .Y(\i43/i46/n420 ));
 NOR3xp33_ASAP7_75t_SL \i43/i46/i121  (.A(\i43/i46/n218 ),
    .B(\i43/i46/n227 ),
    .C(\i43/i46/n196 ),
    .Y(\i43/i46/n418 ));
 NAND3xp33_ASAP7_75t_SL \i43/i46/i122  (.A(\i43/i46/n334 ),
    .B(\i43/i46/n285 ),
    .C(\i43/i46/n239 ),
    .Y(\i43/i46/n417 ));
 NAND2x1_ASAP7_75t_SL \i43/i46/i123  (.A(\i43/i46/n215 ),
    .B(\i43/i46/n300 ),
    .Y(\i43/i46/n415 ));
 NOR3xp33_ASAP7_75t_SL \i43/i46/i124  (.A(\i43/i46/n288 ),
    .B(\i43/i46/n232 ),
    .C(\i43/i46/n272 ),
    .Y(\i43/i46/n413 ));
 INVx1_ASAP7_75t_SL \i43/i46/i125  (.A(\i43/i46/n391 ),
    .Y(\i43/i46/n392 ));
 OAI21xp33_ASAP7_75t_SL \i43/i46/i126  (.A1(\i43/i46/n76 ),
    .A2(\i43/i46/n45 ),
    .B(\i43/i46/n370 ),
    .Y(\i43/i46/n390 ));
 NOR3xp33_ASAP7_75t_SL \i43/i46/i127  (.A(\i43/i46/n329 ),
    .B(\i43/i46/n192 ),
    .C(\i43/i46/n232 ),
    .Y(\i43/i46/n389 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i128  (.A1(\i43/i46/n87 ),
    .A2(\i43/i46/n50 ),
    .B(\i43/i46/n357 ),
    .Y(\i43/i46/n398 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i129  (.A1(\i43/i46/n41 ),
    .A2(\i43/i46/n270 ),
    .B(\i43/i46/n265 ),
    .Y(\i43/i46/n388 ));
 NOR3xp33_ASAP7_75t_SL \i43/i46/i13  (.A(\i43/i46/n480 ),
    .B(\i43/i46/n487 ),
    .C(\i43/i46/n464 ),
    .Y(\i43/i46/n510 ));
 NAND4xp25_ASAP7_75t_SL \i43/i46/i130  (.A(\i43/i46/n245 ),
    .B(\i43/i46/n146 ),
    .C(\i43/i46/n96 ),
    .D(\i43/i46/n99 ),
    .Y(\i43/i46/n387 ));
 NAND5xp2_ASAP7_75t_SL \i43/i46/i131  (.A(\i43/i46/n209 ),
    .B(\i43/i46/n120 ),
    .C(\i43/i46/n165 ),
    .D(\i43/i46/n185 ),
    .E(\i43/i46/n141 ),
    .Y(\i43/i46/n386 ));
 AOI211xp5_ASAP7_75t_SL \i43/i46/i132  (.A1(\i43/i46/n41 ),
    .A2(\i43/i46/n62 ),
    .B(\i43/i46/n284 ),
    .C(\i43/i46/n283 ),
    .Y(\i43/i46/n385 ));
 NOR3xp33_ASAP7_75t_SL \i43/i46/i133  (.A(\i43/i46/n294 ),
    .B(\i43/i46/n207 ),
    .C(\i43/i46/n222 ),
    .Y(\i43/i46/n384 ));
 NOR2xp33_ASAP7_75t_L \i43/i46/i134  (.A(\i43/i46/n336 ),
    .B(\i43/i46/n317 ),
    .Y(\i43/i46/n383 ));
 OAI221xp5_ASAP7_75t_SL \i43/i46/i135  (.A1(\i43/i46/n271 ),
    .A2(\i43/i46/n75 ),
    .B1(\i43/i46/n174 ),
    .B2(\i43/i46/n72 ),
    .C(\i43/i46/n89 ),
    .Y(\i43/i46/n382 ));
 NAND3xp33_ASAP7_75t_SL \i43/i46/i136  (.A(\i43/i46/n290 ),
    .B(\i43/i46/n279 ),
    .C(\i43/i46/n221 ),
    .Y(\i43/i46/n381 ));
 NAND5xp2_ASAP7_75t_SL \i43/i46/i137  (.A(\i43/i46/n247 ),
    .B(\i43/i46/n176 ),
    .C(\i43/i46/n105 ),
    .D(\i43/i46/n113 ),
    .E(\i43/i46/n145 ),
    .Y(\i43/i46/n380 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i138  (.A1(\i43/i46/n45 ),
    .A2(\i43/i46/n40 ),
    .B(\i43/i46/n360 ),
    .Y(\i43/i46/n379 ));
 NOR4xp25_ASAP7_75t_SL \i43/i46/i139  (.A(\i43/i46/n335 ),
    .B(\i43/i46/n268 ),
    .C(\i43/i46/n97 ),
    .D(\i43/i46/n98 ),
    .Y(\i43/i46/n378 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i14  (.A(\i43/i46/n501 ),
    .B(\i43/i46/n490 ),
    .Y(\i43/i46/n509 ));
 OAI211xp5_ASAP7_75t_SL \i43/i46/i140  (.A1(\i43/i46/n40 ),
    .A2(\i43/i46/n261 ),
    .B(\i43/i46/n180 ),
    .C(\i43/i46/n168 ),
    .Y(\i43/i46/n377 ));
 NAND5xp2_ASAP7_75t_SL \i43/i46/i141  (.A(\i43/i46/n258 ),
    .B(\i43/i46/n243 ),
    .C(\i43/i46/n118 ),
    .D(\i43/i46/n181 ),
    .E(\i43/i46/n186 ),
    .Y(\i43/i46/n376 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i142  (.A(\i43/i46/n332 ),
    .B(\i43/i46/n303 ),
    .Y(\i43/i46/n375 ));
 OAI221xp5_ASAP7_75t_SL \i43/i46/i143  (.A1(\i43/i46/n262 ),
    .A2(\i43/i46/n54 ),
    .B1(\i43/i46/n52 ),
    .B2(\i43/i46/n87 ),
    .C(\i43/i46/n223 ),
    .Y(\i43/i46/n374 ));
 NOR3xp33_ASAP7_75t_SL \i43/i46/i144  (.A(\i43/i46/n309 ),
    .B(\i43/i46/n276 ),
    .C(\i43/i46/n274 ),
    .Y(\i43/i46/n397 ));
 NOR2x1_ASAP7_75t_SL \i43/i46/i145  (.A(\i43/i46/n241 ),
    .B(\i43/i46/n361 ),
    .Y(\i43/i46/n396 ));
 OA211x2_ASAP7_75t_SL \i43/i46/i146  (.A1(\i43/i46/n92 ),
    .A2(\i43/i46/n54 ),
    .B(\i43/i46/n369 ),
    .C(\i43/i46/n147 ),
    .Y(\i43/i46/n395 ));
 NOR2xp33_ASAP7_75t_L \i43/i46/i147  (.A(\i43/i46/n191 ),
    .B(\i43/i46/n318 ),
    .Y(\i43/i46/n394 ));
 NOR2xp33_ASAP7_75t_L \i43/i46/i148  (.A(\i43/i46/n201 ),
    .B(\i43/i46/n365 ),
    .Y(\i43/i46/n393 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i149  (.A(\i43/i46/n304 ),
    .B(\i43/i46/n344 ),
    .Y(\i43/i46/n391 ));
 NAND3xp33_ASAP7_75t_SL \i43/i46/i15  (.A(\i43/i46/n475 ),
    .B(\i43/i46/n485 ),
    .C(\i43/i46/n463 ),
    .Y(\i43/i46/n508 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i150  (.A(\i43/i46/n367 ),
    .Y(\i43/i46/n368 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i151  (.A(\i43/i46/n365 ),
    .Y(\i43/i46/n366 ));
 INVx1_ASAP7_75t_SL \i43/i46/i152  (.A(\i43/i46/n363 ),
    .Y(\i43/i46/n364 ));
 INVx1_ASAP7_75t_SL \i43/i46/i153  (.A(\i43/i46/n361 ),
    .Y(\i43/i46/n362 ));
 INVx1_ASAP7_75t_SL \i43/i46/i154  (.A(\i43/i46/n519 ),
    .Y(\i43/i46/n355 ));
 NAND2xp33_ASAP7_75t_L \i43/i46/i155  (.A(\i43/i46/n215 ),
    .B(\i43/i46/n273 ),
    .Y(\i43/i46/n354 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i156  (.A(\i43/i46/n131 ),
    .B(\i43/i46/n221 ),
    .Y(\i43/i46/n353 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i157  (.A(\i43/i46/n193 ),
    .B(\i43/i46/n213 ),
    .Y(\i43/i46/n352 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i46/i158  (.A1(\i43/i46/n34 ),
    .A2(\i43/i46/n65 ),
    .B(\i43/i46/n33 ),
    .C(\i43/i46/n228 ),
    .Y(\i43/i46/n351 ));
 OAI31xp33_ASAP7_75t_SL \i43/i46/i159  (.A1(\i43/i46/n65 ),
    .A2(\i43/i46/n41 ),
    .A3(\i43/i46/n55 ),
    .B(\i43/i46/n79 ),
    .Y(\i43/i46/n350 ));
 NOR2x1_ASAP7_75t_SL \i43/i46/i16  (.A(\i43/i46/n474 ),
    .B(\i43/i46/n470 ),
    .Y(\i43/i46/n505 ));
 NAND3xp33_ASAP7_75t_SL \i43/i46/i160  (.A(\i43/i46/n214 ),
    .B(\i43/i46/n184 ),
    .C(\i43/i46/n129 ),
    .Y(\i43/i46/n349 ));
 AOI21xp5_ASAP7_75t_SL \i43/i46/i161  (.A1(\i43/i46/n38 ),
    .A2(\i43/i46/n74 ),
    .B(\i43/i46/n1 ),
    .Y(\i43/i46/n348 ));
 AOI211xp5_ASAP7_75t_SL \i43/i46/i162  (.A1(\i43/i46/n57 ),
    .A2(\i43/i46/n71 ),
    .B(\i43/i46/n183 ),
    .C(\i43/i46/n121 ),
    .Y(\i43/i46/n373 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i163  (.A1(\i43/i46/n94 ),
    .A2(\i43/i46/n58 ),
    .B(\i43/i46/n217 ),
    .Y(\i43/i46/n347 ));
 OAI31xp33_ASAP7_75t_SL \i43/i46/i164  (.A1(\i43/i46/n47 ),
    .A2(\i43/i46/n95 ),
    .A3(\i43/i46/n51 ),
    .B(\i43/i46/n69 ),
    .Y(\i43/i46/n346 ));
 AO21x1_ASAP7_75t_SL \i43/i46/i165  (.A1(\i43/i46/n67 ),
    .A2(\i43/i46/n151 ),
    .B(\i43/i46/n282 ),
    .Y(\i43/i46/n345 ));
 NOR2xp33_ASAP7_75t_L \i43/i46/i166  (.A(\i43/i46/n229 ),
    .B(\i43/i46/n260 ),
    .Y(\i43/i46/n344 ));
 AO21x1_ASAP7_75t_SL \i43/i46/i167  (.A1(\i43/i46/n149 ),
    .A2(\i43/i46/n174 ),
    .B(\i43/i46/n76 ),
    .Y(\i43/i46/n343 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i43/i46/i168  (.A1(\i43/i46/n70 ),
    .A2(\i43/i46/n78 ),
    .B(\i43/i46/n52 ),
    .C(\i43/i46/n198 ),
    .Y(\i43/i46/n342 ));
 AOI21xp5_ASAP7_75t_SL \i43/i46/i169  (.A1(\i43/i46/n44 ),
    .A2(\i43/i46/n67 ),
    .B(\i43/i46/n220 ),
    .Y(\i43/i46/n341 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i17  (.A(\i43/i46/n476 ),
    .B(\i43/i46/n485 ),
    .Y(\i43/i46/n504 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i43/i46/i170  (.A1(\i43/i46/n42 ),
    .A2(\i43/i46/n35 ),
    .B(\i43/i46/n87 ),
    .C(\i43/i46/n117 ),
    .Y(\i43/i46/n340 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i171  (.A(\i43/i46/n250 ),
    .B(\i43/i46/n237 ),
    .Y(\i43/i46/n339 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i46/i172  (.A1(\i43/i46/n77 ),
    .A2(\i43/i46/n51 ),
    .B(\i43/i46/n33 ),
    .C(\i43/i46/n133 ),
    .Y(\i43/i46/n338 ));
 NAND3xp33_ASAP7_75t_SL \i43/i46/i173  (.A(\i43/i46/n233 ),
    .B(\i43/i46/n173 ),
    .C(\i43/i46/n138 ),
    .Y(\i43/i46/n337 ));
 OAI221xp5_ASAP7_75t_SL \i43/i46/i174  (.A1(\i43/i46/n75 ),
    .A2(\i43/i46/n56 ),
    .B1(\i43/i46/n49 ),
    .B2(\i43/i46/n68 ),
    .C(\i43/i46/n135 ),
    .Y(\i43/i46/n336 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i175  (.A1(\i43/i46/n78 ),
    .A2(\i43/i46/n137 ),
    .B(\i43/i46/n238 ),
    .Y(\i43/i46/n335 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i176  (.A(\i43/i46/n234 ),
    .B(\i43/i46/n210 ),
    .Y(\i43/i46/n334 ));
 AOI221xp5_ASAP7_75t_SL \i43/i46/i177  (.A1(\i43/i46/n34 ),
    .A2(\i43/i46/n79 ),
    .B1(\i43/i46/n67 ),
    .B2(\i43/i46/n83 ),
    .C(\i43/i46/n237 ),
    .Y(\i43/i46/n333 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i178  (.A1(\i43/i46/n59 ),
    .A2(\i43/i46/n155 ),
    .B(\i43/i46/n77 ),
    .Y(\i43/i46/n332 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i46/i179  (.A1(\i43/i46/n62 ),
    .A2(\i43/i46/n44 ),
    .B(\i43/i46/n57 ),
    .C(\i43/i46/n126 ),
    .Y(\i43/i46/n331 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i18  (.A(\i43/i46/n481 ),
    .B(\i43/i46/n473 ),
    .Y(\i43/i46/n503 ));
 OAI221xp5_ASAP7_75t_SL \i43/i46/i180  (.A1(\i43/i46/n46 ),
    .A2(\i43/i46/n87 ),
    .B1(\i43/i46/n52 ),
    .B2(\i43/i46/n80 ),
    .C(\i43/i46/n163 ),
    .Y(\i43/i46/n330 ));
 AOI21xp5_ASAP7_75t_SL \i43/i46/i181  (.A1(\i43/i46/n95 ),
    .A2(\i43/i46/n62 ),
    .B(\i43/i46/n1 ),
    .Y(\i43/i46/n372 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i182  (.A(\i43/i46/n220 ),
    .B(\i43/i46/n252 ),
    .Y(\i43/i46/n371 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i183  (.A(\i43/i46/n254 ),
    .B(\i43/i46/n0 ),
    .Y(\i43/i46/n370 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i184  (.A(\i43/i46/n226 ),
    .B(\i43/i46/n195 ),
    .Y(\i43/i46/n369 ));
 OAI211xp5_ASAP7_75t_SL \i43/i46/i185  (.A1(\i43/i46/n63 ),
    .A2(\i43/i46/n46 ),
    .B(\i43/i46/n177 ),
    .C(\i43/i46/n187 ),
    .Y(\i43/i46/n367 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i186  (.A(\i43/i46/n120 ),
    .B(\i43/i46/n246 ),
    .Y(\i43/i46/n365 ));
 AOI222xp33_ASAP7_75t_SL \i43/i46/i187  (.A1(\i43/i46/n85 ),
    .A2(\i43/i46/n41 ),
    .B1(\i43/i46/n59 ),
    .B2(\i43/i46/n38 ),
    .C1(\i43/i46/n69 ),
    .C2(\i43/i46/n47 ),
    .Y(\i43/i46/n363 ));
 OAI221xp5_ASAP7_75t_SL \i43/i46/i188  (.A1(\i43/i46/n45 ),
    .A2(\i43/i46/n35 ),
    .B1(\i43/i46/n37 ),
    .B2(\i43/i46/n52 ),
    .C(\i43/i46/n180 ),
    .Y(\i43/i46/n361 ));
 AOI222xp33_ASAP7_75t_SL \i43/i46/i189  (.A1(\i43/i46/n34 ),
    .A2(\i43/i46/n90 ),
    .B1(\i43/i46/n33 ),
    .B2(\i43/i46/n67 ),
    .C1(\i43/i46/n83 ),
    .C2(\i43/i46/n73 ),
    .Y(\i43/i46/n360 ));
 NOR4xp75_ASAP7_75t_SL \i43/i46/i19  (.A(\i43/i46/n436 ),
    .B(\i43/i46/n400 ),
    .C(\i43/i46/n375 ),
    .D(\i43/i46/n374 ),
    .Y(\i43/i46/n502 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i190  (.A1(\i43/i46/n39 ),
    .A2(\i43/i46/n91 ),
    .B(\i43/i46/n238 ),
    .Y(\i43/i46/n359 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i191  (.A(\i43/i46/n205 ),
    .B(\i43/i46/n228 ),
    .Y(\i43/i46/n358 ));
 NOR2xp33_ASAP7_75t_L \i43/i46/i192  (.A(\i43/i46/n256 ),
    .B(\i43/i46/n281 ),
    .Y(\i43/i46/n357 ));
 NOR2x1_ASAP7_75t_SL \i43/i46/i193  (.A(\i43/i46/n142 ),
    .B(\i43/i46/n280 ),
    .Y(\i43/i46/n356 ));
 INVxp33_ASAP7_75t_SL \i43/i46/i194  (.A(\i43/i46/n326 ),
    .Y(\i43/i46/n327 ));
 INVx1_ASAP7_75t_SL \i43/i46/i195  (.A(\i43/i46/n323 ),
    .Y(\i43/i46/n324 ));
 INVx1_ASAP7_75t_SL \i43/i46/i196  (.A(\i43/i46/n318 ),
    .Y(\i43/i46/n319 ));
 OAI211xp5_ASAP7_75t_SL \i43/i46/i197  (.A1(\i43/i46/n40 ),
    .A2(\i43/i46/n70 ),
    .B(\i43/i46/n189 ),
    .C(\i43/i46/n188 ),
    .Y(\i43/i46/n317 ));
 AO21x1_ASAP7_75t_SL \i43/i46/i198  (.A1(\i43/i46/n67 ),
    .A2(\i43/i46/n0 ),
    .B(\i43/i46/n225 ),
    .Y(\i43/i46/n316 ));
 OAI221xp5_ASAP7_75t_SL \i43/i46/i199  (.A1(\i43/i46/n72 ),
    .A2(\i43/i46/n70 ),
    .B1(\i43/i46/n42 ),
    .B2(\i43/i46/n63 ),
    .C(\i43/i46/n118 ),
    .Y(\i43/i46/n315 ));
 NOR2x1_ASAP7_75t_SL \i43/i46/i2  (.A(\i43/i46/n515 ),
    .B(\i43/i46/n511 ),
    .Y(\i43/n0 [30]));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i20  (.A(\i43/i46/n461 ),
    .B(\i43/i46/n468 ),
    .Y(\i43/i46/n501 ));
 OA211x2_ASAP7_75t_SL \i43/i46/i200  (.A1(\i43/i46/n37 ),
    .A2(\i43/i46/n137 ),
    .B(\i43/i46/n100 ),
    .C(\i43/i46/n160 ),
    .Y(\i43/i46/n314 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i46/i201  (.A1(\i43/i46/n47 ),
    .A2(\i43/i46/n34 ),
    .B(\i43/i46/n85 ),
    .C(\i43/i46/n242 ),
    .Y(\i43/i46/n313 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i202  (.A(\i43/i46/n267 ),
    .B(\i43/i46/n268 ),
    .Y(\i43/i46/n312 ));
 OAI31xp33_ASAP7_75t_SL \i43/i46/i203  (.A1(\i43/i46/n57 ),
    .A2(\i43/i46/n53 ),
    .A3(\i43/i46/n88 ),
    .B(\i43/i46/n62 ),
    .Y(\i43/i46/n311 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i204  (.A1(\i43/i46/n51 ),
    .A2(\i43/i46/n167 ),
    .B(\i43/i46/n71 ),
    .Y(\i43/i46/n310 ));
 OAI211xp5_ASAP7_75t_SL \i43/i46/i205  (.A1(\i43/i46/n52 ),
    .A2(\i43/i46/n91 ),
    .B(\i43/i46/n139 ),
    .C(\i43/i46/n140 ),
    .Y(\i43/i46/n309 ));
 OAI221xp5_ASAP7_75t_SL \i43/i46/i206  (.A1(\i43/i46/n94 ),
    .A2(\i43/i46/n87 ),
    .B1(\i43/i46/n78 ),
    .B2(\i43/i46/n54 ),
    .C(\i43/i46/n138 ),
    .Y(\i43/i46/n308 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i207  (.A1(\i43/i46/n56 ),
    .A2(\i43/i46/n157 ),
    .B1(\i43/i46/n63 ),
    .B2(\i43/i46/n72 ),
    .Y(\i43/i46/n307 ));
 OAI211xp5_ASAP7_75t_SL \i43/i46/i208  (.A1(\i43/i46/n82 ),
    .A2(\i43/i46/n72 ),
    .B(\i43/i46/n266 ),
    .C(\i43/i46/n179 ),
    .Y(\i43/i46/n306 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i46/i209  (.A1(\i43/i46/n51 ),
    .A2(\i43/i46/n53 ),
    .B(\i43/i46/n85 ),
    .C(\i43/i46/n204 ),
    .Y(\i43/i46/n305 ));
 NAND2x1_ASAP7_75t_SL \i43/i46/i21  (.A(\i43/i46/n467 ),
    .B(\i43/i46/n477 ),
    .Y(\i43/i46/n500 ));
 AOI221xp5_ASAP7_75t_SL \i43/i46/i210  (.A1(\i43/i46/n44 ),
    .A2(\i43/i46/n38 ),
    .B1(\i43/i46/n104 ),
    .B2(\i43/i46/n71 ),
    .C(\i43/i46/n162 ),
    .Y(\i43/i46/n304 ));
 NOR3xp33_ASAP7_75t_SL \i43/i46/i211  (.A(\i43/i46/n251 ),
    .B(\i43/i46/n171 ),
    .C(\i43/i46/n101 ),
    .Y(\i43/i46/n303 ));
 AOI21xp5_ASAP7_75t_SL \i43/i46/i212  (.A1(\i43/i46/n151 ),
    .A2(\i43/i46/n73 ),
    .B(\i43/i46/n263 ),
    .Y(\i43/i46/n302 ));
 OAI211xp5_ASAP7_75t_SL \i43/i46/i213  (.A1(\i43/i46/n89 ),
    .A2(\i43/i46/n158 ),
    .B(\i43/i46/n127 ),
    .C(\i43/i46/n136 ),
    .Y(\i43/i46/n301 ));
 AOI222xp33_ASAP7_75t_SL \i43/i46/i214  (.A1(\i43/i46/n67 ),
    .A2(\i43/i46/n112 ),
    .B1(\i43/i46/n65 ),
    .B2(\i43/i46/n79 ),
    .C1(\i43/i46/n59 ),
    .C2(\i43/i46/n48 ),
    .Y(\i43/i46/n300 ));
 NAND4xp25_ASAP7_75t_SL \i43/i46/i215  (.A(\i43/i46/n134 ),
    .B(\i43/i46/n165 ),
    .C(\i43/i46/n172 ),
    .D(\i43/i46/n111 ),
    .Y(\i43/i46/n299 ));
 AOI221xp5_ASAP7_75t_SL \i43/i46/i216  (.A1(\i43/i46/n48 ),
    .A2(\i43/i46/n81 ),
    .B1(\i43/i46/n41 ),
    .B2(\i43/i46/n85 ),
    .C(\i43/i46/n208 ),
    .Y(\i43/i46/n298 ));
 AOI222xp33_ASAP7_75t_SL \i43/i46/i217  (.A1(\i43/i46/n67 ),
    .A2(\i43/i46/n60 ),
    .B1(\i43/i46/n88 ),
    .B2(\i43/i46/n85 ),
    .C1(\i43/i46/n95 ),
    .C2(\i43/i46/n71 ),
    .Y(\i43/i46/n297 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i46/i218  (.A1(\i43/i46/n44 ),
    .A2(\i43/i46/n36 ),
    .B(\i43/i46/n48 ),
    .C(\i43/i46/n216 ),
    .Y(\i43/i46/n296 ));
 AOI22xp33_ASAP7_75t_SL \i43/i46/i219  (.A1(\i43/i46/n65 ),
    .A2(\i43/i46/n0 ),
    .B1(\i43/i46/n33 ),
    .B2(\i43/i46/n106 ),
    .Y(\i43/i46/n295 ));
 NAND4xp25_ASAP7_75t_SL \i43/i46/i22  (.A(\i43/i46/n430 ),
    .B(\i43/i46/n434 ),
    .C(\i43/i46/n393 ),
    .D(\i43/i46/n451 ),
    .Y(\i43/i46/n499 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i220  (.A1(\i43/i46/n75 ),
    .A2(\i43/i46/n103 ),
    .B1(\i43/i46/n46 ),
    .B2(\i43/i46/n37 ),
    .Y(\i43/i46/n294 ));
 AOI211xp5_ASAP7_75t_SL \i43/i46/i221  (.A1(\i43/i46/n67 ),
    .A2(\i43/i46/n79 ),
    .B(\i43/i46/n255 ),
    .C(\i43/i46/n171 ),
    .Y(\i43/i46/n293 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i222  (.A1(\i43/i46/n87 ),
    .A2(\i43/i46/n114 ),
    .B1(\i43/i46/n76 ),
    .B2(\i43/i46/n37 ),
    .Y(\i43/i46/n292 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i43/i46/i223  (.A1(\i43/i46/n42 ),
    .A2(\i43/i46/n49 ),
    .B(\i43/i46/n80 ),
    .C(\i43/i46/n253 ),
    .Y(\i43/i46/n291 ));
 AOI22xp5_ASAP7_75t_SL \i43/i46/i224  (.A1(\i43/i46/n83 ),
    .A2(\i43/i46/n144 ),
    .B1(\i43/i46/n71 ),
    .B2(\i43/i46/n38 ),
    .Y(\i43/i46/n290 ));
 AOI222xp33_ASAP7_75t_SL \i43/i46/i225  (.A1(\i43/i46/n79 ),
    .A2(\i43/i46/n48 ),
    .B1(\i43/i46/n69 ),
    .B2(\i43/i46/n38 ),
    .C1(\i43/i46/n74 ),
    .C2(\i43/i46/n67 ),
    .Y(\i43/i46/n289 ));
 OAI221xp5_ASAP7_75t_SL \i43/i46/i226  (.A1(\i43/i46/n35 ),
    .A2(\i43/i46/n80 ),
    .B1(\i43/i46/n68 ),
    .B2(\i43/i46/n76 ),
    .C(\i43/i46/n116 ),
    .Y(\i43/i46/n288 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i227  (.A(\i43/i46/n283 ),
    .B(\i43/i46/n284 ),
    .Y(\i43/i46/n287 ));
 AO21x1_ASAP7_75t_SL \i43/i46/i228  (.A1(\i43/i46/n41 ),
    .A2(\i43/i46/n164 ),
    .B(\i43/i46/n199 ),
    .Y(\i43/i46/n329 ));
 AOI21xp5_ASAP7_75t_SL \i43/i46/i229  (.A1(\i43/i46/n155 ),
    .A2(\i43/i46/n88 ),
    .B(\i43/i46/n203 ),
    .Y(\i43/i46/n328 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i23  (.A(\i43/i46/n478 ),
    .B(\i43/i46/n482 ),
    .Y(\i43/i46/n498 ));
 OA211x2_ASAP7_75t_SL \i43/i46/i230  (.A1(\i43/i46/n54 ),
    .A2(\i43/i46/n143 ),
    .B(\i43/i46/n129 ),
    .C(\i43/i46/n163 ),
    .Y(\i43/i46/n326 ));
 AOI22xp5_ASAP7_75t_SL \i43/i46/i231  (.A1(\i43/i46/n41 ),
    .A2(\i43/i46/n148 ),
    .B1(\i43/i46/n60 ),
    .B2(\i43/i46/n77 ),
    .Y(\i43/i46/n325 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i232  (.A(\i43/i46/n285 ),
    .B(\i43/i46/n239 ),
    .Y(\i43/i46/n286 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i233  (.A1(\i43/i46/n80 ),
    .A2(\i43/i46/n166 ),
    .B1(\i43/i46/n84 ),
    .B2(\i43/i46/n64 ),
    .Y(\i43/i46/n323 ));
 AOI21xp5_ASAP7_75t_SL \i43/i46/i234  (.A1(\i43/i46/n48 ),
    .A2(\i43/i46/n71 ),
    .B(\i43/i46/n219 ),
    .Y(\i43/i46/n322 ));
 AOI222xp33_ASAP7_75t_SL \i43/i46/i235  (.A1(\i43/i46/n43 ),
    .A2(\i43/i46/n59 ),
    .B1(\i43/i46/n73 ),
    .B2(\i43/i46/n85 ),
    .C1(\i43/i46/n34 ),
    .C2(\i43/i46/n71 ),
    .Y(\i43/i46/n321 ));
 O2A1O1Ixp5_ASAP7_75t_SL \i43/i46/i236  (.A1(\i43/i46/n41 ),
    .A2(\i43/i46/n48 ),
    .B(\i43/i46/n83 ),
    .C(\i43/i46/n225 ),
    .Y(\i43/i46/n320 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i237  (.A(\i43/i46/n108 ),
    .B(\i43/i46/n275 ),
    .Y(\i43/i46/n318 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i238  (.A(\i43/i46/n277 ),
    .Y(\i43/i46/n278 ));
 INVx1_ASAP7_75t_SL \i43/i46/i239  (.A(\i43/i46/n273 ),
    .Y(\i43/i46/n274 ));
 NOR2x1_ASAP7_75t_SL \i43/i46/i24  (.A(\i43/i46/n453 ),
    .B(\i43/i46/n474 ),
    .Y(\i43/i46/n507 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i240  (.A(\i43/i46/n270 ),
    .Y(\i43/i46/n271 ));
 OAI21xp33_ASAP7_75t_SL \i43/i46/i241  (.A1(\i43/i46/n75 ),
    .A2(\i43/i46/n52 ),
    .B(\i43/i46/n123 ),
    .Y(\i43/i46/n267 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i242  (.A(\i43/i46/n126 ),
    .B(\i43/i46/n153 ),
    .Y(\i43/i46/n266 ));
 NAND2xp33_ASAP7_75t_SL \i43/i46/i243  (.A(\i43/i46/n82 ),
    .B(\i43/i46/n128 ),
    .Y(\i43/i46/n265 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i244  (.A(\i43/i46/n75 ),
    .B(\i43/i46/n158 ),
    .Y(\i43/i46/n264 ));
 NAND2xp33_ASAP7_75t_SL \i43/i46/i245  (.A(\i43/i46/n185 ),
    .B(\i43/i46/n127 ),
    .Y(\i43/i46/n263 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i246  (.A(\i43/i46/n60 ),
    .B(\i43/i46/n148 ),
    .Y(\i43/i46/n262 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i247  (.A(\i43/i46/n55 ),
    .B(\i43/i46/n148 ),
    .Y(\i43/i46/n285 ));
 NOR3xp33_ASAP7_75t_SL \i43/i46/i248  (.A(\i43/i46/n71 ),
    .B(\i43/i46/n33 ),
    .C(\i43/i46/n81 ),
    .Y(\i43/i46/n261 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i249  (.A(\i43/i46/n125 ),
    .B(\i43/i46/n152 ),
    .Y(\i43/i46/n260 ));
 NOR3xp33_ASAP7_75t_SL \i43/i46/i25  (.A(\i43/i46/n455 ),
    .B(\i43/i46/n442 ),
    .C(\i43/i46/n398 ),
    .Y(\i43/i46/n506 ));
 NAND2xp33_ASAP7_75t_L \i43/i46/i250  (.A(\i43/i46/n150 ),
    .B(\i43/i46/n32 ),
    .Y(\i43/i46/n259 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i251  (.A1(\i43/i46/n79 ),
    .A2(\i43/i46/n33 ),
    .B(\i43/i46/n43 ),
    .Y(\i43/i46/n258 ));
 NAND2xp33_ASAP7_75t_SL \i43/i46/i252  (.A(\i43/i46/n42 ),
    .B(\i43/i46/n135 ),
    .Y(\i43/i46/n257 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i253  (.A1(\i43/i46/n87 ),
    .A2(\i43/i46/n64 ),
    .B(\i43/i46/n173 ),
    .Y(\i43/i46/n256 ));
 OAI21xp33_ASAP7_75t_SL \i43/i46/i254  (.A1(\i43/i46/n35 ),
    .A2(\i43/i46/n87 ),
    .B(\i43/i46/n160 ),
    .Y(\i43/i46/n255 ));
 OAI21xp33_ASAP7_75t_SL \i43/i46/i255  (.A1(\i43/i46/n84 ),
    .A2(\i43/i46/n42 ),
    .B(\i43/i46/n52 ),
    .Y(\i43/i46/n254 ));
 OAI21xp33_ASAP7_75t_SL \i43/i46/i256  (.A1(\i43/i46/n95 ),
    .A2(\i43/i46/n53 ),
    .B(\i43/i46/n164 ),
    .Y(\i43/i46/n253 ));
 OAI21xp33_ASAP7_75t_SL \i43/i46/i257  (.A1(\i43/i46/n66 ),
    .A2(\i43/i46/n80 ),
    .B(\i43/i46/n159 ),
    .Y(\i43/i46/n252 ));
 AOI21xp33_ASAP7_75t_SL \i43/i46/i258  (.A1(\i43/i46/n91 ),
    .A2(\i43/i46/n87 ),
    .B(\i43/i46/n49 ),
    .Y(\i43/i46/n251 ));
 OAI21xp33_ASAP7_75t_SL \i43/i46/i259  (.A1(\i43/i46/n58 ),
    .A2(\i43/i46/n35 ),
    .B(\i43/i46/n181 ),
    .Y(\i43/i46/n250 ));
 NAND3xp33_ASAP7_75t_SL \i43/i46/i26  (.A(\i43/i46/n447 ),
    .B(\i43/i46/n448 ),
    .C(\i43/i46/n446 ),
    .Y(\i43/i46/n497 ));
 OAI21xp33_ASAP7_75t_SL \i43/i46/i260  (.A1(\i43/i46/n82 ),
    .A2(\i43/i46/n35 ),
    .B(\i43/i46/n159 ),
    .Y(\i43/i46/n249 ));
 AOI21xp5_ASAP7_75t_SL \i43/i46/i261  (.A1(\i43/i46/n64 ),
    .A2(\i43/i46/n42 ),
    .B(\i43/i46/n91 ),
    .Y(\i43/i46/n284 ));
 AOI21xp5_ASAP7_75t_SL \i43/i46/i262  (.A1(\i43/i46/n83 ),
    .A2(\i43/i46/n65 ),
    .B(\i43/i46/n130 ),
    .Y(\i43/i46/n248 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i263  (.A1(\i43/i46/n74 ),
    .A2(\i43/i46/n86 ),
    .B(\i43/i46/n55 ),
    .Y(\i43/i46/n247 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i264  (.A1(\i43/i46/n77 ),
    .A2(\i43/i46/n34 ),
    .B(\i43/i46/n79 ),
    .Y(\i43/i46/n246 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i265  (.A1(\i43/i46/n66 ),
    .A2(\i43/i46/n84 ),
    .B(\i43/i46/n179 ),
    .Y(\i43/i46/n283 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i266  (.A1(\i43/i46/n81 ),
    .A2(\i43/i46/n62 ),
    .B(\i43/i46/n65 ),
    .Y(\i43/i46/n245 ));
 NAND3xp33_ASAP7_75t_L \i43/i46/i267  (.A(\i43/i46/n37 ),
    .B(\i43/i46/n87 ),
    .C(\i43/i46/n32 ),
    .Y(\i43/i46/n244 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i268  (.A1(\i43/i46/n90 ),
    .A2(\i43/i46/n69 ),
    .B(\i43/i46/n65 ),
    .Y(\i43/i46/n243 ));
 AOI21xp33_ASAP7_75t_SL \i43/i46/i269  (.A1(\i43/i46/n66 ),
    .A2(\i43/i46/n56 ),
    .B(\i43/i46/n75 ),
    .Y(\i43/i46/n242 ));
 NOR3x1_ASAP7_75t_SL \i43/i46/i27  (.A(\i43/i46/n457 ),
    .B(\i43/i46/n460 ),
    .C(\i43/i46/n442 ),
    .Y(\i43/i46/n496 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i270  (.A1(\i43/i46/n91 ),
    .A2(\i43/i46/n72 ),
    .B(\i43/i46/n186 ),
    .Y(\i43/i46/n241 ));
 OAI21xp33_ASAP7_75t_SL \i43/i46/i271  (.A1(\i43/i46/n80 ),
    .A2(\i43/i46/n54 ),
    .B(\i43/i46/n161 ),
    .Y(\i43/i46/n240 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i272  (.A1(\i43/i46/n39 ),
    .A2(\i43/i46/n82 ),
    .B(\i43/i46/n134 ),
    .Y(\i43/i46/n282 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i273  (.A1(\i43/i46/n92 ),
    .A2(\i43/i46/n72 ),
    .B(\i43/i46/n136 ),
    .Y(\i43/i46/n281 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i274  (.A1(\i43/i46/n54 ),
    .A2(\i43/i46/n58 ),
    .B1(\i43/i46/n50 ),
    .B2(\i43/i46/n92 ),
    .Y(\i43/i46/n280 ));
 AOI22xp5_ASAP7_75t_SL \i43/i46/i275  (.A1(\i43/i46/n55 ),
    .A2(\i43/i46/n44 ),
    .B1(\i43/i46/n85 ),
    .B2(\i43/i46/n48 ),
    .Y(\i43/i46/n279 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i276  (.A1(\i43/i46/n39 ),
    .A2(\i43/i46/n37 ),
    .B(\i43/i46/n172 ),
    .Y(\i43/i46/n277 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i277  (.A1(\i43/i46/n91 ),
    .A2(\i43/i46/n89 ),
    .B1(\i43/i46/n61 ),
    .B2(\i43/i46/n42 ),
    .Y(\i43/i46/n276 ));
 AOI22xp5_ASAP7_75t_SL \i43/i46/i278  (.A1(\i43/i46/n38 ),
    .A2(\i43/i46/n86 ),
    .B1(\i43/i46/n73 ),
    .B2(\i43/i46/n44 ),
    .Y(\i43/i46/n275 ));
 AOI22xp5_ASAP7_75t_SL \i43/i46/i279  (.A1(\i43/i46/n90 ),
    .A2(\i43/i46/n57 ),
    .B1(\i43/i46/n38 ),
    .B2(\i43/i46/n93 ),
    .Y(\i43/i46/n273 ));
 AND5x1_ASAP7_75t_SL \i43/i46/i28  (.A(\i43/i46/n454 ),
    .B(\i43/i46/n428 ),
    .C(\i43/i46/n378 ),
    .D(\i43/i46/n416 ),
    .E(\i43/i46/n418 ),
    .Y(\i43/i46/n495 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i280  (.A1(\i43/i46/n80 ),
    .A2(\i43/i46/n89 ),
    .B(\i43/i46/n168 ),
    .Y(\i43/i46/n272 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i281  (.A1(\i43/i46/n89 ),
    .A2(\i43/i46/n45 ),
    .B1(\i43/i46/n40 ),
    .B2(\i43/i46/n68 ),
    .Y(\i43/i46/n1 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i282  (.A(\i43/i46/n46 ),
    .B(\i43/i46/n170 ),
    .Y(\i43/i46/n270 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i283  (.A(\i43/i46/n85 ),
    .B(\i43/i46/n169 ),
    .Y(\i43/i46/n269 ));
 NOR2xp33_ASAP7_75t_L \i43/i46/i284  (.A(\i43/i46/n50 ),
    .B(\i43/i46/n154 ),
    .Y(\i43/i46/n268 ));
 INVx1_ASAP7_75t_SL \i43/i46/i285  (.A(\i43/i46/n235 ),
    .Y(\i43/i46/n236 ));
 INVxp33_ASAP7_75t_SL \i43/i46/i286  (.A(\i43/i46/n233 ),
    .Y(\i43/i46/n234 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i287  (.A(\i43/i46/n229 ),
    .Y(\i43/i46/n230 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i288  (.A(\i43/i46/n222 ),
    .Y(\i43/i46/n223 ));
 INVx1_ASAP7_75t_SL \i43/i46/i289  (.A(\i43/i46/n214 ),
    .Y(\i43/i46/n213 ));
 NOR3xp33_ASAP7_75t_SL \i43/i46/i29  (.A(\i43/i46/n471 ),
    .B(\i43/i46/n445 ),
    .C(\i43/i46/n431 ),
    .Y(\i43/i46/n494 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i290  (.A1(\i43/i46/n61 ),
    .A2(\i43/i46/n39 ),
    .B1(\i43/i46/n49 ),
    .B2(\i43/i46/n45 ),
    .Y(\i43/i46/n212 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i291  (.A1(\i43/i46/n53 ),
    .A2(\i43/i46/n34 ),
    .B(\i43/i46/n44 ),
    .Y(\i43/i46/n211 ));
 OAI22xp33_ASAP7_75t_SL \i43/i46/i292  (.A1(\i43/i46/n94 ),
    .A2(\i43/i46/n91 ),
    .B1(\i43/i46/n52 ),
    .B2(\i43/i46/n61 ),
    .Y(\i43/i46/n210 ));
 OAI21xp5_ASAP7_75t_SL \i43/i46/i293  (.A1(\i43/i46/n77 ),
    .A2(\i43/i46/n65 ),
    .B(\i43/i46/n36 ),
    .Y(\i43/i46/n209 ));
 AOI21xp33_ASAP7_75t_SL \i43/i46/i294  (.A1(\i43/i46/n66 ),
    .A2(\i43/i46/n72 ),
    .B(\i43/i46/n70 ),
    .Y(\i43/i46/n208 ));
 AOI21xp33_ASAP7_75t_SL \i43/i46/i295  (.A1(\i43/i46/n45 ),
    .A2(\i43/i46/n70 ),
    .B(\i43/i46/n52 ),
    .Y(\i43/i46/n207 ));
 AOI21xp5_ASAP7_75t_SL \i43/i46/i296  (.A1(\i43/i46/n57 ),
    .A2(\i43/i46/n60 ),
    .B(\i43/i46/n130 ),
    .Y(\i43/i46/n206 ));
 OAI22xp33_ASAP7_75t_SL \i43/i46/i297  (.A1(\i43/i46/n84 ),
    .A2(\i43/i46/n39 ),
    .B1(\i43/i46/n75 ),
    .B2(\i43/i46/n76 ),
    .Y(\i43/i46/n205 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i298  (.A1(\i43/i46/n75 ),
    .A2(\i43/i46/n54 ),
    .B1(\i43/i46/n40 ),
    .B2(\i43/i46/n61 ),
    .Y(\i43/i46/n204 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i299  (.A1(\i43/i46/n82 ),
    .A2(\i43/i46/n56 ),
    .B1(\i43/i46/n40 ),
    .B2(\i43/i46/n80 ),
    .Y(\i43/i46/n203 ));
 NOR2x1p5_ASAP7_75t_SL \i43/i46/i3  (.A(\i43/i46/n508 ),
    .B(\i43/i46/n513 ),
    .Y(\i43/n0 [28]));
 NOR3xp33_ASAP7_75t_SL \i43/i46/i30  (.A(\i43/i46/n456 ),
    .B(\i43/i46/n444 ),
    .C(\i43/i46/n435 ),
    .Y(\i43/i46/n493 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i300  (.A1(\i43/i46/n63 ),
    .A2(\i43/i46/n49 ),
    .B1(\i43/i46/n84 ),
    .B2(\i43/i46/n46 ),
    .Y(\i43/i46/n202 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i301  (.A1(\i43/i46/n50 ),
    .A2(\i43/i46/n91 ),
    .B1(\i43/i46/n39 ),
    .B2(\i43/i46/n63 ),
    .Y(\i43/i46/n201 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i302  (.A1(\i43/i46/n49 ),
    .A2(\i43/i46/n61 ),
    .B1(\i43/i46/n68 ),
    .B2(\i43/i46/n56 ),
    .Y(\i43/i46/n200 ));
 AOI22xp5_ASAP7_75t_SL \i43/i46/i303  (.A1(\i43/i46/n81 ),
    .A2(\i43/i46/n73 ),
    .B1(\i43/i46/n43 ),
    .B2(\i43/i46/n36 ),
    .Y(\i43/i46/n239 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i304  (.A1(\i43/i46/n82 ),
    .A2(\i43/i46/n89 ),
    .B1(\i43/i46/n75 ),
    .B2(\i43/i46/n46 ),
    .Y(\i43/i46/n199 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i305  (.A1(\i43/i46/n43 ),
    .A2(\i43/i46/n88 ),
    .B1(\i43/i46/n83 ),
    .B2(\i43/i46/n33 ),
    .Y(\i43/i46/n198 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i306  (.A1(\i43/i46/n80 ),
    .A2(\i43/i46/n64 ),
    .B1(\i43/i46/n68 ),
    .B2(\i43/i46/n35 ),
    .Y(\i43/i46/n197 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i307  (.A1(\i43/i46/n89 ),
    .A2(\i43/i46/n58 ),
    .B1(\i43/i46/n50 ),
    .B2(\i43/i46/n68 ),
    .Y(\i43/i46/n196 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i308  (.A1(\i43/i46/n32 ),
    .A2(\i43/i46/n89 ),
    .B1(\i43/i46/n52 ),
    .B2(\i43/i46/n58 ),
    .Y(\i43/i46/n195 ));
 AOI22xp5_ASAP7_75t_SL \i43/i46/i309  (.A1(\i43/i46/n53 ),
    .A2(\i43/i46/n79 ),
    .B1(\i43/i46/n95 ),
    .B2(\i43/i46/n44 ),
    .Y(\i43/i46/n238 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i31  (.A(\i43/i46/n452 ),
    .B(\i43/i46/n482 ),
    .Y(\i43/i46/n492 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i310  (.A1(\i43/i46/n70 ),
    .A2(\i43/i46/n64 ),
    .B1(\i43/i46/n72 ),
    .B2(\i43/i46/n37 ),
    .Y(\i43/i46/n237 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i311  (.A1(\i43/i46/n32 ),
    .A2(\i43/i46/n64 ),
    .B1(\i43/i46/n42 ),
    .B2(\i43/i46/n82 ),
    .Y(\i43/i46/n235 ));
 AOI22xp5_ASAP7_75t_SL \i43/i46/i312  (.A1(\i43/i46/n93 ),
    .A2(\i43/i46/n67 ),
    .B1(\i43/i46/n43 ),
    .B2(\i43/i46/n69 ),
    .Y(\i43/i46/n233 ));
 AO22x1_ASAP7_75t_SL \i43/i46/i313  (.A1(\i43/i46/n33 ),
    .A2(\i43/i46/n34 ),
    .B1(\i43/i46/n57 ),
    .B2(\i43/i46/n81 ),
    .Y(\i43/i46/n232 ));
 AOI22xp5_ASAP7_75t_SL \i43/i46/i314  (.A1(\i43/i46/n73 ),
    .A2(\i43/i46/n79 ),
    .B1(\i43/i46/n53 ),
    .B2(\i43/i46/n69 ),
    .Y(\i43/i46/n231 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i315  (.A1(\i43/i46/n58 ),
    .A2(\i43/i46/n64 ),
    .B1(\i43/i46/n54 ),
    .B2(\i43/i46/n63 ),
    .Y(\i43/i46/n229 ));
 AND2x2_ASAP7_75t_SL \i43/i46/i316  (.A(\i43/i46/n188 ),
    .B(\i43/i46/n189 ),
    .Y(\i43/i46/n194 ));
 NAND2xp33_ASAP7_75t_SL \i43/i46/i317  (.A(\i43/i46/n187 ),
    .B(\i43/i46/n177 ),
    .Y(\i43/i46/n193 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i318  (.A1(\i43/i46/n92 ),
    .A2(\i43/i46/n40 ),
    .B1(\i43/i46/n76 ),
    .B2(\i43/i46/n70 ),
    .Y(\i43/i46/n228 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i319  (.A1(\i43/i46/n35 ),
    .A2(\i43/i46/n63 ),
    .B1(\i43/i46/n72 ),
    .B2(\i43/i46/n68 ),
    .Y(\i43/i46/n227 ));
 NOR5xp2_ASAP7_75t_SL \i43/i46/i32  (.A(\i43/i46/n405 ),
    .B(\i43/i46/n414 ),
    .C(\i43/i46/n307 ),
    .D(\i43/i46/n402 ),
    .E(\i43/i46/n406 ),
    .Y(\i43/i46/n491 ));
 OAI22xp33_ASAP7_75t_SL \i43/i46/i320  (.A1(\i43/i46/n92 ),
    .A2(\i43/i46/n89 ),
    .B1(\i43/i46/n37 ),
    .B2(\i43/i46/n49 ),
    .Y(\i43/i46/n226 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i321  (.A1(\i43/i46/n92 ),
    .A2(\i43/i46/n49 ),
    .B1(\i43/i46/n42 ),
    .B2(\i43/i46/n75 ),
    .Y(\i43/i46/n225 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i322  (.A1(\i43/i46/n35 ),
    .A2(\i43/i46/n75 ),
    .B1(\i43/i46/n46 ),
    .B2(\i43/i46/n45 ),
    .Y(\i43/i46/n224 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i323  (.A1(\i43/i46/n80 ),
    .A2(\i43/i46/n39 ),
    .B1(\i43/i46/n54 ),
    .B2(\i43/i46/n68 ),
    .Y(\i43/i46/n222 ));
 AOI22xp5_ASAP7_75t_SL \i43/i46/i324  (.A1(\i43/i46/n33 ),
    .A2(\i43/i46/n57 ),
    .B1(\i43/i46/n41 ),
    .B2(\i43/i46/n36 ),
    .Y(\i43/i46/n221 ));
 OAI22xp33_ASAP7_75t_SL \i43/i46/i325  (.A1(\i43/i46/n87 ),
    .A2(\i43/i46/n89 ),
    .B1(\i43/i46/n78 ),
    .B2(\i43/i46/n42 ),
    .Y(\i43/i46/n220 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i326  (.A1(\i43/i46/n46 ),
    .A2(\i43/i46/n58 ),
    .B1(\i43/i46/n91 ),
    .B2(\i43/i46/n76 ),
    .Y(\i43/i46/n219 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i327  (.A1(\i43/i46/n68 ),
    .A2(\i43/i46/n64 ),
    .B1(\i43/i46/n50 ),
    .B2(\i43/i46/n37 ),
    .Y(\i43/i46/n218 ));
 AOI22xp5_ASAP7_75t_SL \i43/i46/i328  (.A1(\i43/i46/n79 ),
    .A2(\i43/i46/n57 ),
    .B1(\i43/i46/n95 ),
    .B2(\i43/i46/n69 ),
    .Y(\i43/i46/n217 ));
 OAI22xp5_ASAP7_75t_SL \i43/i46/i329  (.A1(\i43/i46/n78 ),
    .A2(\i43/i46/n89 ),
    .B1(\i43/i46/n50 ),
    .B2(\i43/i46/n32 ),
    .Y(\i43/i46/n216 ));
 NAND5xp2_ASAP7_75t_SL \i43/i46/i33  (.A(\i43/i46/n395 ),
    .B(\i43/i46/n424 ),
    .C(\i43/i46/n355 ),
    .D(\i43/i46/n320 ),
    .E(\i43/i46/n352 ),
    .Y(\i43/i46/n490 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i330  (.A(\i43/i46/n140 ),
    .B(\i43/i46/n139 ),
    .Y(\i43/i46/n192 ));
 AOI22xp5_ASAP7_75t_SL \i43/i46/i331  (.A1(\i43/i46/n93 ),
    .A2(\i43/i46/n34 ),
    .B1(\i43/i46/n77 ),
    .B2(\i43/i46/n62 ),
    .Y(\i43/i46/n215 ));
 OA22x2_ASAP7_75t_SL \i43/i46/i332  (.A1(\i43/i46/n61 ),
    .A2(\i43/i46/n64 ),
    .B1(\i43/i46/n58 ),
    .B2(\i43/i46/n76 ),
    .Y(\i43/i46/n214 ));
 INVx1_ASAP7_75t_SL \i43/i46/i333  (.A(\i43/i46/n190 ),
    .Y(\i43/i46/n191 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i334  (.A(\i43/i46/n183 ),
    .Y(\i43/i46/n184 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i335  (.A(\i43/i46/n177 ),
    .Y(\i43/i46/n178 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i336  (.A(\i43/i46/n175 ),
    .Y(\i43/i46/n176 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i337  (.A(\i43/i46/n169 ),
    .Y(\i43/i46/n170 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i338  (.A(\i43/i46/n166 ),
    .Y(\i43/i46/n167 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i339  (.A(\i43/i46/n161 ),
    .Y(\i43/i46/n162 ));
 NOR2x1_ASAP7_75t_SL \i43/i46/i34  (.A(\i43/i46/n464 ),
    .B(\i43/i46/n487 ),
    .Y(\i43/i46/n489 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i340  (.A(\i43/i46/n156 ),
    .Y(\i43/i46/n157 ));
 INVx1_ASAP7_75t_SL \i43/i46/i341  (.A(\i43/i46/n154 ),
    .Y(\i43/i46/n155 ));
 INVx1_ASAP7_75t_SL \i43/i46/i342  (.A(\i43/i46/n152 ),
    .Y(\i43/i46/n153 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i343  (.A(\i43/i46/n150 ),
    .Y(\i43/i46/n151 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i344  (.A(\i43/i46/n148 ),
    .Y(\i43/i46/n149 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i345  (.A(\i43/i46/n85 ),
    .B(\i43/i46/n51 ),
    .Y(\i43/i46/n147 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i346  (.A(\i43/i46/n77 ),
    .B(\i43/i46/n81 ),
    .Y(\i43/i46/n190 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i347  (.A(\i43/i46/n41 ),
    .B(\i43/i46/n90 ),
    .Y(\i43/i46/n146 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i348  (.A(\i43/i46/n90 ),
    .B(\i43/i46/n48 ),
    .Y(\i43/i46/n145 ));
 NAND2xp33_ASAP7_75t_SL \i43/i46/i349  (.A(\i43/i46/n46 ),
    .B(\i43/i46/n64 ),
    .Y(\i43/i46/n144 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i35  (.A(\i43/i46/n423 ),
    .B(\i43/i46/n486 ),
    .Y(\i43/i46/n488 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i350  (.A(\i43/i46/n36 ),
    .B(\i43/i46/n65 ),
    .Y(\i43/i46/n189 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i351  (.A(\i43/i46/n95 ),
    .B(\i43/i46/n93 ),
    .Y(\i43/i46/n188 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i352  (.A(\i43/i46/n67 ),
    .B(\i43/i46/n59 ),
    .Y(\i43/i46/n187 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i353  (.A(\i43/i46/n85 ),
    .B(\i43/i46/n71 ),
    .Y(\i43/i46/n143 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i354  (.A(\i43/i46/n58 ),
    .B(\i43/i46/n50 ),
    .Y(\i43/i46/n142 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i355  (.A(\i43/i46/n55 ),
    .B(\i43/i46/n83 ),
    .Y(\i43/i46/n186 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i356  (.A(\i43/i46/n69 ),
    .B(\i43/i46/n41 ),
    .Y(\i43/i46/n141 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i357  (.A(\i43/i46/n77 ),
    .B(\i43/i46/n93 ),
    .Y(\i43/i46/n185 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i358  (.A(\i43/i46/n75 ),
    .B(\i43/i46/n40 ),
    .Y(\i43/i46/n183 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i359  (.A(\i43/i46/n69 ),
    .B(\i43/i46/n67 ),
    .Y(\i43/i46/n182 ));
 INVx1_ASAP7_75t_SL \i43/i46/i36  (.A(\i43/i46/n483 ),
    .Y(\i43/i46/n484 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i360  (.A(\i43/i46/n79 ),
    .B(\i43/i46/n51 ),
    .Y(\i43/i46/n181 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i361  (.A(\i43/i46/n93 ),
    .B(\i43/i46/n65 ),
    .Y(\i43/i46/n180 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i362  (.A(\i43/i46/n79 ),
    .B(\i43/i46/n95 ),
    .Y(\i43/i46/n179 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i363  (.A(\i43/i46/n74 ),
    .B(\i43/i46/n65 ),
    .Y(\i43/i46/n177 ));
 AND2x2_ASAP7_75t_SL \i43/i46/i364  (.A(\i43/i46/n86 ),
    .B(\i43/i46/n77 ),
    .Y(\i43/i46/n175 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i365  (.A(\i43/i46/n85 ),
    .B(\i43/i46/n69 ),
    .Y(\i43/i46/n174 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i366  (.A(\i43/i46/n95 ),
    .B(\i43/i46/n36 ),
    .Y(\i43/i46/n173 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i367  (.A(\i43/i46/n44 ),
    .B(\i43/i46/n65 ),
    .Y(\i43/i46/n172 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i368  (.A(\i43/i46/n91 ),
    .B(\i43/i46/n46 ),
    .Y(\i43/i46/n171 ));
 NAND2xp5_ASAP7_75t_L \i43/i46/i369  (.A(\i43/i46/n35 ),
    .B(\i43/i46/n94 ),
    .Y(\i43/i46/n169 ));
 NAND2xp33_ASAP7_75t_L \i43/i46/i37  (.A(\i43/i46/n462 ),
    .B(\i43/i46/n429 ),
    .Y(\i43/i46/n481 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i370  (.A(\i43/i46/n95 ),
    .B(\i43/i46/n33 ),
    .Y(\i43/i46/n168 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i371  (.A(\i43/i46/n95 ),
    .B(\i43/i46/n43 ),
    .Y(\i43/i46/n166 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i372  (.A(\i43/i46/n57 ),
    .B(\i43/i46/n59 ),
    .Y(\i43/i46/n165 ));
 NAND2xp33_ASAP7_75t_SL \i43/i46/i373  (.A(\i43/i46/n61 ),
    .B(\i43/i46/n87 ),
    .Y(\i43/i46/n164 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i374  (.A(\i43/i46/n41 ),
    .B(\i43/i46/n59 ),
    .Y(\i43/i46/n163 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i375  (.A(\i43/i46/n73 ),
    .B(\i43/i46/n59 ),
    .Y(\i43/i46/n161 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i376  (.A(\i43/i46/n77 ),
    .B(\i43/i46/n83 ),
    .Y(\i43/i46/n160 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i377  (.A(\i43/i46/n85 ),
    .B(\i43/i46/n57 ),
    .Y(\i43/i46/n159 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i378  (.A(\i43/i46/n60 ),
    .B(\i43/i46/n69 ),
    .Y(\i43/i46/n158 ));
 NAND2xp5_ASAP7_75t_L \i43/i46/i379  (.A(\i43/i46/n37 ),
    .B(\i43/i46/n68 ),
    .Y(\i43/i46/n156 ));
 NAND2xp5_ASAP7_75t_L \i43/i46/i38  (.A(\i43/i46/n459 ),
    .B(\i43/i46/n411 ),
    .Y(\i43/i46/n480 ));
 NOR2x1_ASAP7_75t_SL \i43/i46/i380  (.A(\i43/i46/n62 ),
    .B(\i43/i46/n71 ),
    .Y(\i43/i46/n154 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i381  (.A(\i43/i46/n88 ),
    .B(\i43/i46/n36 ),
    .Y(\i43/i46/n152 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i382  (.A(\i43/i46/n86 ),
    .B(\i43/i46/n62 ),
    .Y(\i43/i46/n150 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i383  (.A(\i43/i46/n63 ),
    .B(\i43/i46/n84 ),
    .Y(\i43/i46/n0 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i384  (.A(\i43/i46/n32 ),
    .B(\i43/i46/n91 ),
    .Y(\i43/i46/n148 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i385  (.A(\i43/i46/n131 ),
    .Y(\i43/i46/n132 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i386  (.A(\i43/i46/n124 ),
    .Y(\i43/i46/n125 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i387  (.A(\i43/i46/n121 ),
    .Y(\i43/i46/n122 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i388  (.A(\i43/i46/n118 ),
    .Y(\i43/i46/n119 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i389  (.A(\i43/i46/n55 ),
    .B(\i43/i46/n36 ),
    .Y(\i43/i46/n116 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i39  (.A(\i43/i46/n458 ),
    .B(\i43/i46/n439 ),
    .Y(\i43/i46/n479 ));
 NAND2xp33_ASAP7_75t_SL \i43/i46/i390  (.A(\i43/i46/n70 ),
    .B(\i43/i46/n61 ),
    .Y(\i43/i46/n115 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i391  (.A(\i43/i46/n48 ),
    .B(\i43/i46/n57 ),
    .Y(\i43/i46/n114 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i392  (.A(\i43/i46/n51 ),
    .B(\i43/i46/n83 ),
    .Y(\i43/i46/n113 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i393  (.A(\i43/i46/n57 ),
    .B(\i43/i46/n36 ),
    .Y(\i43/i46/n140 ));
 NAND2xp33_ASAP7_75t_SL \i43/i46/i394  (.A(\i43/i46/n82 ),
    .B(\i43/i46/n45 ),
    .Y(\i43/i46/n112 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i395  (.A(\i43/i46/n71 ),
    .B(\i43/i46/n55 ),
    .Y(\i43/i46/n111 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i396  (.A(\i43/i46/n33 ),
    .B(\i43/i46/n38 ),
    .Y(\i43/i46/n110 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i397  (.A(\i43/i46/n75 ),
    .B(\i43/i46/n82 ),
    .Y(\i43/i46/n109 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i398  (.A(\i43/i46/n93 ),
    .B(\i43/i46/n53 ),
    .Y(\i43/i46/n108 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i399  (.A(\i43/i46/n44 ),
    .B(\i43/i46/n43 ),
    .Y(\i43/i46/n139 ));
 AND5x1_ASAP7_75t_SL \i43/i46/i4  (.A(\i43/i46/n509 ),
    .B(\i43/i46/n506 ),
    .C(\i43/i46/n486 ),
    .D(\i43/i46/n507 ),
    .E(\i43/i46/n476 ),
    .Y(\i43/n0 [27]));
 NAND4xp25_ASAP7_75t_SL \i43/i46/i40  (.A(\i43/i46/n422 ),
    .B(\i43/i46/n310 ),
    .C(\i43/i46/n313 ),
    .D(\i43/i46/n346 ),
    .Y(\i43/i46/n478 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i400  (.A(\i43/i46/n60 ),
    .B(\i43/i46/n34 ),
    .Y(\i43/i46/n107 ));
 NAND2xp33_ASAP7_75t_SL \i43/i46/i401  (.A(\i43/i46/n39 ),
    .B(\i43/i46/n66 ),
    .Y(\i43/i46/n106 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i402  (.A(\i43/i46/n47 ),
    .B(\i43/i46/n33 ),
    .Y(\i43/i46/n105 ));
 NAND2xp5_ASAP7_75t_L \i43/i46/i403  (.A(\i43/i46/n42 ),
    .B(\i43/i46/n66 ),
    .Y(\i43/i46/n104 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i404  (.A(\i43/i46/n38 ),
    .B(\i43/i46/n73 ),
    .Y(\i43/i46/n103 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i405  (.A(\i43/i46/n73 ),
    .B(\i43/i46/n60 ),
    .Y(\i43/i46/n138 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i406  (.A(\i43/i46/n41 ),
    .B(\i43/i46/n73 ),
    .Y(\i43/i46/n137 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i407  (.A(\i43/i46/n74 ),
    .B(\i43/i46/n48 ),
    .Y(\i43/i46/n136 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i408  (.A(\i43/i46/n72 ),
    .B(\i43/i46/n45 ),
    .Y(\i43/i46/n102 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i409  (.A(\i43/i46/n67 ),
    .B(\i43/i46/n36 ),
    .Y(\i43/i46/n135 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i41  (.A(\i43/i46/n441 ),
    .B(\i43/i46/n450 ),
    .Y(\i43/i46/n487 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i410  (.A(\i43/i46/n47 ),
    .B(\i43/i46/n93 ),
    .Y(\i43/i46/n134 ));
 NOR2xp33_ASAP7_75t_L \i43/i46/i411  (.A(\i43/i46/n35 ),
    .B(\i43/i46/n37 ),
    .Y(\i43/i46/n133 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i412  (.A(\i43/i46/n42 ),
    .B(\i43/i46/n75 ),
    .Y(\i43/i46/n101 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i413  (.A(\i43/i46/n71 ),
    .B(\i43/i46/n34 ),
    .Y(\i43/i46/n100 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i414  (.A(\i43/i46/n51 ),
    .B(\i43/i46/n44 ),
    .Y(\i43/i46/n131 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i415  (.A(\i43/i46/n92 ),
    .B(\i43/i46/n42 ),
    .Y(\i43/i46/n130 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i416  (.A(\i43/i46/n47 ),
    .B(\i43/i46/n81 ),
    .Y(\i43/i46/n129 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i417  (.A(\i43/i46/n47 ),
    .B(\i43/i46/n60 ),
    .Y(\i43/i46/n128 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i418  (.A(\i43/i46/n74 ),
    .B(\i43/i46/n51 ),
    .Y(\i43/i46/n127 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i419  (.A(\i43/i46/n38 ),
    .B(\i43/i46/n93 ),
    .Y(\i43/i46/n99 ));
 AND4x1_ASAP7_75t_SL \i43/i46/i42  (.A(\i43/i46/n443 ),
    .B(\i43/i46/n422 ),
    .C(\i43/i46/n356 ),
    .D(\i43/i46/n194 ),
    .Y(\i43/i46/n477 ));
 NOR2xp67_ASAP7_75t_SL \i43/i46/i420  (.A(\i43/i46/n50 ),
    .B(\i43/i46/n80 ),
    .Y(\i43/i46/n126 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i421  (.A(\i43/i46/n50 ),
    .B(\i43/i46/n92 ),
    .Y(\i43/i46/n98 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i422  (.A(\i43/i46/n61 ),
    .B(\i43/i46/n42 ),
    .Y(\i43/i46/n97 ));
 AND2x2_ASAP7_75t_SL \i43/i46/i423  (.A(\i43/i46/n93 ),
    .B(\i43/i46/n57 ),
    .Y(\i43/i46/n124 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i424  (.A(\i43/i46/n55 ),
    .B(\i43/i46/n44 ),
    .Y(\i43/i46/n96 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i425  (.A(\i43/i46/n79 ),
    .B(\i43/i46/n38 ),
    .Y(\i43/i46/n123 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i426  (.A(\i43/i46/n49 ),
    .B(\i43/i46/n32 ),
    .Y(\i43/i46/n121 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i427  (.A(\i43/i46/n33 ),
    .B(\i43/i46/n53 ),
    .Y(\i43/i46/n120 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i428  (.A(\i43/i46/n83 ),
    .B(\i43/i46/n53 ),
    .Y(\i43/i46/n118 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i429  (.A(\i43/i46/n60 ),
    .B(\i43/i46/n51 ),
    .Y(\i43/i46/n117 ));
 AND4x1_ASAP7_75t_SL \i43/i46/i43  (.A(\i43/i46/n384 ),
    .B(\i43/i46/n319 ),
    .C(\i43/i46/n371 ),
    .D(\i43/i46/n190 ),
    .Y(\i43/i46/n486 ));
 INVx1_ASAP7_75t_SL \i43/i46/i430  (.A(\i43/i46/n95 ),
    .Y(\i43/i46/n94 ));
 INVx3_ASAP7_75t_SL \i43/i46/i431  (.A(\i43/i46/n93 ),
    .Y(\i43/i46/n92 ));
 INVx1_ASAP7_75t_SL \i43/i46/i432  (.A(\i43/i46/n91 ),
    .Y(\i43/i46/n90 ));
 INVx2_ASAP7_75t_SL \i43/i46/i433  (.A(\i43/i46/n89 ),
    .Y(\i43/i46/n88 ));
 INVx2_ASAP7_75t_SL \i43/i46/i434  (.A(\i43/i46/n87 ),
    .Y(\i43/i46/n86 ));
 INVx2_ASAP7_75t_SL \i43/i46/i435  (.A(\i43/i46/n85 ),
    .Y(\i43/i46/n84 ));
 INVx4_ASAP7_75t_SL \i43/i46/i436  (.A(\i43/i46/n83 ),
    .Y(\i43/i46/n82 ));
 INVx3_ASAP7_75t_SL \i43/i46/i437  (.A(\i43/i46/n81 ),
    .Y(\i43/i46/n80 ));
 INVx1_ASAP7_75t_SL \i43/i46/i438  (.A(\i43/i46/n79 ),
    .Y(\i43/i46/n78 ));
 INVx2_ASAP7_75t_SL \i43/i46/i439  (.A(\i43/i46/n77 ),
    .Y(\i43/i46/n76 ));
 NOR2x1_ASAP7_75t_SL \i43/i46/i44  (.A(\i43/i46/n308 ),
    .B(\i43/i46/n460 ),
    .Y(\i43/i46/n485 ));
 INVx3_ASAP7_75t_SL \i43/i46/i440  (.A(\i43/i46/n75 ),
    .Y(\i43/i46/n74 ));
 INVx2_ASAP7_75t_SL \i43/i46/i441  (.A(\i43/i46/n73 ),
    .Y(\i43/i46/n72 ));
 INVx3_ASAP7_75t_SL \i43/i46/i442  (.A(\i43/i46/n71 ),
    .Y(\i43/i46/n70 ));
 INVx2_ASAP7_75t_SL \i43/i46/i443  (.A(\i43/i46/n69 ),
    .Y(\i43/i46/n68 ));
 INVx2_ASAP7_75t_SL \i43/i46/i444  (.A(\i43/i46/n67 ),
    .Y(\i43/i46/n66 ));
 INVx2_ASAP7_75t_SL \i43/i46/i445  (.A(\i43/i46/n65 ),
    .Y(\i43/i46/n64 ));
 AND2x4_ASAP7_75t_SL \i43/i46/i446  (.A(\i43/i46/n25 ),
    .B(\i43/i46/n15 ),
    .Y(\i43/i46/n95 ));
 AND2x4_ASAP7_75t_SL \i43/i46/i447  (.A(\i43/i46/n5 ),
    .B(\i43/i46/n6 ),
    .Y(\i43/i46/n93 ));
 OR2x2_ASAP7_75t_SL \i43/i46/i448  (.A(\i43/i46/n27 ),
    .B(\i43/i46/n11 ),
    .Y(\i43/i46/n91 ));
 OR2x2_ASAP7_75t_SL \i43/i46/i449  (.A(\i43/i46/n28 ),
    .B(\i43/i46/n9 ),
    .Y(\i43/i46/n89 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i45  (.A(\i43/i46/n461 ),
    .B(\i43/i46/n440 ),
    .Y(\i43/i46/n483 ));
 OR2x6_ASAP7_75t_SL \i43/i46/i450  (.A(\i43/i46/n7 ),
    .B(\i43/i46/n11 ),
    .Y(\i43/i46/n87 ));
 AND2x4_ASAP7_75t_SL \i43/i46/i451  (.A(\i43/i46/n4 ),
    .B(\i43/i46/n19 ),
    .Y(\i43/i46/n85 ));
 AND2x4_ASAP7_75t_SL \i43/i46/i452  (.A(\i43/i46/n10 ),
    .B(\i43/i46/n22 ),
    .Y(\i43/i46/n83 ));
 AND2x2_ASAP7_75t_SL \i43/i46/i453  (.A(\i43/i46/n6 ),
    .B(\i43/i46/n19 ),
    .Y(\i43/i46/n81 ));
 AND2x4_ASAP7_75t_SL \i43/i46/i454  (.A(\i43/i46/n5 ),
    .B(\i43/i46/n26 ),
    .Y(\i43/i46/n79 ));
 AND2x2_ASAP7_75t_SL \i43/i46/i455  (.A(\i43/i46/n16 ),
    .B(\i43/i46/n15 ),
    .Y(\i43/i46/n77 ));
 OR2x4_ASAP7_75t_SL \i43/i46/i456  (.A(\i43/i46/n3 ),
    .B(\i43/i46/n31 ),
    .Y(\i43/i46/n75 ));
 AND2x4_ASAP7_75t_SL \i43/i46/i457  (.A(\i43/i46/n25 ),
    .B(\i43/i46/n12 ),
    .Y(\i43/i46/n73 ));
 AND2x2_ASAP7_75t_SL \i43/i46/i458  (.A(\i43/i46/n4 ),
    .B(\i43/i46/n10 ),
    .Y(\i43/i46/n71 ));
 AND2x2_ASAP7_75t_SL \i43/i46/i459  (.A(\i43/i46/n5 ),
    .B(\i43/i46/n4 ),
    .Y(\i43/i46/n69 ));
 NAND2x1_ASAP7_75t_SL \i43/i46/i46  (.A(\i43/i46/n433 ),
    .B(\i43/i46/n397 ),
    .Y(\i43/i46/n482 ));
 AND2x4_ASAP7_75t_SL \i43/i46/i460  (.A(\i43/i46/n16 ),
    .B(\i43/i46/n29 ),
    .Y(\i43/i46/n67 ));
 AND2x4_ASAP7_75t_SL \i43/i46/i461  (.A(\i43/i46/n8 ),
    .B(\i43/i46/n12 ),
    .Y(\i43/i46/n65 ));
 INVx3_ASAP7_75t_SL \i43/i46/i462  (.A(\i43/i46/n63 ),
    .Y(\i43/i46/n62 ));
 INVx3_ASAP7_75t_SL \i43/i46/i463  (.A(\i43/i46/n61 ),
    .Y(\i43/i46/n60 ));
 INVx2_ASAP7_75t_SL \i43/i46/i464  (.A(\i43/i46/n59 ),
    .Y(\i43/i46/n58 ));
 INVx1_ASAP7_75t_SL \i43/i46/i465  (.A(\i43/i46/n57 ),
    .Y(\i43/i46/n56 ));
 INVx3_ASAP7_75t_SL \i43/i46/i466  (.A(\i43/i46/n55 ),
    .Y(\i43/i46/n54 ));
 INVx2_ASAP7_75t_SL \i43/i46/i467  (.A(\i43/i46/n53 ),
    .Y(\i43/i46/n52 ));
 INVx3_ASAP7_75t_SL \i43/i46/i468  (.A(\i43/i46/n51 ),
    .Y(\i43/i46/n50 ));
 INVx3_ASAP7_75t_SL \i43/i46/i469  (.A(\i43/i46/n49 ),
    .Y(\i43/i46/n48 ));
 NAND2xp5_ASAP7_75t_L \i43/i46/i47  (.A(\i43/i46/n443 ),
    .B(\i43/i46/n426 ),
    .Y(\i43/i46/n473 ));
 INVx3_ASAP7_75t_SL \i43/i46/i470  (.A(\i43/i46/n47 ),
    .Y(\i43/i46/n46 ));
 INVx3_ASAP7_75t_SL \i43/i46/i471  (.A(\i43/i46/n45 ),
    .Y(\i43/i46/n44 ));
 INVx3_ASAP7_75t_SL \i43/i46/i472  (.A(\i43/i46/n43 ),
    .Y(\i43/i46/n42 ));
 INVx2_ASAP7_75t_SL \i43/i46/i473  (.A(\i43/i46/n41 ),
    .Y(\i43/i46/n40 ));
 INVx3_ASAP7_75t_SL \i43/i46/i474  (.A(\i43/i46/n39 ),
    .Y(\i43/i46/n38 ));
 INVx2_ASAP7_75t_SL \i43/i46/i475  (.A(\i43/i46/n37 ),
    .Y(\i43/i46/n36 ));
 INVx4_ASAP7_75t_SL \i43/i46/i476  (.A(\i43/i46/n35 ),
    .Y(\i43/i46/n34 ));
 INVx3_ASAP7_75t_SL \i43/i46/i477  (.A(\i43/i46/n33 ),
    .Y(\i43/i46/n32 ));
 NAND2x1p5_ASAP7_75t_SL \i43/i46/i478  (.A(\i43/i46/n22 ),
    .B(\i43/i46/n5 ),
    .Y(\i43/i46/n63 ));
 OR2x2_ASAP7_75t_SL \i43/i46/i479  (.A(\i43/i46/n27 ),
    .B(\i43/i46/n20 ),
    .Y(\i43/i46/n61 ));
 AND3x1_ASAP7_75t_SL \i43/i46/i48  (.A(\i43/i46/n427 ),
    .B(\i43/i46/n410 ),
    .C(\i43/i46/n396 ),
    .Y(\i43/i46/n472 ));
 AND2x4_ASAP7_75t_SL \i43/i46/i480  (.A(\i43/i46/n6 ),
    .B(\i43/i46/n30 ),
    .Y(\i43/i46/n59 ));
 AND2x4_ASAP7_75t_SL \i43/i46/i481  (.A(\i43/i46/n25 ),
    .B(\i43/i46/n18 ),
    .Y(\i43/i46/n57 ));
 AND2x2_ASAP7_75t_SL \i43/i46/i482  (.A(\i43/i46/n8 ),
    .B(\i43/i46/n18 ),
    .Y(\i43/i46/n55 ));
 AND2x4_ASAP7_75t_SL \i43/i46/i483  (.A(\i43/i46/n16 ),
    .B(\i43/i46/n12 ),
    .Y(\i43/i46/n53 ));
 AND2x4_ASAP7_75t_SL \i43/i46/i484  (.A(\i43/i46/n25 ),
    .B(\i43/i46/n29 ),
    .Y(\i43/i46/n51 ));
 OR2x2_ASAP7_75t_SL \i43/i46/i485  (.A(\i43/i46/n17 ),
    .B(\i43/i46/n24 ),
    .Y(\i43/i46/n49 ));
 AND2x4_ASAP7_75t_SL \i43/i46/i486  (.A(\i43/i46/n23 ),
    .B(\i43/i46/n15 ),
    .Y(\i43/i46/n47 ));
 OR2x2_ASAP7_75t_SL \i43/i46/i487  (.A(\i43/i46/n27 ),
    .B(\i43/i46/n31 ),
    .Y(\i43/i46/n45 ));
 AND2x4_ASAP7_75t_SL \i43/i46/i488  (.A(\i43/i46/n23 ),
    .B(\i43/i46/n29 ),
    .Y(\i43/i46/n43 ));
 AND2x4_ASAP7_75t_SL \i43/i46/i489  (.A(\i43/i46/n16 ),
    .B(\i43/i46/n18 ),
    .Y(\i43/i46/n41 ));
 NAND4xp25_ASAP7_75t_SL \i43/i46/i49  (.A(\i43/i46/n425 ),
    .B(\i43/i46/n388 ),
    .C(\i43/i46/n314 ),
    .D(\i43/i46/n311 ),
    .Y(\i43/i46/n471 ));
 OR2x2_ASAP7_75t_SL \i43/i46/i490  (.A(\i43/i46/n14 ),
    .B(\i43/i46/n9 ),
    .Y(\i43/i46/n39 ));
 OR2x6_ASAP7_75t_SL \i43/i46/i491  (.A(\i43/i46/n20 ),
    .B(\i43/i46/n21 ),
    .Y(\i43/i46/n37 ));
 OR2x6_ASAP7_75t_SL \i43/i46/i492  (.A(\i43/i46/n24 ),
    .B(\i43/i46/n13 ),
    .Y(\i43/i46/n35 ));
 AND2x4_ASAP7_75t_SL \i43/i46/i493  (.A(\i43/i46/n30 ),
    .B(\i43/i46/n22 ),
    .Y(\i43/i46/n33 ));
 INVx2_ASAP7_75t_SL \i43/i46/i494  (.A(\i43/i46/n31 ),
    .Y(\i43/i46/n30 ));
 INVx1_ASAP7_75t_SL \i43/i46/i495  (.A(\i43/i46/n28 ),
    .Y(\i43/i46/n29 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i496  (.A(\i43/i46/n27 ),
    .Y(\i43/i46/n26 ));
 INVx1_ASAP7_75t_SL \i43/i46/i497  (.A(\i43/i46/n24 ),
    .Y(\i43/i46/n23 ));
 INVx3_ASAP7_75t_SL \i43/i46/i498  (.A(\i43/i46/n21 ),
    .Y(\i43/i46/n22 ));
 INVx1_ASAP7_75t_SL \i43/i46/i499  (.A(\i43/i46/n20 ),
    .Y(\i43/i46/n19 ));
 NAND5xp2_ASAP7_75t_SL \i43/i46/i5  (.A(\i43/i46/n475 ),
    .B(\i43/i46/n485 ),
    .C(\i43/i46/n479 ),
    .D(\i43/i46/n469 ),
    .E(\i43/i46/n463 ),
    .Y(\i43/i46/n515 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i50  (.A(\i43/i46/n248 ),
    .B(\i43/i46/n517 ),
    .Y(\i43/i46/n470 ));
 INVx1_ASAP7_75t_SL \i43/i46/i500  (.A(\i43/i46/n17 ),
    .Y(\i43/i46/n18 ));
 OR2x2_ASAP7_75t_SL \i43/i46/i501  (.A(n66),
    .B(n34[21]),
    .Y(\i43/i46/n31 ));
 OR2x2_ASAP7_75t_SL \i43/i46/i502  (.A(n67),
    .B(n34[16]),
    .Y(\i43/i46/n28 ));
 OR2x2_ASAP7_75t_SL \i43/i46/i503  (.A(n64),
    .B(n34[23]),
    .Y(\i43/i46/n27 ));
 AND2x2_ASAP7_75t_SL \i43/i46/i504  (.A(n34[17]),
    .B(\i43/i46/n2 ),
    .Y(\i43/i46/n25 ));
 NAND2x1p5_ASAP7_75t_SL \i43/i46/i505  (.A(n34[18]),
    .B(n68),
    .Y(\i43/i46/n24 ));
 OR2x2_ASAP7_75t_SL \i43/i46/i506  (.A(n63),
    .B(n34[22]),
    .Y(\i43/i46/n21 ));
 OR2x2_ASAP7_75t_SL \i43/i46/i507  (.A(n65),
    .B(n34[20]),
    .Y(\i43/i46/n20 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i508  (.A(n34[16]),
    .B(n67),
    .Y(\i43/i46/n17 ));
 INVx1_ASAP7_75t_SL \i43/i46/i509  (.A(\i43/i46/n14 ),
    .Y(\i43/i46/n15 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i51  (.A(\i43/i46/n417 ),
    .B(\i43/i46/n449 ),
    .Y(\i43/i46/n469 ));
 INVx2_ASAP7_75t_SL \i43/i46/i510  (.A(\i43/i46/n12 ),
    .Y(\i43/i46/n13 ));
 INVx1_ASAP7_75t_SL \i43/i46/i511  (.A(\i43/i46/n11 ),
    .Y(\i43/i46/n10 ));
 INVx1_ASAP7_75t_SL \i43/i46/i512  (.A(\i43/i46/n9 ),
    .Y(\i43/i46/n8 ));
 INVx1_ASAP7_75t_SL \i43/i46/i513  (.A(\i43/i46/n6 ),
    .Y(\i43/i46/n7 ));
 INVx2_ASAP7_75t_SL \i43/i46/i514  (.A(\i43/i46/n3 ),
    .Y(\i43/i46/n4 ));
 AND2x2_ASAP7_75t_SL \i43/i46/i515  (.A(n34[18]),
    .B(n34[17]),
    .Y(\i43/i46/n16 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i516  (.A(n34[19]),
    .B(n34[16]),
    .Y(\i43/i46/n14 ));
 AND2x2_ASAP7_75t_SL \i43/i46/i517  (.A(n67),
    .B(n69),
    .Y(\i43/i46/n12 ));
 OR2x2_ASAP7_75t_SL \i43/i46/i518  (.A(n34[21]),
    .B(n34[20]),
    .Y(\i43/i46/n11 ));
 OR2x2_ASAP7_75t_SL \i43/i46/i519  (.A(n34[18]),
    .B(n34[17]),
    .Y(\i43/i46/n9 ));
 NOR3xp33_ASAP7_75t_SL \i43/i46/i52  (.A(\i43/i46/n387 ),
    .B(\i43/i46/n403 ),
    .C(\i43/i46/n306 ),
    .Y(\i43/i46/n468 ));
 AND2x2_ASAP7_75t_SL \i43/i46/i520  (.A(n63),
    .B(n64),
    .Y(\i43/i46/n6 ));
 AND2x2_ASAP7_75t_SL \i43/i46/i521  (.A(n34[21]),
    .B(n34[20]),
    .Y(\i43/i46/n5 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i522  (.A(n34[23]),
    .B(n34[22]),
    .Y(\i43/i46/n3 ));
 INVxp67_ASAP7_75t_SL \i43/i46/i523  (.A(n34[18]),
    .Y(\i43/i46/n2 ));
 AND3x1_ASAP7_75t_SL \i43/i46/i524  (.A(\i43/i46/n462 ),
    .B(\i43/i46/n441 ),
    .C(\i43/i46/n475 ),
    .Y(\i43/i46/n516 ));
 AND3x1_ASAP7_75t_SL \i43/i46/i525  (.A(\i43/i46/n328 ),
    .B(\i43/i46/n269 ),
    .C(\i43/i46/n331 ),
    .Y(\i43/i46/n517 ));
 OR3x1_ASAP7_75t_SL \i43/i46/i526  (.A(\i43/i46/n224 ),
    .B(\i43/i46/n133 ),
    .C(\i43/i46/n200 ),
    .Y(\i43/i46/n518 ));
 NAND3xp33_ASAP7_75t_SL \i43/i46/i527  (.A(\i43/i46/n231 ),
    .B(\i43/i46/n117 ),
    .C(\i43/i46/n107 ),
    .Y(\i43/i46/n519 ));
 AOI211xp5_ASAP7_75t_SL \i43/i46/i53  (.A1(\i43/i46/n382 ),
    .A2(\i43/i46/n4 ),
    .B(\i43/i46/n399 ),
    .C(\i43/i46/n401 ),
    .Y(\i43/i46/n467 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i54  (.A(\i43/i46/n432 ),
    .B(\i43/i46/n438 ),
    .Y(\i43/i46/n466 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i55  (.A(\i43/i46/n398 ),
    .B(\i43/i46/n442 ),
    .Y(\i43/i46/n465 ));
 NOR2xp33_ASAP7_75t_L \i43/i46/i56  (.A(\i43/i46/n417 ),
    .B(\i43/i46/n437 ),
    .Y(\i43/i46/n476 ));
 OA211x2_ASAP7_75t_SL \i43/i46/i57  (.A1(\i43/i46/n91 ),
    .A2(\i43/i46/n66 ),
    .B(\i43/i46/n396 ),
    .C(\i43/i46/n373 ),
    .Y(\i43/i46/n475 ));
 NAND3xp33_ASAP7_75t_SL \i43/i46/i58  (.A(\i43/i46/n356 ),
    .B(\i43/i46/n383 ),
    .C(\i43/i46/n322 ),
    .Y(\i43/i46/n474 ));
 INVx1_ASAP7_75t_SL \i43/i46/i59  (.A(\i43/i46/n458 ),
    .Y(\i43/i46/n459 ));
 AND4x1_ASAP7_75t_SL \i43/i46/i6  (.A(\i43/i46/n503 ),
    .B(\i43/i46/n507 ),
    .C(\i43/i46/n493 ),
    .D(\i43/i46/n466 ),
    .Y(\i43/n0 [24]));
 INVxp67_ASAP7_75t_SL \i43/i46/i60  (.A(\i43/i46/n517 ),
    .Y(\i43/i46/n457 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i61  (.A(\i43/i46/n413 ),
    .B(\i43/i46/n397 ),
    .Y(\i43/i46/n456 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i62  (.A(\i43/i46/n302 ),
    .B(\i43/i46/n413 ),
    .Y(\i43/i46/n455 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i63  (.A(\i43/i46/n395 ),
    .B(\i43/i46/n392 ),
    .Y(\i43/i46/n464 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i64  (.A(\i43/i46/n518 ),
    .B(\i43/i46/n386 ),
    .Y(\i43/i46/n454 ));
 NAND2xp5_ASAP7_75t_L \i43/i46/i65  (.A(\i43/i46/n393 ),
    .B(\i43/i46/n312 ),
    .Y(\i43/i46/n453 ));
 NOR3xp33_ASAP7_75t_SL \i43/i46/i66  (.A(\i43/i46/n419 ),
    .B(\i43/i46/n345 ),
    .C(\i43/i46/n347 ),
    .Y(\i43/i46/n463 ));
 NAND3xp33_ASAP7_75t_SL \i43/i46/i67  (.A(\i43/i46/n394 ),
    .B(\i43/i46/n343 ),
    .C(\i43/i46/n217 ),
    .Y(\i43/i46/n452 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i68  (.A(\i43/i46/n301 ),
    .B(\i43/i46/n377 ),
    .Y(\i43/i46/n451 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i69  (.A(\i43/i46/n390 ),
    .B(\i43/i46/n519 ),
    .Y(\i43/i46/n450 ));
 AND4x2_ASAP7_75t_SL \i43/i46/i7  (.A(\i43/i46/n494 ),
    .B(\i43/i46/n498 ),
    .C(\i43/i46/n506 ),
    .D(\i43/i46/n516 ),
    .Y(\i43/n0 [31]));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i70  (.A(\i43/i46/n356 ),
    .B(\i43/i46/n404 ),
    .Y(\i43/i46/n449 ));
 OA211x2_ASAP7_75t_SL \i43/i46/i71  (.A1(\i43/i46/n66 ),
    .A2(\i43/i46/n87 ),
    .B(\i43/i46/n368 ),
    .C(\i43/i46/n371 ),
    .Y(\i43/i46/n448 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i72  (.A(\i43/i46/n391 ),
    .B(\i43/i46/n408 ),
    .Y(\i43/i46/n447 ));
 AND3x1_ASAP7_75t_SL \i43/i46/i73  (.A(\i43/i46/n355 ),
    .B(\i43/i46/n366 ),
    .C(\i43/i46/n351 ),
    .Y(\i43/i46/n446 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i74  (.A(\i43/i46/n380 ),
    .B(\i43/i46/n367 ),
    .Y(\i43/i46/n462 ));
 NOR3xp33_ASAP7_75t_SL \i43/i46/i75  (.A(\i43/i46/n329 ),
    .B(\i43/i46/n364 ),
    .C(\i43/i46/n202 ),
    .Y(\i43/i46/n461 ));
 NAND2x1_ASAP7_75t_SL \i43/i46/i76  (.A(\i43/i46/n385 ),
    .B(\i43/i46/n325 ),
    .Y(\i43/i46/n460 ));
 NAND2xp33_ASAP7_75t_SL \i43/i46/i77  (.A(\i43/i46/n371 ),
    .B(\i43/i46/n394 ),
    .Y(\i43/i46/n445 ));
 NAND3xp33_ASAP7_75t_SL \i43/i46/i78  (.A(\i43/i46/n320 ),
    .B(\i43/i46/n358 ),
    .C(\i43/i46/n297 ),
    .Y(\i43/i46/n458 ));
 NAND2xp33_ASAP7_75t_SL \i43/i46/i79  (.A(\i43/i46/n373 ),
    .B(\i43/i46/n396 ),
    .Y(\i43/i46/n444 ));
 NAND4xp75_ASAP7_75t_SL \i43/i46/i8  (.A(\i43/i46/n495 ),
    .B(\i43/i46/n496 ),
    .C(\i43/i46/n484 ),
    .D(\i43/i46/n472 ),
    .Y(\i43/i46/n514 ));
 NOR2x1_ASAP7_75t_SL \i43/i46/i80  (.A(\i43/i46/n381 ),
    .B(\i43/i46/n421 ),
    .Y(\i43/i46/n440 ));
 NAND2xp33_ASAP7_75t_SL \i43/i46/i81  (.A(\i43/i46/n412 ),
    .B(\i43/i46/n420 ),
    .Y(\i43/i46/n439 ));
 NAND4xp25_ASAP7_75t_SL \i43/i46/i82  (.A(\i43/i46/n325 ),
    .B(\i43/i46/n328 ),
    .C(\i43/i46/n296 ),
    .D(\i43/i46/n363 ),
    .Y(\i43/i46/n438 ));
 NAND3xp33_ASAP7_75t_SL \i43/i46/i83  (.A(\i43/i46/n324 ),
    .B(\i43/i46/n293 ),
    .C(\i43/i46/n278 ),
    .Y(\i43/i46/n437 ));
 NAND2xp5_ASAP7_75t_SL \i43/i46/i84  (.A(\i43/i46/n319 ),
    .B(\i43/i46/n389 ),
    .Y(\i43/i46/n436 ));
 NAND5xp2_ASAP7_75t_SL \i43/i46/i85  (.A(\i43/i46/n358 ),
    .B(\i43/i46/n215 ),
    .C(\i43/i46/n341 ),
    .D(\i43/i46/n236 ),
    .E(\i43/i46/n230 ),
    .Y(\i43/i46/n435 ));
 AOI211xp5_ASAP7_75t_SL \i43/i46/i86  (.A1(\i43/i46/n244 ),
    .A2(\i43/i46/n47 ),
    .B(\i43/i46/n286 ),
    .C(\i43/i46/n277 ),
    .Y(\i43/i46/n434 ));
 NOR2x1_ASAP7_75t_SL \i43/i46/i87  (.A(\i43/i46/n379 ),
    .B(\i43/i46/n415 ),
    .Y(\i43/i46/n433 ));
 NAND5xp2_ASAP7_75t_SL \i43/i46/i88  (.A(\i43/i46/n321 ),
    .B(\i43/i46/n370 ),
    .C(\i43/i46/n231 ),
    .D(\i43/i46/n128 ),
    .E(\i43/i46/n110 ),
    .Y(\i43/i46/n432 ));
 NAND4xp25_ASAP7_75t_SL \i43/i46/i89  (.A(\i43/i46/n355 ),
    .B(\i43/i46/n369 ),
    .C(\i43/i46/n348 ),
    .D(\i43/i46/n287 ),
    .Y(\i43/i46/n431 ));
 NAND4xp75_ASAP7_75t_SL \i43/i46/i9  (.A(\i43/i46/n489 ),
    .B(\i43/i46/n505 ),
    .C(\i43/i46/n502 ),
    .D(\i43/i46/n465 ),
    .Y(\i43/i46/n513 ));
 NOR2xp33_ASAP7_75t_SL \i43/i46/i90  (.A(\i43/i46/n349 ),
    .B(\i43/i46/n376 ),
    .Y(\i43/i46/n430 ));
 NOR5xp2_ASAP7_75t_SL \i43/i46/i91  (.A(\i43/i46/n337 ),
    .B(\i43/i46/n340 ),
    .C(\i43/i46/n119 ),
    .D(\i43/i46/n153 ),
    .E(\i43/i46/n102 ),
    .Y(\i43/i46/n429 ));
 AOI221xp5_ASAP7_75t_SL \i43/i46/i92  (.A1(\i43/i46/n259 ),
    .A2(\i43/i46/n55 ),
    .B1(\i43/i46/n156 ),
    .B2(\i43/i46/n257 ),
    .C(\i43/i46/n212 ),
    .Y(\i43/i46/n428 ));
 NOR5xp2_ASAP7_75t_SL \i43/i46/i93  (.A(\i43/i46/n213 ),
    .B(\i43/i46/n272 ),
    .C(\i43/i46/n240 ),
    .D(\i43/i46/n219 ),
    .E(\i43/i46/n178 ),
    .Y(\i43/i46/n427 ));
 NOR5xp2_ASAP7_75t_SL \i43/i46/i94  (.A(\i43/i46/n316 ),
    .B(\i43/i46/n353 ),
    .C(\i43/i46/n342 ),
    .D(\i43/i46/n218 ),
    .E(\i43/i46/n224 ),
    .Y(\i43/i46/n426 ));
 AOI211xp5_ASAP7_75t_SL \i43/i46/i95  (.A1(\i43/i46/n0 ),
    .A2(\i43/i46/n38 ),
    .B(\i43/i46/n299 ),
    .C(\i43/i46/n291 ),
    .Y(\i43/i46/n425 ));
 NOR5xp2_ASAP7_75t_SL \i43/i46/i96  (.A(\i43/i46/n330 ),
    .B(\i43/i46/n276 ),
    .C(\i43/i46/n282 ),
    .D(\i43/i46/n124 ),
    .E(\i43/i46/n175 ),
    .Y(\i43/i46/n424 ));
 NOR2xp67_ASAP7_75t_SL \i43/i46/i97  (.A(\i43/i46/n407 ),
    .B(\i43/i46/n409 ),
    .Y(\i43/i46/n443 ));
 AO211x2_ASAP7_75t_SL \i43/i46/i98  (.A1(\i43/i46/n88 ),
    .A2(\i43/i46/n264 ),
    .B(\i43/i46/n235 ),
    .C(\i43/i46/n315 ),
    .Y(\i43/i46/n442 ));
 AOI21xp5_ASAP7_75t_SL \i43/i46/i99  (.A1(\i43/i46/n33 ),
    .A2(\i43/i46/n73 ),
    .B(\i43/i46/n518 ),
    .Y(\i43/i46/n441 ));
 INVx1_ASAP7_75t_SL \i43/i460  (.A(\i43/n0 [13]),
    .Y(\i43/n171 ));
 INVxp67_ASAP7_75t_SL \i43/i461  (.A(\i43/n0 [6]),
    .Y(\i43/n170 ));
 INVx1_ASAP7_75t_SL \i43/i462  (.A(\i43/n0 [5]),
    .Y(\i43/n169 ));
 INVx1_ASAP7_75t_SL \i43/i463  (.A(n36[27]),
    .Y(\i43/n168 ));
 INVxp67_ASAP7_75t_SL \i43/i464  (.A(n37[12]),
    .Y(\i43/n167 ));
 INVx1_ASAP7_75t_SL \i43/i465  (.A(n36[29]),
    .Y(\i43/n166 ));
 INVxp67_ASAP7_75t_SL \i43/i466  (.A(n37[2]),
    .Y(\i43/n68 ));
 INVxp67_ASAP7_75t_SL \i43/i467  (.A(n37[27]),
    .Y(\i43/n165 ));
 INVxp67_ASAP7_75t_SL \i43/i468  (.A(net116),
    .Y(\i43/n164 ));
 INVxp67_ASAP7_75t_SL \i43/i469  (.A(net35),
    .Y(\i43/n163 ));
 NOR2x1_ASAP7_75t_SL \i43/i47/i0  (.A(\i43/i47/n479 ),
    .B(\i43/i47/n506 ),
    .Y(\i43/n0 [17]));
 AND3x1_ASAP7_75t_SL \i43/i47/i1  (.A(\i43/i47/n502 ),
    .B(\i43/i47/n504 ),
    .C(\i43/i47/n483 ),
    .Y(\i43/n0 [21]));
 NOR4xp75_ASAP7_75t_SL \i43/i47/i10  (.A(\i43/i47/n492 ),
    .B(\i43/i47/n496 ),
    .C(\i43/i47/n474 ),
    .D(\i43/i47/n489 ),
    .Y(\i43/n0 [18]));
 INVx1_ASAP7_75t_SL \i43/i47/i100  (.A(\i43/i47/n409 ),
    .Y(\i43/i47/n410 ));
 INVx1_ASAP7_75t_SL \i43/i47/i101  (.A(\i43/i47/n407 ),
    .Y(\i43/i47/n408 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i102  (.A(\i43/i47/n356 ),
    .B(\i43/i47/n351 ),
    .Y(\i43/i47/n406 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i103  (.A(\i43/i47/n325 ),
    .B(\i43/i47/n321 ),
    .Y(\i43/i47/n405 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i104  (.A(\i43/i47/n369 ),
    .B(\i43/i47/n324 ),
    .Y(\i43/i47/n404 ));
 NAND3xp33_ASAP7_75t_L \i43/i47/i105  (.A(\i43/i47/n267 ),
    .B(\i43/i47/n273 ),
    .C(\i43/i47/n354 ),
    .Y(\i43/i47/n403 ));
 NAND2xp5_ASAP7_75t_L \i43/i47/i106  (.A(\i43/i47/n337 ),
    .B(\i43/i47/n213 ),
    .Y(\i43/i47/n402 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i107  (.A(\i43/i47/n357 ),
    .B(\i43/i47/n331 ),
    .Y(\i43/i47/n401 ));
 NAND5xp2_ASAP7_75t_SL \i43/i47/i108  (.A(\i43/i47/n296 ),
    .B(\i43/i47/n120 ),
    .C(\i43/i47/n181 ),
    .D(\i43/i47/n123 ),
    .E(\i43/i47/n117 ),
    .Y(\i43/i47/n400 ));
 NOR4xp25_ASAP7_75t_SL \i43/i47/i109  (.A(\i43/i47/n279 ),
    .B(\i43/i47/n196 ),
    .C(\i43/i47/n131 ),
    .D(\i43/i47/n225 ),
    .Y(\i43/i47/n399 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i11  (.A(\i43/i47/n509 ),
    .B(\i43/i47/n491 ),
    .Y(\i43/i47/n504 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i110  (.A(\i43/i47/n347 ),
    .B(\i43/i47/n359 ),
    .Y(\i43/i47/n398 ));
 NAND2xp33_ASAP7_75t_SL \i43/i47/i111  (.A(\i43/i47/n320 ),
    .B(\i43/i47/n303 ),
    .Y(\i43/i47/n397 ));
 AOI221xp5_ASAP7_75t_SL \i43/i47/i112  (.A1(\i43/i47/n109 ),
    .A2(\i43/i47/n95 ),
    .B1(\i43/i47/n115 ),
    .B2(\i43/i47/n47 ),
    .C(\i43/i47/n215 ),
    .Y(\i43/i47/n416 ));
 NAND5xp2_ASAP7_75t_SL \i43/i47/i113  (.A(\i43/i47/n277 ),
    .B(\i43/i47/n205 ),
    .C(\i43/i47/n210 ),
    .D(\i43/i47/n181 ),
    .E(\i43/i47/n122 ),
    .Y(\i43/i47/n396 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i114  (.A(\i43/i47/n293 ),
    .B(\i43/i47/n369 ),
    .Y(\i43/i47/n395 ));
 OAI221xp5_ASAP7_75t_SL \i43/i47/i115  (.A1(\i43/i47/n156 ),
    .A2(\i43/i47/n54 ),
    .B1(\i43/i47/n157 ),
    .B2(\i43/i47/n39 ),
    .C(\i43/i47/n336 ),
    .Y(\i43/i47/n394 ));
 NOR2xp33_ASAP7_75t_L \i43/i47/i116  (.A(\i43/i47/n290 ),
    .B(\i43/i47/n356 ),
    .Y(\i43/i47/n415 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i117  (.A(\i43/i47/n287 ),
    .B(\i43/i47/n319 ),
    .Y(\i43/i47/n414 ));
 NOR3xp33_ASAP7_75t_SL \i43/i47/i118  (.A(\i43/i47/n217 ),
    .B(\i43/i47/n226 ),
    .C(\i43/i47/n195 ),
    .Y(\i43/i47/n412 ));
 NAND3xp33_ASAP7_75t_SL \i43/i47/i119  (.A(\i43/i47/n332 ),
    .B(\i43/i47/n283 ),
    .C(\i43/i47/n238 ),
    .Y(\i43/i47/n411 ));
 NAND3xp33_ASAP7_75t_SL \i43/i47/i12  (.A(\i43/i47/n477 ),
    .B(\i43/i47/n482 ),
    .C(\i43/i47/n416 ),
    .Y(\i43/i47/n503 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i120  (.A(\i43/i47/n214 ),
    .B(\i43/i47/n298 ),
    .Y(\i43/i47/n409 ));
 NOR3xp33_ASAP7_75t_SL \i43/i47/i121  (.A(\i43/i47/n286 ),
    .B(\i43/i47/n231 ),
    .C(\i43/i47/n270 ),
    .Y(\i43/i47/n407 ));
 INVx1_ASAP7_75t_SL \i43/i47/i122  (.A(\i43/i47/n514 ),
    .Y(\i43/i47/n387 ));
 OAI21xp33_ASAP7_75t_SL \i43/i47/i123  (.A1(\i43/i47/n76 ),
    .A2(\i43/i47/n45 ),
    .B(\i43/i47/n367 ),
    .Y(\i43/i47/n386 ));
 NOR3xp33_ASAP7_75t_SL \i43/i47/i124  (.A(\i43/i47/n327 ),
    .B(\i43/i47/n191 ),
    .C(\i43/i47/n231 ),
    .Y(\i43/i47/n385 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i125  (.A1(\i43/i47/n87 ),
    .A2(\i43/i47/n50 ),
    .B(\i43/i47/n354 ),
    .Y(\i43/i47/n393 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i126  (.A1(\i43/i47/n41 ),
    .A2(\i43/i47/n268 ),
    .B(\i43/i47/n263 ),
    .Y(\i43/i47/n384 ));
 NAND4xp25_ASAP7_75t_SL \i43/i47/i127  (.A(\i43/i47/n244 ),
    .B(\i43/i47/n145 ),
    .C(\i43/i47/n96 ),
    .D(\i43/i47/n99 ),
    .Y(\i43/i47/n383 ));
 NAND5xp2_ASAP7_75t_SL \i43/i47/i128  (.A(\i43/i47/n208 ),
    .B(\i43/i47/n120 ),
    .C(\i43/i47/n164 ),
    .D(\i43/i47/n184 ),
    .E(\i43/i47/n140 ),
    .Y(\i43/i47/n382 ));
 AOI211xp5_ASAP7_75t_SL \i43/i47/i129  (.A1(\i43/i47/n41 ),
    .A2(\i43/i47/n62 ),
    .B(\i43/i47/n282 ),
    .C(\i43/i47/n281 ),
    .Y(\i43/i47/n381 ));
 NOR3xp33_ASAP7_75t_SL \i43/i47/i13  (.A(\i43/i47/n508 ),
    .B(\i43/i47/n478 ),
    .C(\i43/i47/n455 ),
    .Y(\i43/i47/n502 ));
 NOR3xp33_ASAP7_75t_SL \i43/i47/i130  (.A(\i43/i47/n292 ),
    .B(\i43/i47/n206 ),
    .C(\i43/i47/n221 ),
    .Y(\i43/i47/n380 ));
 NOR2xp33_ASAP7_75t_L \i43/i47/i131  (.A(\i43/i47/n334 ),
    .B(\i43/i47/n315 ),
    .Y(\i43/i47/n379 ));
 OAI221xp5_ASAP7_75t_SL \i43/i47/i132  (.A1(\i43/i47/n269 ),
    .A2(\i43/i47/n75 ),
    .B1(\i43/i47/n173 ),
    .B2(\i43/i47/n72 ),
    .C(\i43/i47/n89 ),
    .Y(\i43/i47/n378 ));
 NAND5xp2_ASAP7_75t_SL \i43/i47/i133  (.A(\i43/i47/n246 ),
    .B(\i43/i47/n175 ),
    .C(\i43/i47/n105 ),
    .D(\i43/i47/n113 ),
    .E(\i43/i47/n144 ),
    .Y(\i43/i47/n377 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i134  (.A1(\i43/i47/n45 ),
    .A2(\i43/i47/n40 ),
    .B(\i43/i47/n357 ),
    .Y(\i43/i47/n376 ));
 NOR4xp25_ASAP7_75t_SL \i43/i47/i135  (.A(\i43/i47/n333 ),
    .B(\i43/i47/n266 ),
    .C(\i43/i47/n97 ),
    .D(\i43/i47/n98 ),
    .Y(\i43/i47/n375 ));
 OAI211xp5_ASAP7_75t_SL \i43/i47/i136  (.A1(\i43/i47/n40 ),
    .A2(\i43/i47/n259 ),
    .B(\i43/i47/n179 ),
    .C(\i43/i47/n167 ),
    .Y(\i43/i47/n374 ));
 NAND5xp2_ASAP7_75t_SL \i43/i47/i137  (.A(\i43/i47/n257 ),
    .B(\i43/i47/n242 ),
    .C(\i43/i47/n118 ),
    .D(\i43/i47/n180 ),
    .E(\i43/i47/n185 ),
    .Y(\i43/i47/n373 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i138  (.A(\i43/i47/n330 ),
    .B(\i43/i47/n301 ),
    .Y(\i43/i47/n372 ));
 OAI221xp5_ASAP7_75t_SL \i43/i47/i139  (.A1(\i43/i47/n260 ),
    .A2(\i43/i47/n54 ),
    .B1(\i43/i47/n52 ),
    .B2(\i43/i47/n87 ),
    .C(\i43/i47/n222 ),
    .Y(\i43/i47/n371 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i14  (.A(\i43/i47/n493 ),
    .B(\i43/i47/n481 ),
    .Y(\i43/i47/n501 ));
 NOR3xp33_ASAP7_75t_SL \i43/i47/i140  (.A(\i43/i47/n307 ),
    .B(\i43/i47/n274 ),
    .C(\i43/i47/n272 ),
    .Y(\i43/i47/n392 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i141  (.A(\i43/i47/n240 ),
    .B(\i43/i47/n358 ),
    .Y(\i43/i47/n391 ));
 OA211x2_ASAP7_75t_SL \i43/i47/i142  (.A1(\i43/i47/n92 ),
    .A2(\i43/i47/n54 ),
    .B(\i43/i47/n366 ),
    .C(\i43/i47/n146 ),
    .Y(\i43/i47/n390 ));
 NOR2xp33_ASAP7_75t_L \i43/i47/i143  (.A(\i43/i47/n190 ),
    .B(\i43/i47/n316 ),
    .Y(\i43/i47/n389 ));
 NOR2xp33_ASAP7_75t_L \i43/i47/i144  (.A(\i43/i47/n200 ),
    .B(\i43/i47/n362 ),
    .Y(\i43/i47/n388 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i145  (.A(\i43/i47/n364 ),
    .Y(\i43/i47/n365 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i146  (.A(\i43/i47/n362 ),
    .Y(\i43/i47/n363 ));
 INVx1_ASAP7_75t_SL \i43/i47/i147  (.A(\i43/i47/n360 ),
    .Y(\i43/i47/n361 ));
 INVx1_ASAP7_75t_SL \i43/i47/i148  (.A(\i43/i47/n358 ),
    .Y(\i43/i47/n359 ));
 INVx1_ASAP7_75t_SL \i43/i47/i149  (.A(\i43/i47/n512 ),
    .Y(\i43/i47/n352 ));
 NAND3xp33_ASAP7_75t_SL \i43/i47/i15  (.A(\i43/i47/n466 ),
    .B(\i43/i47/n476 ),
    .C(\i43/i47/n454 ),
    .Y(\i43/i47/n500 ));
 NAND2xp33_ASAP7_75t_L \i43/i47/i150  (.A(\i43/i47/n214 ),
    .B(\i43/i47/n271 ),
    .Y(\i43/i47/n351 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i151  (.A(\i43/i47/n130 ),
    .B(\i43/i47/n220 ),
    .Y(\i43/i47/n350 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i152  (.A(\i43/i47/n192 ),
    .B(\i43/i47/n212 ),
    .Y(\i43/i47/n349 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i47/i153  (.A1(\i43/i47/n34 ),
    .A2(\i43/i47/n65 ),
    .B(\i43/i47/n33 ),
    .C(\i43/i47/n227 ),
    .Y(\i43/i47/n348 ));
 OAI31xp33_ASAP7_75t_SL \i43/i47/i154  (.A1(\i43/i47/n65 ),
    .A2(\i43/i47/n41 ),
    .A3(\i43/i47/n55 ),
    .B(\i43/i47/n79 ),
    .Y(\i43/i47/n347 ));
 NAND3xp33_ASAP7_75t_SL \i43/i47/i155  (.A(\i43/i47/n213 ),
    .B(\i43/i47/n183 ),
    .C(\i43/i47/n128 ),
    .Y(\i43/i47/n346 ));
 AOI21xp5_ASAP7_75t_SL \i43/i47/i156  (.A1(\i43/i47/n38 ),
    .A2(\i43/i47/n74 ),
    .B(\i43/i47/n1 ),
    .Y(\i43/i47/n345 ));
 AOI211xp5_ASAP7_75t_SL \i43/i47/i157  (.A1(\i43/i47/n57 ),
    .A2(\i43/i47/n71 ),
    .B(\i43/i47/n182 ),
    .C(\i43/i47/n121 ),
    .Y(\i43/i47/n370 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i158  (.A1(\i43/i47/n94 ),
    .A2(\i43/i47/n58 ),
    .B(\i43/i47/n216 ),
    .Y(\i43/i47/n344 ));
 OAI31xp33_ASAP7_75t_SL \i43/i47/i159  (.A1(\i43/i47/n47 ),
    .A2(\i43/i47/n95 ),
    .A3(\i43/i47/n51 ),
    .B(\i43/i47/n69 ),
    .Y(\i43/i47/n343 ));
 NOR2xp33_ASAP7_75t_L \i43/i47/i16  (.A(\i43/i47/n465 ),
    .B(\i43/i47/n461 ),
    .Y(\i43/i47/n497 ));
 AO21x1_ASAP7_75t_SL \i43/i47/i160  (.A1(\i43/i47/n67 ),
    .A2(\i43/i47/n150 ),
    .B(\i43/i47/n280 ),
    .Y(\i43/i47/n342 ));
 AO21x1_ASAP7_75t_SL \i43/i47/i161  (.A1(\i43/i47/n148 ),
    .A2(\i43/i47/n173 ),
    .B(\i43/i47/n76 ),
    .Y(\i43/i47/n341 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i43/i47/i162  (.A1(\i43/i47/n70 ),
    .A2(\i43/i47/n78 ),
    .B(\i43/i47/n52 ),
    .C(\i43/i47/n197 ),
    .Y(\i43/i47/n340 ));
 AOI21xp5_ASAP7_75t_SL \i43/i47/i163  (.A1(\i43/i47/n44 ),
    .A2(\i43/i47/n67 ),
    .B(\i43/i47/n219 ),
    .Y(\i43/i47/n339 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i43/i47/i164  (.A1(\i43/i47/n42 ),
    .A2(\i43/i47/n35 ),
    .B(\i43/i47/n87 ),
    .C(\i43/i47/n117 ),
    .Y(\i43/i47/n338 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i165  (.A(\i43/i47/n249 ),
    .B(\i43/i47/n236 ),
    .Y(\i43/i47/n337 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i47/i166  (.A1(\i43/i47/n77 ),
    .A2(\i43/i47/n51 ),
    .B(\i43/i47/n33 ),
    .C(\i43/i47/n132 ),
    .Y(\i43/i47/n336 ));
 NAND3xp33_ASAP7_75t_SL \i43/i47/i167  (.A(\i43/i47/n232 ),
    .B(\i43/i47/n172 ),
    .C(\i43/i47/n137 ),
    .Y(\i43/i47/n335 ));
 OAI221xp5_ASAP7_75t_SL \i43/i47/i168  (.A1(\i43/i47/n75 ),
    .A2(\i43/i47/n56 ),
    .B1(\i43/i47/n49 ),
    .B2(\i43/i47/n68 ),
    .C(\i43/i47/n134 ),
    .Y(\i43/i47/n334 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i169  (.A1(\i43/i47/n78 ),
    .A2(\i43/i47/n136 ),
    .B(\i43/i47/n237 ),
    .Y(\i43/i47/n333 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i17  (.A(\i43/i47/n468 ),
    .B(\i43/i47/n476 ),
    .Y(\i43/i47/n496 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i170  (.A(\i43/i47/n233 ),
    .B(\i43/i47/n209 ),
    .Y(\i43/i47/n332 ));
 AOI221xp5_ASAP7_75t_SL \i43/i47/i171  (.A1(\i43/i47/n34 ),
    .A2(\i43/i47/n79 ),
    .B1(\i43/i47/n67 ),
    .B2(\i43/i47/n83 ),
    .C(\i43/i47/n236 ),
    .Y(\i43/i47/n331 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i172  (.A1(\i43/i47/n59 ),
    .A2(\i43/i47/n154 ),
    .B(\i43/i47/n77 ),
    .Y(\i43/i47/n330 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i47/i173  (.A1(\i43/i47/n62 ),
    .A2(\i43/i47/n44 ),
    .B(\i43/i47/n57 ),
    .C(\i43/i47/n125 ),
    .Y(\i43/i47/n329 ));
 OAI221xp5_ASAP7_75t_SL \i43/i47/i174  (.A1(\i43/i47/n46 ),
    .A2(\i43/i47/n87 ),
    .B1(\i43/i47/n52 ),
    .B2(\i43/i47/n80 ),
    .C(\i43/i47/n162 ),
    .Y(\i43/i47/n328 ));
 AOI21xp5_ASAP7_75t_SL \i43/i47/i175  (.A1(\i43/i47/n95 ),
    .A2(\i43/i47/n62 ),
    .B(\i43/i47/n1 ),
    .Y(\i43/i47/n369 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i176  (.A(\i43/i47/n219 ),
    .B(\i43/i47/n251 ),
    .Y(\i43/i47/n368 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i177  (.A(\i43/i47/n253 ),
    .B(\i43/i47/n0 ),
    .Y(\i43/i47/n367 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i178  (.A(\i43/i47/n225 ),
    .B(\i43/i47/n194 ),
    .Y(\i43/i47/n366 ));
 OAI211xp5_ASAP7_75t_SL \i43/i47/i179  (.A1(\i43/i47/n63 ),
    .A2(\i43/i47/n46 ),
    .B(\i43/i47/n176 ),
    .C(\i43/i47/n186 ),
    .Y(\i43/i47/n364 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i18  (.A(\i43/i47/n473 ),
    .B(\i43/i47/n464 ),
    .Y(\i43/i47/n495 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i180  (.A(\i43/i47/n120 ),
    .B(\i43/i47/n245 ),
    .Y(\i43/i47/n362 ));
 AOI222xp33_ASAP7_75t_SL \i43/i47/i181  (.A1(\i43/i47/n85 ),
    .A2(\i43/i47/n41 ),
    .B1(\i43/i47/n59 ),
    .B2(\i43/i47/n38 ),
    .C1(\i43/i47/n69 ),
    .C2(\i43/i47/n47 ),
    .Y(\i43/i47/n360 ));
 OAI221xp5_ASAP7_75t_SL \i43/i47/i182  (.A1(\i43/i47/n45 ),
    .A2(\i43/i47/n35 ),
    .B1(\i43/i47/n37 ),
    .B2(\i43/i47/n52 ),
    .C(\i43/i47/n179 ),
    .Y(\i43/i47/n358 ));
 AOI222xp33_ASAP7_75t_SL \i43/i47/i183  (.A1(\i43/i47/n34 ),
    .A2(\i43/i47/n90 ),
    .B1(\i43/i47/n33 ),
    .B2(\i43/i47/n67 ),
    .C1(\i43/i47/n83 ),
    .C2(\i43/i47/n73 ),
    .Y(\i43/i47/n357 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i184  (.A1(\i43/i47/n39 ),
    .A2(\i43/i47/n91 ),
    .B(\i43/i47/n237 ),
    .Y(\i43/i47/n356 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i185  (.A(\i43/i47/n204 ),
    .B(\i43/i47/n227 ),
    .Y(\i43/i47/n355 ));
 NOR2xp67_ASAP7_75t_SL \i43/i47/i186  (.A(\i43/i47/n255 ),
    .B(\i43/i47/n279 ),
    .Y(\i43/i47/n354 ));
 NOR2x1_ASAP7_75t_SL \i43/i47/i187  (.A(\i43/i47/n141 ),
    .B(\i43/i47/n278 ),
    .Y(\i43/i47/n353 ));
 INVxp33_ASAP7_75t_SL \i43/i47/i188  (.A(\i43/i47/n324 ),
    .Y(\i43/i47/n325 ));
 INVx1_ASAP7_75t_SL \i43/i47/i189  (.A(\i43/i47/n321 ),
    .Y(\i43/i47/n322 ));
 NOR4xp25_ASAP7_75t_SL \i43/i47/i19  (.A(\i43/i47/n429 ),
    .B(\i43/i47/n395 ),
    .C(\i43/i47/n372 ),
    .D(\i43/i47/n371 ),
    .Y(\i43/i47/n494 ));
 INVx1_ASAP7_75t_SL \i43/i47/i190  (.A(\i43/i47/n316 ),
    .Y(\i43/i47/n317 ));
 OAI211xp5_ASAP7_75t_SL \i43/i47/i191  (.A1(\i43/i47/n40 ),
    .A2(\i43/i47/n70 ),
    .B(\i43/i47/n188 ),
    .C(\i43/i47/n187 ),
    .Y(\i43/i47/n315 ));
 AO21x1_ASAP7_75t_SL \i43/i47/i192  (.A1(\i43/i47/n67 ),
    .A2(\i43/i47/n0 ),
    .B(\i43/i47/n224 ),
    .Y(\i43/i47/n314 ));
 OAI221xp5_ASAP7_75t_SL \i43/i47/i193  (.A1(\i43/i47/n72 ),
    .A2(\i43/i47/n70 ),
    .B1(\i43/i47/n42 ),
    .B2(\i43/i47/n63 ),
    .C(\i43/i47/n118 ),
    .Y(\i43/i47/n313 ));
 OA211x2_ASAP7_75t_SL \i43/i47/i194  (.A1(\i43/i47/n37 ),
    .A2(\i43/i47/n136 ),
    .B(\i43/i47/n100 ),
    .C(\i43/i47/n159 ),
    .Y(\i43/i47/n312 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i47/i195  (.A1(\i43/i47/n47 ),
    .A2(\i43/i47/n34 ),
    .B(\i43/i47/n85 ),
    .C(\i43/i47/n241 ),
    .Y(\i43/i47/n311 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i196  (.A(\i43/i47/n265 ),
    .B(\i43/i47/n266 ),
    .Y(\i43/i47/n310 ));
 OAI31xp33_ASAP7_75t_SL \i43/i47/i197  (.A1(\i43/i47/n57 ),
    .A2(\i43/i47/n53 ),
    .A3(\i43/i47/n88 ),
    .B(\i43/i47/n62 ),
    .Y(\i43/i47/n309 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i198  (.A1(\i43/i47/n51 ),
    .A2(\i43/i47/n166 ),
    .B(\i43/i47/n71 ),
    .Y(\i43/i47/n308 ));
 OAI211xp5_ASAP7_75t_SL \i43/i47/i199  (.A1(\i43/i47/n52 ),
    .A2(\i43/i47/n91 ),
    .B(\i43/i47/n138 ),
    .C(\i43/i47/n139 ),
    .Y(\i43/i47/n307 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i2  (.A(\i43/i47/n507 ),
    .B(\i43/i47/n503 ),
    .Y(\i43/n0 [22]));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i20  (.A(\i43/i47/n452 ),
    .B(\i43/i47/n459 ),
    .Y(\i43/i47/n493 ));
 OAI221xp5_ASAP7_75t_SL \i43/i47/i200  (.A1(\i43/i47/n94 ),
    .A2(\i43/i47/n87 ),
    .B1(\i43/i47/n78 ),
    .B2(\i43/i47/n54 ),
    .C(\i43/i47/n137 ),
    .Y(\i43/i47/n306 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i201  (.A1(\i43/i47/n56 ),
    .A2(\i43/i47/n156 ),
    .B1(\i43/i47/n63 ),
    .B2(\i43/i47/n72 ),
    .Y(\i43/i47/n305 ));
 OAI211xp5_ASAP7_75t_SL \i43/i47/i202  (.A1(\i43/i47/n82 ),
    .A2(\i43/i47/n72 ),
    .B(\i43/i47/n264 ),
    .C(\i43/i47/n178 ),
    .Y(\i43/i47/n304 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i47/i203  (.A1(\i43/i47/n51 ),
    .A2(\i43/i47/n53 ),
    .B(\i43/i47/n85 ),
    .C(\i43/i47/n203 ),
    .Y(\i43/i47/n303 ));
 AOI221xp5_ASAP7_75t_SL \i43/i47/i204  (.A1(\i43/i47/n44 ),
    .A2(\i43/i47/n38 ),
    .B1(\i43/i47/n104 ),
    .B2(\i43/i47/n71 ),
    .C(\i43/i47/n161 ),
    .Y(\i43/i47/n302 ));
 NOR3xp33_ASAP7_75t_SL \i43/i47/i205  (.A(\i43/i47/n250 ),
    .B(\i43/i47/n170 ),
    .C(\i43/i47/n101 ),
    .Y(\i43/i47/n301 ));
 AOI21xp5_ASAP7_75t_SL \i43/i47/i206  (.A1(\i43/i47/n150 ),
    .A2(\i43/i47/n73 ),
    .B(\i43/i47/n261 ),
    .Y(\i43/i47/n300 ));
 OAI211xp5_ASAP7_75t_SL \i43/i47/i207  (.A1(\i43/i47/n89 ),
    .A2(\i43/i47/n157 ),
    .B(\i43/i47/n126 ),
    .C(\i43/i47/n135 ),
    .Y(\i43/i47/n299 ));
 AOI222xp33_ASAP7_75t_SL \i43/i47/i208  (.A1(\i43/i47/n112 ),
    .A2(\i43/i47/n67 ),
    .B1(\i43/i47/n65 ),
    .B2(\i43/i47/n79 ),
    .C1(\i43/i47/n59 ),
    .C2(\i43/i47/n48 ),
    .Y(\i43/i47/n298 ));
 NAND4xp25_ASAP7_75t_SL \i43/i47/i209  (.A(\i43/i47/n133 ),
    .B(\i43/i47/n164 ),
    .C(\i43/i47/n171 ),
    .D(\i43/i47/n111 ),
    .Y(\i43/i47/n297 ));
 NAND2x1_ASAP7_75t_SL \i43/i47/i21  (.A(\i43/i47/n458 ),
    .B(\i43/i47/n469 ),
    .Y(\i43/i47/n492 ));
 AOI221xp5_ASAP7_75t_SL \i43/i47/i210  (.A1(\i43/i47/n48 ),
    .A2(\i43/i47/n81 ),
    .B1(\i43/i47/n41 ),
    .B2(\i43/i47/n85 ),
    .C(\i43/i47/n207 ),
    .Y(\i43/i47/n296 ));
 AOI222xp33_ASAP7_75t_SL \i43/i47/i211  (.A1(\i43/i47/n67 ),
    .A2(\i43/i47/n60 ),
    .B1(\i43/i47/n88 ),
    .B2(\i43/i47/n85 ),
    .C1(\i43/i47/n95 ),
    .C2(\i43/i47/n71 ),
    .Y(\i43/i47/n295 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i47/i212  (.A1(\i43/i47/n44 ),
    .A2(\i43/i47/n36 ),
    .B(\i43/i47/n48 ),
    .C(\i43/i47/n215 ),
    .Y(\i43/i47/n294 ));
 AOI22xp33_ASAP7_75t_SL \i43/i47/i213  (.A1(\i43/i47/n65 ),
    .A2(\i43/i47/n0 ),
    .B1(\i43/i47/n33 ),
    .B2(\i43/i47/n106 ),
    .Y(\i43/i47/n293 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i214  (.A1(\i43/i47/n75 ),
    .A2(\i43/i47/n103 ),
    .B1(\i43/i47/n46 ),
    .B2(\i43/i47/n37 ),
    .Y(\i43/i47/n292 ));
 AOI211xp5_ASAP7_75t_SL \i43/i47/i215  (.A1(\i43/i47/n67 ),
    .A2(\i43/i47/n79 ),
    .B(\i43/i47/n254 ),
    .C(\i43/i47/n170 ),
    .Y(\i43/i47/n291 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i216  (.A1(\i43/i47/n87 ),
    .A2(\i43/i47/n114 ),
    .B1(\i43/i47/n76 ),
    .B2(\i43/i47/n37 ),
    .Y(\i43/i47/n290 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i43/i47/i217  (.A1(\i43/i47/n42 ),
    .A2(\i43/i47/n49 ),
    .B(\i43/i47/n80 ),
    .C(\i43/i47/n252 ),
    .Y(\i43/i47/n289 ));
 AOI22xp5_ASAP7_75t_SL \i43/i47/i218  (.A1(\i43/i47/n83 ),
    .A2(\i43/i47/n143 ),
    .B1(\i43/i47/n71 ),
    .B2(\i43/i47/n38 ),
    .Y(\i43/i47/n288 ));
 AOI222xp33_ASAP7_75t_SL \i43/i47/i219  (.A1(\i43/i47/n79 ),
    .A2(\i43/i47/n48 ),
    .B1(\i43/i47/n69 ),
    .B2(\i43/i47/n38 ),
    .C1(\i43/i47/n74 ),
    .C2(\i43/i47/n67 ),
    .Y(\i43/i47/n287 ));
 NAND4xp25_ASAP7_75t_SL \i43/i47/i22  (.A(\i43/i47/n423 ),
    .B(\i43/i47/n427 ),
    .C(\i43/i47/n388 ),
    .D(\i43/i47/n443 ),
    .Y(\i43/i47/n491 ));
 OAI221xp5_ASAP7_75t_SL \i43/i47/i220  (.A1(\i43/i47/n35 ),
    .A2(\i43/i47/n80 ),
    .B1(\i43/i47/n68 ),
    .B2(\i43/i47/n76 ),
    .C(\i43/i47/n116 ),
    .Y(\i43/i47/n286 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i221  (.A(\i43/i47/n281 ),
    .B(\i43/i47/n282 ),
    .Y(\i43/i47/n285 ));
 AO21x1_ASAP7_75t_L \i43/i47/i222  (.A1(\i43/i47/n41 ),
    .A2(\i43/i47/n163 ),
    .B(\i43/i47/n198 ),
    .Y(\i43/i47/n327 ));
 AOI21xp5_ASAP7_75t_SL \i43/i47/i223  (.A1(\i43/i47/n154 ),
    .A2(\i43/i47/n88 ),
    .B(\i43/i47/n202 ),
    .Y(\i43/i47/n326 ));
 OA211x2_ASAP7_75t_SL \i43/i47/i224  (.A1(\i43/i47/n54 ),
    .A2(\i43/i47/n142 ),
    .B(\i43/i47/n128 ),
    .C(\i43/i47/n162 ),
    .Y(\i43/i47/n324 ));
 AOI22xp5_ASAP7_75t_SL \i43/i47/i225  (.A1(\i43/i47/n41 ),
    .A2(\i43/i47/n147 ),
    .B1(\i43/i47/n60 ),
    .B2(\i43/i47/n77 ),
    .Y(\i43/i47/n323 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i226  (.A(\i43/i47/n283 ),
    .B(\i43/i47/n238 ),
    .Y(\i43/i47/n284 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i227  (.A1(\i43/i47/n80 ),
    .A2(\i43/i47/n165 ),
    .B1(\i43/i47/n84 ),
    .B2(\i43/i47/n64 ),
    .Y(\i43/i47/n321 ));
 AOI21xp5_ASAP7_75t_SL \i43/i47/i228  (.A1(\i43/i47/n48 ),
    .A2(\i43/i47/n71 ),
    .B(\i43/i47/n218 ),
    .Y(\i43/i47/n320 ));
 AOI222xp33_ASAP7_75t_SL \i43/i47/i229  (.A1(\i43/i47/n43 ),
    .A2(\i43/i47/n59 ),
    .B1(\i43/i47/n73 ),
    .B2(\i43/i47/n85 ),
    .C1(\i43/i47/n34 ),
    .C2(\i43/i47/n71 ),
    .Y(\i43/i47/n319 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i23  (.A(\i43/i47/n470 ),
    .B(\i43/i47/n474 ),
    .Y(\i43/i47/n490 ));
 O2A1O1Ixp33_ASAP7_75t_L \i43/i47/i230  (.A1(\i43/i47/n41 ),
    .A2(\i43/i47/n48 ),
    .B(\i43/i47/n83 ),
    .C(\i43/i47/n224 ),
    .Y(\i43/i47/n318 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i231  (.A(\i43/i47/n108 ),
    .B(\i43/i47/n273 ),
    .Y(\i43/i47/n316 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i232  (.A(\i43/i47/n275 ),
    .Y(\i43/i47/n276 ));
 INVx1_ASAP7_75t_SL \i43/i47/i233  (.A(\i43/i47/n271 ),
    .Y(\i43/i47/n272 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i234  (.A(\i43/i47/n268 ),
    .Y(\i43/i47/n269 ));
 OAI21xp33_ASAP7_75t_SL \i43/i47/i235  (.A1(\i43/i47/n75 ),
    .A2(\i43/i47/n52 ),
    .B(\i43/i47/n123 ),
    .Y(\i43/i47/n265 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i236  (.A(\i43/i47/n125 ),
    .B(\i43/i47/n152 ),
    .Y(\i43/i47/n264 ));
 NAND2xp33_ASAP7_75t_SL \i43/i47/i237  (.A(\i43/i47/n82 ),
    .B(\i43/i47/n127 ),
    .Y(\i43/i47/n263 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i238  (.A(\i43/i47/n75 ),
    .B(\i43/i47/n157 ),
    .Y(\i43/i47/n262 ));
 NAND2xp33_ASAP7_75t_SL \i43/i47/i239  (.A(\i43/i47/n184 ),
    .B(\i43/i47/n126 ),
    .Y(\i43/i47/n261 ));
 NOR2x1_ASAP7_75t_SL \i43/i47/i24  (.A(\i43/i47/n445 ),
    .B(\i43/i47/n465 ),
    .Y(\i43/i47/n499 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i240  (.A(\i43/i47/n60 ),
    .B(\i43/i47/n147 ),
    .Y(\i43/i47/n260 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i241  (.A(\i43/i47/n55 ),
    .B(\i43/i47/n147 ),
    .Y(\i43/i47/n283 ));
 NOR3xp33_ASAP7_75t_SL \i43/i47/i242  (.A(\i43/i47/n71 ),
    .B(\i43/i47/n33 ),
    .C(\i43/i47/n81 ),
    .Y(\i43/i47/n259 ));
 NAND2xp33_ASAP7_75t_L \i43/i47/i243  (.A(\i43/i47/n149 ),
    .B(\i43/i47/n32 ),
    .Y(\i43/i47/n258 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i244  (.A1(\i43/i47/n79 ),
    .A2(\i43/i47/n33 ),
    .B(\i43/i47/n43 ),
    .Y(\i43/i47/n257 ));
 NAND2xp33_ASAP7_75t_SL \i43/i47/i245  (.A(\i43/i47/n42 ),
    .B(\i43/i47/n134 ),
    .Y(\i43/i47/n256 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i246  (.A1(\i43/i47/n87 ),
    .A2(\i43/i47/n64 ),
    .B(\i43/i47/n172 ),
    .Y(\i43/i47/n255 ));
 OAI21xp33_ASAP7_75t_SL \i43/i47/i247  (.A1(\i43/i47/n35 ),
    .A2(\i43/i47/n87 ),
    .B(\i43/i47/n159 ),
    .Y(\i43/i47/n254 ));
 OAI21xp33_ASAP7_75t_SL \i43/i47/i248  (.A1(\i43/i47/n84 ),
    .A2(\i43/i47/n42 ),
    .B(\i43/i47/n52 ),
    .Y(\i43/i47/n253 ));
 OAI21xp33_ASAP7_75t_SL \i43/i47/i249  (.A1(\i43/i47/n95 ),
    .A2(\i43/i47/n53 ),
    .B(\i43/i47/n163 ),
    .Y(\i43/i47/n252 ));
 NOR3xp33_ASAP7_75t_SL \i43/i47/i25  (.A(\i43/i47/n447 ),
    .B(\i43/i47/n434 ),
    .C(\i43/i47/n393 ),
    .Y(\i43/i47/n498 ));
 OAI21xp33_ASAP7_75t_SL \i43/i47/i250  (.A1(\i43/i47/n66 ),
    .A2(\i43/i47/n80 ),
    .B(\i43/i47/n158 ),
    .Y(\i43/i47/n251 ));
 AOI21xp33_ASAP7_75t_SL \i43/i47/i251  (.A1(\i43/i47/n91 ),
    .A2(\i43/i47/n87 ),
    .B(\i43/i47/n49 ),
    .Y(\i43/i47/n250 ));
 OAI21xp33_ASAP7_75t_SL \i43/i47/i252  (.A1(\i43/i47/n58 ),
    .A2(\i43/i47/n35 ),
    .B(\i43/i47/n180 ),
    .Y(\i43/i47/n249 ));
 OAI21xp33_ASAP7_75t_SL \i43/i47/i253  (.A1(\i43/i47/n82 ),
    .A2(\i43/i47/n35 ),
    .B(\i43/i47/n158 ),
    .Y(\i43/i47/n248 ));
 AOI21xp5_ASAP7_75t_SL \i43/i47/i254  (.A1(\i43/i47/n64 ),
    .A2(\i43/i47/n42 ),
    .B(\i43/i47/n91 ),
    .Y(\i43/i47/n282 ));
 AOI21xp5_ASAP7_75t_SL \i43/i47/i255  (.A1(\i43/i47/n83 ),
    .A2(\i43/i47/n65 ),
    .B(\i43/i47/n129 ),
    .Y(\i43/i47/n247 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i256  (.A1(\i43/i47/n74 ),
    .A2(\i43/i47/n86 ),
    .B(\i43/i47/n55 ),
    .Y(\i43/i47/n246 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i257  (.A1(\i43/i47/n77 ),
    .A2(\i43/i47/n34 ),
    .B(\i43/i47/n79 ),
    .Y(\i43/i47/n245 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i258  (.A1(\i43/i47/n66 ),
    .A2(\i43/i47/n84 ),
    .B(\i43/i47/n178 ),
    .Y(\i43/i47/n281 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i259  (.A1(\i43/i47/n81 ),
    .A2(\i43/i47/n62 ),
    .B(\i43/i47/n65 ),
    .Y(\i43/i47/n244 ));
 NAND3xp33_ASAP7_75t_SL \i43/i47/i26  (.A(\i43/i47/n438 ),
    .B(\i43/i47/n440 ),
    .C(\i43/i47/n439 ),
    .Y(\i43/i47/n489 ));
 NAND3xp33_ASAP7_75t_L \i43/i47/i260  (.A(\i43/i47/n37 ),
    .B(\i43/i47/n87 ),
    .C(\i43/i47/n32 ),
    .Y(\i43/i47/n243 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i261  (.A1(\i43/i47/n90 ),
    .A2(\i43/i47/n69 ),
    .B(\i43/i47/n65 ),
    .Y(\i43/i47/n242 ));
 AOI21xp33_ASAP7_75t_SL \i43/i47/i262  (.A1(\i43/i47/n66 ),
    .A2(\i43/i47/n56 ),
    .B(\i43/i47/n75 ),
    .Y(\i43/i47/n241 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i263  (.A1(\i43/i47/n91 ),
    .A2(\i43/i47/n72 ),
    .B(\i43/i47/n185 ),
    .Y(\i43/i47/n240 ));
 OAI21xp33_ASAP7_75t_SL \i43/i47/i264  (.A1(\i43/i47/n80 ),
    .A2(\i43/i47/n54 ),
    .B(\i43/i47/n160 ),
    .Y(\i43/i47/n239 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i265  (.A1(\i43/i47/n39 ),
    .A2(\i43/i47/n82 ),
    .B(\i43/i47/n133 ),
    .Y(\i43/i47/n280 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i266  (.A1(\i43/i47/n92 ),
    .A2(\i43/i47/n72 ),
    .B(\i43/i47/n135 ),
    .Y(\i43/i47/n279 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i267  (.A1(\i43/i47/n54 ),
    .A2(\i43/i47/n58 ),
    .B1(\i43/i47/n50 ),
    .B2(\i43/i47/n92 ),
    .Y(\i43/i47/n278 ));
 AOI22xp5_ASAP7_75t_SL \i43/i47/i268  (.A1(\i43/i47/n55 ),
    .A2(\i43/i47/n44 ),
    .B1(\i43/i47/n85 ),
    .B2(\i43/i47/n48 ),
    .Y(\i43/i47/n277 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i269  (.A1(\i43/i47/n39 ),
    .A2(\i43/i47/n37 ),
    .B(\i43/i47/n171 ),
    .Y(\i43/i47/n275 ));
 NOR3xp33_ASAP7_75t_SL \i43/i47/i27  (.A(\i43/i47/n449 ),
    .B(\i43/i47/n451 ),
    .C(\i43/i47/n434 ),
    .Y(\i43/i47/n488 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i270  (.A1(\i43/i47/n91 ),
    .A2(\i43/i47/n89 ),
    .B1(\i43/i47/n61 ),
    .B2(\i43/i47/n42 ),
    .Y(\i43/i47/n274 ));
 AOI22xp5_ASAP7_75t_SL \i43/i47/i271  (.A1(\i43/i47/n38 ),
    .A2(\i43/i47/n86 ),
    .B1(\i43/i47/n73 ),
    .B2(\i43/i47/n44 ),
    .Y(\i43/i47/n273 ));
 AOI22xp5_ASAP7_75t_SL \i43/i47/i272  (.A1(\i43/i47/n90 ),
    .A2(\i43/i47/n57 ),
    .B1(\i43/i47/n38 ),
    .B2(\i43/i47/n93 ),
    .Y(\i43/i47/n271 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i273  (.A1(\i43/i47/n80 ),
    .A2(\i43/i47/n89 ),
    .B(\i43/i47/n167 ),
    .Y(\i43/i47/n270 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i274  (.A1(\i43/i47/n89 ),
    .A2(\i43/i47/n45 ),
    .B1(\i43/i47/n40 ),
    .B2(\i43/i47/n68 ),
    .Y(\i43/i47/n1 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i275  (.A(\i43/i47/n46 ),
    .B(\i43/i47/n169 ),
    .Y(\i43/i47/n268 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i276  (.A(\i43/i47/n85 ),
    .B(\i43/i47/n168 ),
    .Y(\i43/i47/n267 ));
 NOR2xp33_ASAP7_75t_L \i43/i47/i277  (.A(\i43/i47/n50 ),
    .B(\i43/i47/n153 ),
    .Y(\i43/i47/n266 ));
 INVx1_ASAP7_75t_SL \i43/i47/i278  (.A(\i43/i47/n234 ),
    .Y(\i43/i47/n235 ));
 INVxp33_ASAP7_75t_SL \i43/i47/i279  (.A(\i43/i47/n232 ),
    .Y(\i43/i47/n233 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i28  (.A(\i43/i47/n472 ),
    .B(\i43/i47/n467 ),
    .Y(\i43/i47/n487 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i280  (.A(\i43/i47/n228 ),
    .Y(\i43/i47/n229 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i281  (.A(\i43/i47/n221 ),
    .Y(\i43/i47/n222 ));
 INVx1_ASAP7_75t_SL \i43/i47/i282  (.A(\i43/i47/n213 ),
    .Y(\i43/i47/n212 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i283  (.A1(\i43/i47/n61 ),
    .A2(\i43/i47/n39 ),
    .B1(\i43/i47/n49 ),
    .B2(\i43/i47/n45 ),
    .Y(\i43/i47/n211 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i284  (.A1(\i43/i47/n53 ),
    .A2(\i43/i47/n34 ),
    .B(\i43/i47/n44 ),
    .Y(\i43/i47/n210 ));
 OAI22xp33_ASAP7_75t_SL \i43/i47/i285  (.A1(\i43/i47/n94 ),
    .A2(\i43/i47/n91 ),
    .B1(\i43/i47/n52 ),
    .B2(\i43/i47/n61 ),
    .Y(\i43/i47/n209 ));
 OAI21xp5_ASAP7_75t_SL \i43/i47/i286  (.A1(\i43/i47/n77 ),
    .A2(\i43/i47/n65 ),
    .B(\i43/i47/n36 ),
    .Y(\i43/i47/n208 ));
 AOI21xp33_ASAP7_75t_SL \i43/i47/i287  (.A1(\i43/i47/n66 ),
    .A2(\i43/i47/n72 ),
    .B(\i43/i47/n70 ),
    .Y(\i43/i47/n207 ));
 AOI21xp33_ASAP7_75t_SL \i43/i47/i288  (.A1(\i43/i47/n45 ),
    .A2(\i43/i47/n70 ),
    .B(\i43/i47/n52 ),
    .Y(\i43/i47/n206 ));
 AOI21xp5_ASAP7_75t_SL \i43/i47/i289  (.A1(\i43/i47/n57 ),
    .A2(\i43/i47/n60 ),
    .B(\i43/i47/n129 ),
    .Y(\i43/i47/n205 ));
 AND5x1_ASAP7_75t_SL \i43/i47/i29  (.A(\i43/i47/n446 ),
    .B(\i43/i47/n421 ),
    .C(\i43/i47/n375 ),
    .D(\i43/i47/n410 ),
    .E(\i43/i47/n412 ),
    .Y(\i43/i47/n486 ));
 OAI22xp33_ASAP7_75t_SL \i43/i47/i290  (.A1(\i43/i47/n84 ),
    .A2(\i43/i47/n39 ),
    .B1(\i43/i47/n75 ),
    .B2(\i43/i47/n76 ),
    .Y(\i43/i47/n204 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i291  (.A1(\i43/i47/n75 ),
    .A2(\i43/i47/n54 ),
    .B1(\i43/i47/n40 ),
    .B2(\i43/i47/n61 ),
    .Y(\i43/i47/n203 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i292  (.A1(\i43/i47/n82 ),
    .A2(\i43/i47/n56 ),
    .B1(\i43/i47/n40 ),
    .B2(\i43/i47/n80 ),
    .Y(\i43/i47/n202 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i293  (.A1(\i43/i47/n63 ),
    .A2(\i43/i47/n49 ),
    .B1(\i43/i47/n84 ),
    .B2(\i43/i47/n46 ),
    .Y(\i43/i47/n201 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i294  (.A1(\i43/i47/n50 ),
    .A2(\i43/i47/n91 ),
    .B1(\i43/i47/n39 ),
    .B2(\i43/i47/n63 ),
    .Y(\i43/i47/n200 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i295  (.A1(\i43/i47/n49 ),
    .A2(\i43/i47/n61 ),
    .B1(\i43/i47/n68 ),
    .B2(\i43/i47/n56 ),
    .Y(\i43/i47/n199 ));
 AOI22xp5_ASAP7_75t_SL \i43/i47/i296  (.A1(\i43/i47/n81 ),
    .A2(\i43/i47/n73 ),
    .B1(\i43/i47/n43 ),
    .B2(\i43/i47/n36 ),
    .Y(\i43/i47/n238 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i297  (.A1(\i43/i47/n82 ),
    .A2(\i43/i47/n89 ),
    .B1(\i43/i47/n75 ),
    .B2(\i43/i47/n46 ),
    .Y(\i43/i47/n198 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i298  (.A1(\i43/i47/n43 ),
    .A2(\i43/i47/n88 ),
    .B1(\i43/i47/n83 ),
    .B2(\i43/i47/n33 ),
    .Y(\i43/i47/n197 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i299  (.A1(\i43/i47/n80 ),
    .A2(\i43/i47/n64 ),
    .B1(\i43/i47/n68 ),
    .B2(\i43/i47/n35 ),
    .Y(\i43/i47/n196 ));
 NOR2x1_ASAP7_75t_SL \i43/i47/i3  (.A(\i43/i47/n500 ),
    .B(\i43/i47/n505 ),
    .Y(\i43/n0 [20]));
 NOR3xp33_ASAP7_75t_SL \i43/i47/i30  (.A(\i43/i47/n462 ),
    .B(\i43/i47/n437 ),
    .C(\i43/i47/n424 ),
    .Y(\i43/i47/n485 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i300  (.A1(\i43/i47/n89 ),
    .A2(\i43/i47/n58 ),
    .B1(\i43/i47/n50 ),
    .B2(\i43/i47/n68 ),
    .Y(\i43/i47/n195 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i301  (.A1(\i43/i47/n32 ),
    .A2(\i43/i47/n89 ),
    .B1(\i43/i47/n52 ),
    .B2(\i43/i47/n58 ),
    .Y(\i43/i47/n194 ));
 AOI22xp5_ASAP7_75t_SL \i43/i47/i302  (.A1(\i43/i47/n53 ),
    .A2(\i43/i47/n79 ),
    .B1(\i43/i47/n95 ),
    .B2(\i43/i47/n44 ),
    .Y(\i43/i47/n237 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i303  (.A1(\i43/i47/n70 ),
    .A2(\i43/i47/n64 ),
    .B1(\i43/i47/n72 ),
    .B2(\i43/i47/n37 ),
    .Y(\i43/i47/n236 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i304  (.A1(\i43/i47/n32 ),
    .A2(\i43/i47/n64 ),
    .B1(\i43/i47/n42 ),
    .B2(\i43/i47/n82 ),
    .Y(\i43/i47/n234 ));
 AOI22xp5_ASAP7_75t_SL \i43/i47/i305  (.A1(\i43/i47/n93 ),
    .A2(\i43/i47/n67 ),
    .B1(\i43/i47/n43 ),
    .B2(\i43/i47/n69 ),
    .Y(\i43/i47/n232 ));
 AO22x1_ASAP7_75t_SL \i43/i47/i306  (.A1(\i43/i47/n33 ),
    .A2(\i43/i47/n34 ),
    .B1(\i43/i47/n57 ),
    .B2(\i43/i47/n81 ),
    .Y(\i43/i47/n231 ));
 AOI22xp5_ASAP7_75t_SL \i43/i47/i307  (.A1(\i43/i47/n73 ),
    .A2(\i43/i47/n79 ),
    .B1(\i43/i47/n53 ),
    .B2(\i43/i47/n69 ),
    .Y(\i43/i47/n230 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i308  (.A1(\i43/i47/n58 ),
    .A2(\i43/i47/n64 ),
    .B1(\i43/i47/n54 ),
    .B2(\i43/i47/n63 ),
    .Y(\i43/i47/n228 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i309  (.A(\i43/i47/n187 ),
    .B(\i43/i47/n188 ),
    .Y(\i43/i47/n193 ));
 NOR3xp33_ASAP7_75t_SL \i43/i47/i31  (.A(\i43/i47/n448 ),
    .B(\i43/i47/n436 ),
    .C(\i43/i47/n428 ),
    .Y(\i43/i47/n484 ));
 NAND2xp33_ASAP7_75t_SL \i43/i47/i310  (.A(\i43/i47/n186 ),
    .B(\i43/i47/n176 ),
    .Y(\i43/i47/n192 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i311  (.A1(\i43/i47/n92 ),
    .A2(\i43/i47/n40 ),
    .B1(\i43/i47/n76 ),
    .B2(\i43/i47/n70 ),
    .Y(\i43/i47/n227 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i312  (.A1(\i43/i47/n35 ),
    .A2(\i43/i47/n63 ),
    .B1(\i43/i47/n72 ),
    .B2(\i43/i47/n68 ),
    .Y(\i43/i47/n226 ));
 OAI22xp33_ASAP7_75t_SL \i43/i47/i313  (.A1(\i43/i47/n92 ),
    .A2(\i43/i47/n89 ),
    .B1(\i43/i47/n37 ),
    .B2(\i43/i47/n49 ),
    .Y(\i43/i47/n225 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i314  (.A1(\i43/i47/n92 ),
    .A2(\i43/i47/n49 ),
    .B1(\i43/i47/n42 ),
    .B2(\i43/i47/n75 ),
    .Y(\i43/i47/n224 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i315  (.A1(\i43/i47/n35 ),
    .A2(\i43/i47/n75 ),
    .B1(\i43/i47/n46 ),
    .B2(\i43/i47/n45 ),
    .Y(\i43/i47/n223 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i316  (.A1(\i43/i47/n80 ),
    .A2(\i43/i47/n39 ),
    .B1(\i43/i47/n54 ),
    .B2(\i43/i47/n68 ),
    .Y(\i43/i47/n221 ));
 AOI22xp5_ASAP7_75t_SL \i43/i47/i317  (.A1(\i43/i47/n33 ),
    .A2(\i43/i47/n57 ),
    .B1(\i43/i47/n41 ),
    .B2(\i43/i47/n36 ),
    .Y(\i43/i47/n220 ));
 OAI22xp33_ASAP7_75t_SL \i43/i47/i318  (.A1(\i43/i47/n87 ),
    .A2(\i43/i47/n89 ),
    .B1(\i43/i47/n78 ),
    .B2(\i43/i47/n42 ),
    .Y(\i43/i47/n219 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i319  (.A1(\i43/i47/n46 ),
    .A2(\i43/i47/n58 ),
    .B1(\i43/i47/n91 ),
    .B2(\i43/i47/n76 ),
    .Y(\i43/i47/n218 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i32  (.A(\i43/i47/n444 ),
    .B(\i43/i47/n474 ),
    .Y(\i43/i47/n483 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i320  (.A1(\i43/i47/n68 ),
    .A2(\i43/i47/n64 ),
    .B1(\i43/i47/n50 ),
    .B2(\i43/i47/n37 ),
    .Y(\i43/i47/n217 ));
 AOI22xp5_ASAP7_75t_SL \i43/i47/i321  (.A1(\i43/i47/n79 ),
    .A2(\i43/i47/n57 ),
    .B1(\i43/i47/n95 ),
    .B2(\i43/i47/n69 ),
    .Y(\i43/i47/n216 ));
 OAI22xp5_ASAP7_75t_SL \i43/i47/i322  (.A1(\i43/i47/n78 ),
    .A2(\i43/i47/n89 ),
    .B1(\i43/i47/n50 ),
    .B2(\i43/i47/n32 ),
    .Y(\i43/i47/n215 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i323  (.A(\i43/i47/n139 ),
    .B(\i43/i47/n138 ),
    .Y(\i43/i47/n191 ));
 AOI22xp5_ASAP7_75t_SL \i43/i47/i324  (.A1(\i43/i47/n93 ),
    .A2(\i43/i47/n34 ),
    .B1(\i43/i47/n77 ),
    .B2(\i43/i47/n62 ),
    .Y(\i43/i47/n214 ));
 OA22x2_ASAP7_75t_SL \i43/i47/i325  (.A1(\i43/i47/n61 ),
    .A2(\i43/i47/n64 ),
    .B1(\i43/i47/n58 ),
    .B2(\i43/i47/n76 ),
    .Y(\i43/i47/n213 ));
 INVx1_ASAP7_75t_SL \i43/i47/i326  (.A(\i43/i47/n189 ),
    .Y(\i43/i47/n190 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i327  (.A(\i43/i47/n182 ),
    .Y(\i43/i47/n183 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i328  (.A(\i43/i47/n176 ),
    .Y(\i43/i47/n177 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i329  (.A(\i43/i47/n174 ),
    .Y(\i43/i47/n175 ));
 NOR5xp2_ASAP7_75t_SL \i43/i47/i33  (.A(\i43/i47/n400 ),
    .B(\i43/i47/n408 ),
    .C(\i43/i47/n305 ),
    .D(\i43/i47/n397 ),
    .E(\i43/i47/n401 ),
    .Y(\i43/i47/n482 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i330  (.A(\i43/i47/n168 ),
    .Y(\i43/i47/n169 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i331  (.A(\i43/i47/n165 ),
    .Y(\i43/i47/n166 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i332  (.A(\i43/i47/n160 ),
    .Y(\i43/i47/n161 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i333  (.A(\i43/i47/n155 ),
    .Y(\i43/i47/n156 ));
 INVx1_ASAP7_75t_SL \i43/i47/i334  (.A(\i43/i47/n153 ),
    .Y(\i43/i47/n154 ));
 INVx1_ASAP7_75t_SL \i43/i47/i335  (.A(\i43/i47/n151 ),
    .Y(\i43/i47/n152 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i336  (.A(\i43/i47/n149 ),
    .Y(\i43/i47/n150 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i337  (.A(\i43/i47/n147 ),
    .Y(\i43/i47/n148 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i338  (.A(\i43/i47/n85 ),
    .B(\i43/i47/n51 ),
    .Y(\i43/i47/n146 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i339  (.A(\i43/i47/n77 ),
    .B(\i43/i47/n81 ),
    .Y(\i43/i47/n189 ));
 NAND5xp2_ASAP7_75t_SL \i43/i47/i34  (.A(\i43/i47/n390 ),
    .B(\i43/i47/n417 ),
    .C(\i43/i47/n352 ),
    .D(\i43/i47/n318 ),
    .E(\i43/i47/n349 ),
    .Y(\i43/i47/n481 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i340  (.A(\i43/i47/n41 ),
    .B(\i43/i47/n90 ),
    .Y(\i43/i47/n145 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i341  (.A(\i43/i47/n90 ),
    .B(\i43/i47/n48 ),
    .Y(\i43/i47/n144 ));
 NAND2xp33_ASAP7_75t_SL \i43/i47/i342  (.A(\i43/i47/n46 ),
    .B(\i43/i47/n64 ),
    .Y(\i43/i47/n143 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i343  (.A(\i43/i47/n36 ),
    .B(\i43/i47/n65 ),
    .Y(\i43/i47/n188 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i344  (.A(\i43/i47/n95 ),
    .B(\i43/i47/n93 ),
    .Y(\i43/i47/n187 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i345  (.A(\i43/i47/n67 ),
    .B(\i43/i47/n59 ),
    .Y(\i43/i47/n186 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i346  (.A(\i43/i47/n85 ),
    .B(\i43/i47/n71 ),
    .Y(\i43/i47/n142 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i347  (.A(\i43/i47/n58 ),
    .B(\i43/i47/n50 ),
    .Y(\i43/i47/n141 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i348  (.A(\i43/i47/n55 ),
    .B(\i43/i47/n83 ),
    .Y(\i43/i47/n185 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i349  (.A(\i43/i47/n69 ),
    .B(\i43/i47/n41 ),
    .Y(\i43/i47/n140 ));
 NOR2xp33_ASAP7_75t_L \i43/i47/i35  (.A(\i43/i47/n455 ),
    .B(\i43/i47/n478 ),
    .Y(\i43/i47/n480 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i350  (.A(\i43/i47/n77 ),
    .B(\i43/i47/n93 ),
    .Y(\i43/i47/n184 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i351  (.A(\i43/i47/n75 ),
    .B(\i43/i47/n40 ),
    .Y(\i43/i47/n182 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i352  (.A(\i43/i47/n69 ),
    .B(\i43/i47/n67 ),
    .Y(\i43/i47/n181 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i353  (.A(\i43/i47/n79 ),
    .B(\i43/i47/n51 ),
    .Y(\i43/i47/n180 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i354  (.A(\i43/i47/n93 ),
    .B(\i43/i47/n65 ),
    .Y(\i43/i47/n179 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i355  (.A(\i43/i47/n79 ),
    .B(\i43/i47/n95 ),
    .Y(\i43/i47/n178 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i356  (.A(\i43/i47/n74 ),
    .B(\i43/i47/n65 ),
    .Y(\i43/i47/n176 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i357  (.A(\i43/i47/n86 ),
    .B(\i43/i47/n77 ),
    .Y(\i43/i47/n174 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i358  (.A(\i43/i47/n85 ),
    .B(\i43/i47/n69 ),
    .Y(\i43/i47/n173 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i359  (.A(\i43/i47/n95 ),
    .B(\i43/i47/n36 ),
    .Y(\i43/i47/n172 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i36  (.A(\i43/i47/n416 ),
    .B(\i43/i47/n477 ),
    .Y(\i43/i47/n479 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i360  (.A(\i43/i47/n44 ),
    .B(\i43/i47/n65 ),
    .Y(\i43/i47/n171 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i361  (.A(\i43/i47/n91 ),
    .B(\i43/i47/n46 ),
    .Y(\i43/i47/n170 ));
 NAND2xp5_ASAP7_75t_L \i43/i47/i362  (.A(\i43/i47/n35 ),
    .B(\i43/i47/n94 ),
    .Y(\i43/i47/n168 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i363  (.A(\i43/i47/n95 ),
    .B(\i43/i47/n33 ),
    .Y(\i43/i47/n167 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i364  (.A(\i43/i47/n95 ),
    .B(\i43/i47/n43 ),
    .Y(\i43/i47/n165 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i365  (.A(\i43/i47/n57 ),
    .B(\i43/i47/n59 ),
    .Y(\i43/i47/n164 ));
 NAND2xp33_ASAP7_75t_SL \i43/i47/i366  (.A(\i43/i47/n61 ),
    .B(\i43/i47/n87 ),
    .Y(\i43/i47/n163 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i367  (.A(\i43/i47/n59 ),
    .B(\i43/i47/n41 ),
    .Y(\i43/i47/n162 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i368  (.A(\i43/i47/n73 ),
    .B(\i43/i47/n59 ),
    .Y(\i43/i47/n160 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i369  (.A(\i43/i47/n77 ),
    .B(\i43/i47/n83 ),
    .Y(\i43/i47/n159 ));
 INVx1_ASAP7_75t_SL \i43/i47/i37  (.A(\i43/i47/n509 ),
    .Y(\i43/i47/n475 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i370  (.A(\i43/i47/n85 ),
    .B(\i43/i47/n57 ),
    .Y(\i43/i47/n158 ));
 NOR2xp33_ASAP7_75t_L \i43/i47/i371  (.A(\i43/i47/n60 ),
    .B(\i43/i47/n69 ),
    .Y(\i43/i47/n157 ));
 NAND2xp5_ASAP7_75t_L \i43/i47/i372  (.A(\i43/i47/n37 ),
    .B(\i43/i47/n68 ),
    .Y(\i43/i47/n155 ));
 NOR2x1_ASAP7_75t_SL \i43/i47/i373  (.A(\i43/i47/n62 ),
    .B(\i43/i47/n71 ),
    .Y(\i43/i47/n153 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i374  (.A(\i43/i47/n88 ),
    .B(\i43/i47/n36 ),
    .Y(\i43/i47/n151 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i375  (.A(\i43/i47/n86 ),
    .B(\i43/i47/n62 ),
    .Y(\i43/i47/n149 ));
 NAND2x1_ASAP7_75t_SL \i43/i47/i376  (.A(\i43/i47/n84 ),
    .B(\i43/i47/n63 ),
    .Y(\i43/i47/n0 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i377  (.A(\i43/i47/n32 ),
    .B(\i43/i47/n91 ),
    .Y(\i43/i47/n147 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i378  (.A(\i43/i47/n130 ),
    .Y(\i43/i47/n131 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i379  (.A(\i43/i47/n121 ),
    .Y(\i43/i47/n122 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i38  (.A(\i43/i47/n453 ),
    .B(\i43/i47/n422 ),
    .Y(\i43/i47/n473 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i380  (.A(\i43/i47/n118 ),
    .Y(\i43/i47/n119 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i381  (.A(\i43/i47/n55 ),
    .B(\i43/i47/n36 ),
    .Y(\i43/i47/n116 ));
 NAND2xp33_ASAP7_75t_SL \i43/i47/i382  (.A(\i43/i47/n70 ),
    .B(\i43/i47/n61 ),
    .Y(\i43/i47/n115 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i383  (.A(\i43/i47/n48 ),
    .B(\i43/i47/n57 ),
    .Y(\i43/i47/n114 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i384  (.A(\i43/i47/n51 ),
    .B(\i43/i47/n83 ),
    .Y(\i43/i47/n113 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i385  (.A(\i43/i47/n57 ),
    .B(\i43/i47/n36 ),
    .Y(\i43/i47/n139 ));
 NAND2xp33_ASAP7_75t_SL \i43/i47/i386  (.A(\i43/i47/n82 ),
    .B(\i43/i47/n45 ),
    .Y(\i43/i47/n112 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i387  (.A(\i43/i47/n71 ),
    .B(\i43/i47/n55 ),
    .Y(\i43/i47/n111 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i388  (.A(\i43/i47/n33 ),
    .B(\i43/i47/n38 ),
    .Y(\i43/i47/n110 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i389  (.A(\i43/i47/n75 ),
    .B(\i43/i47/n82 ),
    .Y(\i43/i47/n109 ));
 NAND2xp33_ASAP7_75t_L \i43/i47/i39  (.A(\i43/i47/n453 ),
    .B(\i43/i47/n433 ),
    .Y(\i43/i47/n472 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i390  (.A(\i43/i47/n93 ),
    .B(\i43/i47/n53 ),
    .Y(\i43/i47/n108 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i391  (.A(\i43/i47/n44 ),
    .B(\i43/i47/n43 ),
    .Y(\i43/i47/n138 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i392  (.A(\i43/i47/n60 ),
    .B(\i43/i47/n34 ),
    .Y(\i43/i47/n107 ));
 NAND2xp33_ASAP7_75t_SL \i43/i47/i393  (.A(\i43/i47/n39 ),
    .B(\i43/i47/n66 ),
    .Y(\i43/i47/n106 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i394  (.A(\i43/i47/n47 ),
    .B(\i43/i47/n33 ),
    .Y(\i43/i47/n105 ));
 NAND2xp5_ASAP7_75t_L \i43/i47/i395  (.A(\i43/i47/n42 ),
    .B(\i43/i47/n66 ),
    .Y(\i43/i47/n104 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i396  (.A(\i43/i47/n38 ),
    .B(\i43/i47/n73 ),
    .Y(\i43/i47/n103 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i397  (.A(\i43/i47/n73 ),
    .B(\i43/i47/n60 ),
    .Y(\i43/i47/n137 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i398  (.A(\i43/i47/n41 ),
    .B(\i43/i47/n73 ),
    .Y(\i43/i47/n136 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i399  (.A(\i43/i47/n74 ),
    .B(\i43/i47/n48 ),
    .Y(\i43/i47/n135 ));
 AND5x1_ASAP7_75t_SL \i43/i47/i4  (.A(\i43/i47/n501 ),
    .B(\i43/i47/n498 ),
    .C(\i43/i47/n477 ),
    .D(\i43/i47/n499 ),
    .E(\i43/i47/n468 ),
    .Y(\i43/n0 [19]));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i40  (.A(\i43/i47/n450 ),
    .B(\i43/i47/n432 ),
    .Y(\i43/i47/n471 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i400  (.A(\i43/i47/n72 ),
    .B(\i43/i47/n45 ),
    .Y(\i43/i47/n102 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i401  (.A(\i43/i47/n67 ),
    .B(\i43/i47/n36 ),
    .Y(\i43/i47/n134 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i402  (.A(\i43/i47/n47 ),
    .B(\i43/i47/n93 ),
    .Y(\i43/i47/n133 ));
 NOR2xp33_ASAP7_75t_L \i43/i47/i403  (.A(\i43/i47/n35 ),
    .B(\i43/i47/n37 ),
    .Y(\i43/i47/n132 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i404  (.A(\i43/i47/n42 ),
    .B(\i43/i47/n75 ),
    .Y(\i43/i47/n101 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i405  (.A(\i43/i47/n71 ),
    .B(\i43/i47/n34 ),
    .Y(\i43/i47/n100 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i406  (.A(\i43/i47/n51 ),
    .B(\i43/i47/n44 ),
    .Y(\i43/i47/n130 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i407  (.A(\i43/i47/n92 ),
    .B(\i43/i47/n42 ),
    .Y(\i43/i47/n129 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i408  (.A(\i43/i47/n47 ),
    .B(\i43/i47/n81 ),
    .Y(\i43/i47/n128 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i409  (.A(\i43/i47/n47 ),
    .B(\i43/i47/n60 ),
    .Y(\i43/i47/n127 ));
 NAND4xp25_ASAP7_75t_SL \i43/i47/i41  (.A(\i43/i47/n415 ),
    .B(\i43/i47/n308 ),
    .C(\i43/i47/n311 ),
    .D(\i43/i47/n343 ),
    .Y(\i43/i47/n470 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i410  (.A(\i43/i47/n74 ),
    .B(\i43/i47/n51 ),
    .Y(\i43/i47/n126 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i411  (.A(\i43/i47/n38 ),
    .B(\i43/i47/n93 ),
    .Y(\i43/i47/n99 ));
 NOR2xp33_ASAP7_75t_L \i43/i47/i412  (.A(\i43/i47/n50 ),
    .B(\i43/i47/n80 ),
    .Y(\i43/i47/n125 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i413  (.A(\i43/i47/n50 ),
    .B(\i43/i47/n92 ),
    .Y(\i43/i47/n98 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i414  (.A(\i43/i47/n61 ),
    .B(\i43/i47/n42 ),
    .Y(\i43/i47/n97 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i415  (.A(\i43/i47/n93 ),
    .B(\i43/i47/n57 ),
    .Y(\i43/i47/n124 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i416  (.A(\i43/i47/n55 ),
    .B(\i43/i47/n44 ),
    .Y(\i43/i47/n96 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i417  (.A(\i43/i47/n79 ),
    .B(\i43/i47/n38 ),
    .Y(\i43/i47/n123 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i418  (.A(\i43/i47/n49 ),
    .B(\i43/i47/n32 ),
    .Y(\i43/i47/n121 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i419  (.A(\i43/i47/n33 ),
    .B(\i43/i47/n53 ),
    .Y(\i43/i47/n120 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i42  (.A(\i43/i47/n433 ),
    .B(\i43/i47/n442 ),
    .Y(\i43/i47/n478 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i420  (.A(\i43/i47/n83 ),
    .B(\i43/i47/n53 ),
    .Y(\i43/i47/n118 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i421  (.A(\i43/i47/n60 ),
    .B(\i43/i47/n51 ),
    .Y(\i43/i47/n117 ));
 INVx1_ASAP7_75t_SL \i43/i47/i422  (.A(\i43/i47/n95 ),
    .Y(\i43/i47/n94 ));
 INVx2_ASAP7_75t_SL \i43/i47/i423  (.A(\i43/i47/n93 ),
    .Y(\i43/i47/n92 ));
 INVx1_ASAP7_75t_SL \i43/i47/i424  (.A(\i43/i47/n91 ),
    .Y(\i43/i47/n90 ));
 INVx2_ASAP7_75t_SL \i43/i47/i425  (.A(\i43/i47/n89 ),
    .Y(\i43/i47/n88 ));
 INVx2_ASAP7_75t_SL \i43/i47/i426  (.A(\i43/i47/n87 ),
    .Y(\i43/i47/n86 ));
 INVx2_ASAP7_75t_SL \i43/i47/i427  (.A(\i43/i47/n85 ),
    .Y(\i43/i47/n84 ));
 INVx3_ASAP7_75t_SL \i43/i47/i428  (.A(\i43/i47/n83 ),
    .Y(\i43/i47/n82 ));
 INVx2_ASAP7_75t_SL \i43/i47/i429  (.A(\i43/i47/n81 ),
    .Y(\i43/i47/n80 ));
 AND4x1_ASAP7_75t_SL \i43/i47/i43  (.A(\i43/i47/n435 ),
    .B(\i43/i47/n415 ),
    .C(\i43/i47/n353 ),
    .D(\i43/i47/n193 ),
    .Y(\i43/i47/n469 ));
 INVx2_ASAP7_75t_SL \i43/i47/i430  (.A(\i43/i47/n79 ),
    .Y(\i43/i47/n78 ));
 INVx2_ASAP7_75t_SL \i43/i47/i431  (.A(\i43/i47/n77 ),
    .Y(\i43/i47/n76 ));
 INVx2_ASAP7_75t_SL \i43/i47/i432  (.A(\i43/i47/n75 ),
    .Y(\i43/i47/n74 ));
 INVx2_ASAP7_75t_SL \i43/i47/i433  (.A(\i43/i47/n73 ),
    .Y(\i43/i47/n72 ));
 INVx2_ASAP7_75t_SL \i43/i47/i434  (.A(\i43/i47/n71 ),
    .Y(\i43/i47/n70 ));
 INVx2_ASAP7_75t_SL \i43/i47/i435  (.A(\i43/i47/n69 ),
    .Y(\i43/i47/n68 ));
 INVx2_ASAP7_75t_SL \i43/i47/i436  (.A(\i43/i47/n67 ),
    .Y(\i43/i47/n66 ));
 INVx2_ASAP7_75t_SL \i43/i47/i437  (.A(\i43/i47/n65 ),
    .Y(\i43/i47/n64 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i438  (.A(\i43/i47/n25 ),
    .B(\i43/i47/n15 ),
    .Y(\i43/i47/n95 ));
 AND2x4_ASAP7_75t_SL \i43/i47/i439  (.A(\i43/i47/n5 ),
    .B(\i43/i47/n6 ),
    .Y(\i43/i47/n93 ));
 AND4x1_ASAP7_75t_SL \i43/i47/i44  (.A(\i43/i47/n380 ),
    .B(\i43/i47/n317 ),
    .C(\i43/i47/n368 ),
    .D(\i43/i47/n189 ),
    .Y(\i43/i47/n477 ));
 OR2x2_ASAP7_75t_SL \i43/i47/i440  (.A(\i43/i47/n27 ),
    .B(\i43/i47/n11 ),
    .Y(\i43/i47/n91 ));
 OR2x2_ASAP7_75t_SL \i43/i47/i441  (.A(\i43/i47/n28 ),
    .B(\i43/i47/n9 ),
    .Y(\i43/i47/n89 ));
 OR2x6_ASAP7_75t_SL \i43/i47/i442  (.A(\i43/i47/n7 ),
    .B(\i43/i47/n11 ),
    .Y(\i43/i47/n87 ));
 AND2x4_ASAP7_75t_SL \i43/i47/i443  (.A(\i43/i47/n4 ),
    .B(\i43/i47/n19 ),
    .Y(\i43/i47/n85 ));
 AND2x4_ASAP7_75t_SL \i43/i47/i444  (.A(\i43/i47/n10 ),
    .B(\i43/i47/n22 ),
    .Y(\i43/i47/n83 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i445  (.A(\i43/i47/n6 ),
    .B(\i43/i47/n19 ),
    .Y(\i43/i47/n81 ));
 AND2x4_ASAP7_75t_SL \i43/i47/i446  (.A(\i43/i47/n5 ),
    .B(\i43/i47/n26 ),
    .Y(\i43/i47/n79 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i447  (.A(\i43/i47/n16 ),
    .B(\i43/i47/n15 ),
    .Y(\i43/i47/n77 ));
 OR2x2_ASAP7_75t_SL \i43/i47/i448  (.A(\i43/i47/n3 ),
    .B(\i43/i47/n31 ),
    .Y(\i43/i47/n75 ));
 AND2x4_ASAP7_75t_SL \i43/i47/i449  (.A(\i43/i47/n25 ),
    .B(\i43/i47/n12 ),
    .Y(\i43/i47/n73 ));
 NOR2x1_ASAP7_75t_SL \i43/i47/i45  (.A(\i43/i47/n306 ),
    .B(\i43/i47/n451 ),
    .Y(\i43/i47/n476 ));
 AND2x4_ASAP7_75t_SL \i43/i47/i450  (.A(\i43/i47/n4 ),
    .B(\i43/i47/n10 ),
    .Y(\i43/i47/n71 ));
 AND2x4_ASAP7_75t_SL \i43/i47/i451  (.A(\i43/i47/n5 ),
    .B(\i43/i47/n4 ),
    .Y(\i43/i47/n69 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i452  (.A(\i43/i47/n16 ),
    .B(\i43/i47/n29 ),
    .Y(\i43/i47/n67 ));
 AND2x4_ASAP7_75t_SL \i43/i47/i453  (.A(\i43/i47/n8 ),
    .B(\i43/i47/n12 ),
    .Y(\i43/i47/n65 ));
 INVx2_ASAP7_75t_SL \i43/i47/i454  (.A(\i43/i47/n63 ),
    .Y(\i43/i47/n62 ));
 INVx3_ASAP7_75t_SL \i43/i47/i455  (.A(\i43/i47/n61 ),
    .Y(\i43/i47/n60 ));
 INVx2_ASAP7_75t_SL \i43/i47/i456  (.A(\i43/i47/n59 ),
    .Y(\i43/i47/n58 ));
 INVx1_ASAP7_75t_SL \i43/i47/i457  (.A(\i43/i47/n57 ),
    .Y(\i43/i47/n56 ));
 INVx2_ASAP7_75t_SL \i43/i47/i458  (.A(\i43/i47/n55 ),
    .Y(\i43/i47/n54 ));
 INVx3_ASAP7_75t_SL \i43/i47/i459  (.A(\i43/i47/n53 ),
    .Y(\i43/i47/n52 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i46  (.A(\i43/i47/n392 ),
    .B(\i43/i47/n426 ),
    .Y(\i43/i47/n474 ));
 INVx2_ASAP7_75t_SL \i43/i47/i460  (.A(\i43/i47/n51 ),
    .Y(\i43/i47/n50 ));
 INVx2_ASAP7_75t_SL \i43/i47/i461  (.A(\i43/i47/n49 ),
    .Y(\i43/i47/n48 ));
 INVx2_ASAP7_75t_SL \i43/i47/i462  (.A(\i43/i47/n47 ),
    .Y(\i43/i47/n46 ));
 INVx4_ASAP7_75t_SL \i43/i47/i463  (.A(\i43/i47/n45 ),
    .Y(\i43/i47/n44 ));
 INVx4_ASAP7_75t_SL \i43/i47/i464  (.A(\i43/i47/n43 ),
    .Y(\i43/i47/n42 ));
 INVx2_ASAP7_75t_SL \i43/i47/i465  (.A(\i43/i47/n41 ),
    .Y(\i43/i47/n40 ));
 INVx2_ASAP7_75t_SL \i43/i47/i466  (.A(\i43/i47/n39 ),
    .Y(\i43/i47/n38 ));
 INVx2_ASAP7_75t_SL \i43/i47/i467  (.A(\i43/i47/n37 ),
    .Y(\i43/i47/n36 ));
 INVx3_ASAP7_75t_SL \i43/i47/i468  (.A(\i43/i47/n35 ),
    .Y(\i43/i47/n34 ));
 INVx2_ASAP7_75t_SL \i43/i47/i469  (.A(\i43/i47/n33 ),
    .Y(\i43/i47/n32 ));
 INVx1_ASAP7_75t_SL \i43/i47/i47  (.A(\i43/i47/n466 ),
    .Y(\i43/i47/n467 ));
 NAND2x1p5_ASAP7_75t_SL \i43/i47/i470  (.A(\i43/i47/n22 ),
    .B(\i43/i47/n5 ),
    .Y(\i43/i47/n63 ));
 OR2x2_ASAP7_75t_SL \i43/i47/i471  (.A(\i43/i47/n27 ),
    .B(\i43/i47/n20 ),
    .Y(\i43/i47/n61 ));
 AND2x4_ASAP7_75t_SL \i43/i47/i472  (.A(\i43/i47/n6 ),
    .B(\i43/i47/n30 ),
    .Y(\i43/i47/n59 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i473  (.A(\i43/i47/n25 ),
    .B(\i43/i47/n18 ),
    .Y(\i43/i47/n57 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i474  (.A(\i43/i47/n8 ),
    .B(\i43/i47/n18 ),
    .Y(\i43/i47/n55 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i475  (.A(\i43/i47/n16 ),
    .B(\i43/i47/n12 ),
    .Y(\i43/i47/n53 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i476  (.A(\i43/i47/n25 ),
    .B(\i43/i47/n29 ),
    .Y(\i43/i47/n51 ));
 OR2x2_ASAP7_75t_SL \i43/i47/i477  (.A(\i43/i47/n17 ),
    .B(\i43/i47/n24 ),
    .Y(\i43/i47/n49 ));
 AND2x4_ASAP7_75t_SL \i43/i47/i478  (.A(\i43/i47/n23 ),
    .B(\i43/i47/n15 ),
    .Y(\i43/i47/n47 ));
 OR2x2_ASAP7_75t_SL \i43/i47/i479  (.A(\i43/i47/n27 ),
    .B(\i43/i47/n31 ),
    .Y(\i43/i47/n45 ));
 NAND2xp5_ASAP7_75t_L \i43/i47/i48  (.A(\i43/i47/n435 ),
    .B(\i43/i47/n419 ),
    .Y(\i43/i47/n464 ));
 AND2x4_ASAP7_75t_SL \i43/i47/i480  (.A(\i43/i47/n23 ),
    .B(\i43/i47/n29 ),
    .Y(\i43/i47/n43 ));
 AND2x4_ASAP7_75t_SL \i43/i47/i481  (.A(\i43/i47/n16 ),
    .B(\i43/i47/n18 ),
    .Y(\i43/i47/n41 ));
 OR2x2_ASAP7_75t_SL \i43/i47/i482  (.A(\i43/i47/n14 ),
    .B(\i43/i47/n9 ),
    .Y(\i43/i47/n39 ));
 OR2x6_ASAP7_75t_SL \i43/i47/i483  (.A(\i43/i47/n20 ),
    .B(\i43/i47/n21 ),
    .Y(\i43/i47/n37 ));
 OR2x6_ASAP7_75t_SL \i43/i47/i484  (.A(\i43/i47/n24 ),
    .B(\i43/i47/n13 ),
    .Y(\i43/i47/n35 ));
 AND2x4_ASAP7_75t_SL \i43/i47/i485  (.A(\i43/i47/n30 ),
    .B(\i43/i47/n22 ),
    .Y(\i43/i47/n33 ));
 INVx2_ASAP7_75t_SL \i43/i47/i486  (.A(\i43/i47/n31 ),
    .Y(\i43/i47/n30 ));
 INVx2_ASAP7_75t_SL \i43/i47/i487  (.A(\i43/i47/n28 ),
    .Y(\i43/i47/n29 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i488  (.A(\i43/i47/n27 ),
    .Y(\i43/i47/n26 ));
 INVx2_ASAP7_75t_SL \i43/i47/i489  (.A(\i43/i47/n24 ),
    .Y(\i43/i47/n23 ));
 AND3x1_ASAP7_75t_SL \i43/i47/i49  (.A(\i43/i47/n420 ),
    .B(\i43/i47/n405 ),
    .C(\i43/i47/n391 ),
    .Y(\i43/i47/n463 ));
 INVx3_ASAP7_75t_SL \i43/i47/i490  (.A(\i43/i47/n21 ),
    .Y(\i43/i47/n22 ));
 INVx2_ASAP7_75t_SL \i43/i47/i491  (.A(\i43/i47/n20 ),
    .Y(\i43/i47/n19 ));
 INVx1_ASAP7_75t_SL \i43/i47/i492  (.A(\i43/i47/n17 ),
    .Y(\i43/i47/n18 ));
 OR2x2_ASAP7_75t_SL \i43/i47/i493  (.A(n72),
    .B(n34[13]),
    .Y(\i43/i47/n31 ));
 OR2x2_ASAP7_75t_SL \i43/i47/i494  (.A(n73),
    .B(n34[8]),
    .Y(\i43/i47/n28 ));
 OR2x2_ASAP7_75t_SL \i43/i47/i495  (.A(n71),
    .B(n34[15]),
    .Y(\i43/i47/n27 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i496  (.A(n34[9]),
    .B(n74),
    .Y(\i43/i47/n25 ));
 NAND2x1_ASAP7_75t_SL \i43/i47/i497  (.A(n34[10]),
    .B(n75),
    .Y(\i43/i47/n24 ));
 OR2x2_ASAP7_75t_SL \i43/i47/i498  (.A(n70),
    .B(n34[14]),
    .Y(\i43/i47/n21 ));
 OR2x2_ASAP7_75t_SL \i43/i47/i499  (.A(\i43/i47/n2 ),
    .B(n34[12]),
    .Y(\i43/i47/n20 ));
 NAND5xp2_ASAP7_75t_SL \i43/i47/i5  (.A(\i43/i47/n466 ),
    .B(\i43/i47/n476 ),
    .C(\i43/i47/n471 ),
    .D(\i43/i47/n460 ),
    .E(\i43/i47/n454 ),
    .Y(\i43/i47/n507 ));
 NAND4xp25_ASAP7_75t_SL \i43/i47/i50  (.A(\i43/i47/n418 ),
    .B(\i43/i47/n384 ),
    .C(\i43/i47/n312 ),
    .D(\i43/i47/n309 ),
    .Y(\i43/i47/n462 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i500  (.A(n34[8]),
    .B(n73),
    .Y(\i43/i47/n17 ));
 INVx1_ASAP7_75t_SL \i43/i47/i501  (.A(\i43/i47/n14 ),
    .Y(\i43/i47/n15 ));
 INVx2_ASAP7_75t_SL \i43/i47/i502  (.A(\i43/i47/n12 ),
    .Y(\i43/i47/n13 ));
 INVx1_ASAP7_75t_SL \i43/i47/i503  (.A(\i43/i47/n11 ),
    .Y(\i43/i47/n10 ));
 INVx1_ASAP7_75t_SL \i43/i47/i504  (.A(\i43/i47/n9 ),
    .Y(\i43/i47/n8 ));
 INVx1_ASAP7_75t_SL \i43/i47/i505  (.A(\i43/i47/n6 ),
    .Y(\i43/i47/n7 ));
 INVx2_ASAP7_75t_SL \i43/i47/i506  (.A(\i43/i47/n3 ),
    .Y(\i43/i47/n4 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i507  (.A(n34[10]),
    .B(n34[9]),
    .Y(\i43/i47/n16 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i508  (.A(n34[11]),
    .B(n34[8]),
    .Y(\i43/i47/n14 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i509  (.A(n73),
    .B(n76),
    .Y(\i43/i47/n12 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i51  (.A(\i43/i47/n247 ),
    .B(\i43/i47/n510 ),
    .Y(\i43/i47/n461 ));
 OR2x2_ASAP7_75t_SL \i43/i47/i510  (.A(n34[13]),
    .B(n34[12]),
    .Y(\i43/i47/n11 ));
 OR2x2_ASAP7_75t_SL \i43/i47/i511  (.A(n34[10]),
    .B(n34[9]),
    .Y(\i43/i47/n9 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i512  (.A(n70),
    .B(n71),
    .Y(\i43/i47/n6 ));
 AND2x2_ASAP7_75t_SL \i43/i47/i513  (.A(n34[13]),
    .B(n34[12]),
    .Y(\i43/i47/n5 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i514  (.A(n34[15]),
    .B(n34[14]),
    .Y(\i43/i47/n3 ));
 INVxp67_ASAP7_75t_SL \i43/i47/i515  (.A(n34[13]),
    .Y(\i43/i47/n2 ));
 OR4x1_ASAP7_75t_SL \i43/i47/i516  (.A(\i43/i47/n450 ),
    .B(\i43/i47/n278 ),
    .C(\i43/i47/n248 ),
    .D(\i43/i47/n226 ),
    .Y(\i43/i47/n508 ));
 NAND5xp2_ASAP7_75t_SL \i43/i47/i517  (.A(\i43/i47/n452 ),
    .B(\i43/i47/n288 ),
    .C(\i43/i47/n277 ),
    .D(\i43/i47/n220 ),
    .E(\i43/i47/n414 ),
    .Y(\i43/i47/n509 ));
 AND3x1_ASAP7_75t_SL \i43/i47/i518  (.A(\i43/i47/n326 ),
    .B(\i43/i47/n267 ),
    .C(\i43/i47/n329 ),
    .Y(\i43/i47/n510 ));
 OR3x1_ASAP7_75t_SL \i43/i47/i519  (.A(\i43/i47/n223 ),
    .B(\i43/i47/n132 ),
    .C(\i43/i47/n199 ),
    .Y(\i43/i47/n511 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i52  (.A(\i43/i47/n411 ),
    .B(\i43/i47/n441 ),
    .Y(\i43/i47/n460 ));
 NAND3xp33_ASAP7_75t_SL \i43/i47/i520  (.A(\i43/i47/n230 ),
    .B(\i43/i47/n117 ),
    .C(\i43/i47/n107 ),
    .Y(\i43/i47/n512 ));
 NAND3xp33_ASAP7_75t_SL \i43/i47/i521  (.A(\i43/i47/n513 ),
    .B(\i43/i47/n302 ),
    .C(\i43/i47/n151 ),
    .Y(\i43/i47/n514 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i522  (.A(\i43/i47/n228 ),
    .B(\i43/i47/n124 ),
    .Y(\i43/i47/n513 ));
 NOR3xp33_ASAP7_75t_SL \i43/i47/i53  (.A(\i43/i47/n383 ),
    .B(\i43/i47/n398 ),
    .C(\i43/i47/n304 ),
    .Y(\i43/i47/n459 ));
 AOI211xp5_ASAP7_75t_SL \i43/i47/i54  (.A1(\i43/i47/n378 ),
    .A2(\i43/i47/n4 ),
    .B(\i43/i47/n394 ),
    .C(\i43/i47/n396 ),
    .Y(\i43/i47/n458 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i55  (.A(\i43/i47/n425 ),
    .B(\i43/i47/n431 ),
    .Y(\i43/i47/n457 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i56  (.A(\i43/i47/n393 ),
    .B(\i43/i47/n434 ),
    .Y(\i43/i47/n456 ));
 NOR2xp33_ASAP7_75t_L \i43/i47/i57  (.A(\i43/i47/n411 ),
    .B(\i43/i47/n430 ),
    .Y(\i43/i47/n468 ));
 OA211x2_ASAP7_75t_SL \i43/i47/i58  (.A1(\i43/i47/n91 ),
    .A2(\i43/i47/n66 ),
    .B(\i43/i47/n391 ),
    .C(\i43/i47/n370 ),
    .Y(\i43/i47/n466 ));
 NAND3xp33_ASAP7_75t_SL \i43/i47/i59  (.A(\i43/i47/n353 ),
    .B(\i43/i47/n379 ),
    .C(\i43/i47/n320 ),
    .Y(\i43/i47/n465 ));
 AND4x1_ASAP7_75t_SL \i43/i47/i6  (.A(\i43/i47/n495 ),
    .B(\i43/i47/n499 ),
    .C(\i43/i47/n484 ),
    .D(\i43/i47/n457 ),
    .Y(\i43/n0 [16]));
 INVxp67_ASAP7_75t_SL \i43/i47/i60  (.A(\i43/i47/n510 ),
    .Y(\i43/i47/n449 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i61  (.A(\i43/i47/n407 ),
    .B(\i43/i47/n392 ),
    .Y(\i43/i47/n448 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i62  (.A(\i43/i47/n300 ),
    .B(\i43/i47/n407 ),
    .Y(\i43/i47/n447 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i63  (.A(\i43/i47/n390 ),
    .B(\i43/i47/n387 ),
    .Y(\i43/i47/n455 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i64  (.A(\i43/i47/n511 ),
    .B(\i43/i47/n382 ),
    .Y(\i43/i47/n446 ));
 NAND2xp5_ASAP7_75t_L \i43/i47/i65  (.A(\i43/i47/n388 ),
    .B(\i43/i47/n310 ),
    .Y(\i43/i47/n445 ));
 NOR3xp33_ASAP7_75t_SL \i43/i47/i66  (.A(\i43/i47/n413 ),
    .B(\i43/i47/n342 ),
    .C(\i43/i47/n344 ),
    .Y(\i43/i47/n454 ));
 NAND3xp33_ASAP7_75t_SL \i43/i47/i67  (.A(\i43/i47/n389 ),
    .B(\i43/i47/n341 ),
    .C(\i43/i47/n216 ),
    .Y(\i43/i47/n444 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i68  (.A(\i43/i47/n299 ),
    .B(\i43/i47/n374 ),
    .Y(\i43/i47/n443 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i69  (.A(\i43/i47/n386 ),
    .B(\i43/i47/n512 ),
    .Y(\i43/i47/n442 ));
 AND4x1_ASAP7_75t_L \i43/i47/i7  (.A(\i43/i47/n485 ),
    .B(\i43/i47/n490 ),
    .C(\i43/i47/n498 ),
    .D(\i43/i47/n487 ),
    .Y(\i43/n0 [23]));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i70  (.A(\i43/i47/n353 ),
    .B(\i43/i47/n399 ),
    .Y(\i43/i47/n441 ));
 OA211x2_ASAP7_75t_SL \i43/i47/i71  (.A1(\i43/i47/n66 ),
    .A2(\i43/i47/n87 ),
    .B(\i43/i47/n365 ),
    .C(\i43/i47/n368 ),
    .Y(\i43/i47/n440 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i72  (.A(\i43/i47/n514 ),
    .B(\i43/i47/n403 ),
    .Y(\i43/i47/n439 ));
 AND3x1_ASAP7_75t_SL \i43/i47/i73  (.A(\i43/i47/n352 ),
    .B(\i43/i47/n363 ),
    .C(\i43/i47/n348 ),
    .Y(\i43/i47/n438 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i74  (.A(\i43/i47/n377 ),
    .B(\i43/i47/n364 ),
    .Y(\i43/i47/n453 ));
 NOR3xp33_ASAP7_75t_SL \i43/i47/i75  (.A(\i43/i47/n327 ),
    .B(\i43/i47/n361 ),
    .C(\i43/i47/n201 ),
    .Y(\i43/i47/n452 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i76  (.A(\i43/i47/n323 ),
    .B(\i43/i47/n381 ),
    .Y(\i43/i47/n451 ));
 NAND2xp33_ASAP7_75t_SL \i43/i47/i77  (.A(\i43/i47/n368 ),
    .B(\i43/i47/n389 ),
    .Y(\i43/i47/n437 ));
 NAND3xp33_ASAP7_75t_SL \i43/i47/i78  (.A(\i43/i47/n318 ),
    .B(\i43/i47/n355 ),
    .C(\i43/i47/n295 ),
    .Y(\i43/i47/n450 ));
 NAND2xp33_ASAP7_75t_SL \i43/i47/i79  (.A(\i43/i47/n370 ),
    .B(\i43/i47/n391 ),
    .Y(\i43/i47/n436 ));
 NAND4xp25_ASAP7_75t_SL \i43/i47/i8  (.A(\i43/i47/n486 ),
    .B(\i43/i47/n488 ),
    .C(\i43/i47/n475 ),
    .D(\i43/i47/n463 ),
    .Y(\i43/i47/n506 ));
 NAND2xp33_ASAP7_75t_SL \i43/i47/i80  (.A(\i43/i47/n406 ),
    .B(\i43/i47/n414 ),
    .Y(\i43/i47/n432 ));
 NAND4xp25_ASAP7_75t_SL \i43/i47/i81  (.A(\i43/i47/n323 ),
    .B(\i43/i47/n326 ),
    .C(\i43/i47/n294 ),
    .D(\i43/i47/n360 ),
    .Y(\i43/i47/n431 ));
 NAND3xp33_ASAP7_75t_SL \i43/i47/i82  (.A(\i43/i47/n322 ),
    .B(\i43/i47/n291 ),
    .C(\i43/i47/n276 ),
    .Y(\i43/i47/n430 ));
 NAND2xp5_ASAP7_75t_SL \i43/i47/i83  (.A(\i43/i47/n317 ),
    .B(\i43/i47/n385 ),
    .Y(\i43/i47/n429 ));
 NAND5xp2_ASAP7_75t_SL \i43/i47/i84  (.A(\i43/i47/n355 ),
    .B(\i43/i47/n214 ),
    .C(\i43/i47/n339 ),
    .D(\i43/i47/n235 ),
    .E(\i43/i47/n229 ),
    .Y(\i43/i47/n428 ));
 AOI211xp5_ASAP7_75t_SL \i43/i47/i85  (.A1(\i43/i47/n243 ),
    .A2(\i43/i47/n47 ),
    .B(\i43/i47/n284 ),
    .C(\i43/i47/n275 ),
    .Y(\i43/i47/n427 ));
 NOR2xp33_ASAP7_75t_L \i43/i47/i86  (.A(\i43/i47/n376 ),
    .B(\i43/i47/n409 ),
    .Y(\i43/i47/n426 ));
 NAND5xp2_ASAP7_75t_SL \i43/i47/i87  (.A(\i43/i47/n319 ),
    .B(\i43/i47/n367 ),
    .C(\i43/i47/n230 ),
    .D(\i43/i47/n127 ),
    .E(\i43/i47/n110 ),
    .Y(\i43/i47/n425 ));
 NAND4xp25_ASAP7_75t_SL \i43/i47/i88  (.A(\i43/i47/n352 ),
    .B(\i43/i47/n366 ),
    .C(\i43/i47/n345 ),
    .D(\i43/i47/n285 ),
    .Y(\i43/i47/n424 ));
 NOR2xp33_ASAP7_75t_SL \i43/i47/i89  (.A(\i43/i47/n346 ),
    .B(\i43/i47/n373 ),
    .Y(\i43/i47/n423 ));
 NAND4xp25_ASAP7_75t_SL \i43/i47/i9  (.A(\i43/i47/n480 ),
    .B(\i43/i47/n497 ),
    .C(\i43/i47/n494 ),
    .D(\i43/i47/n456 ),
    .Y(\i43/i47/n505 ));
 NOR5xp2_ASAP7_75t_SL \i43/i47/i90  (.A(\i43/i47/n335 ),
    .B(\i43/i47/n338 ),
    .C(\i43/i47/n119 ),
    .D(\i43/i47/n152 ),
    .E(\i43/i47/n102 ),
    .Y(\i43/i47/n422 ));
 AOI221xp5_ASAP7_75t_SL \i43/i47/i91  (.A1(\i43/i47/n258 ),
    .A2(\i43/i47/n55 ),
    .B1(\i43/i47/n155 ),
    .B2(\i43/i47/n256 ),
    .C(\i43/i47/n211 ),
    .Y(\i43/i47/n421 ));
 NOR5xp2_ASAP7_75t_SL \i43/i47/i92  (.A(\i43/i47/n212 ),
    .B(\i43/i47/n270 ),
    .C(\i43/i47/n239 ),
    .D(\i43/i47/n218 ),
    .E(\i43/i47/n177 ),
    .Y(\i43/i47/n420 ));
 NOR5xp2_ASAP7_75t_SL \i43/i47/i93  (.A(\i43/i47/n314 ),
    .B(\i43/i47/n350 ),
    .C(\i43/i47/n340 ),
    .D(\i43/i47/n217 ),
    .E(\i43/i47/n223 ),
    .Y(\i43/i47/n419 ));
 AOI211xp5_ASAP7_75t_SL \i43/i47/i94  (.A1(\i43/i47/n0 ),
    .A2(\i43/i47/n38 ),
    .B(\i43/i47/n297 ),
    .C(\i43/i47/n289 ),
    .Y(\i43/i47/n418 ));
 NOR5xp2_ASAP7_75t_SL \i43/i47/i95  (.A(\i43/i47/n328 ),
    .B(\i43/i47/n274 ),
    .C(\i43/i47/n280 ),
    .D(\i43/i47/n124 ),
    .E(\i43/i47/n174 ),
    .Y(\i43/i47/n417 ));
 NOR2xp67_ASAP7_75t_SL \i43/i47/i96  (.A(\i43/i47/n402 ),
    .B(\i43/i47/n404 ),
    .Y(\i43/i47/n435 ));
 AO211x2_ASAP7_75t_SL \i43/i47/i97  (.A1(\i43/i47/n88 ),
    .A2(\i43/i47/n262 ),
    .B(\i43/i47/n234 ),
    .C(\i43/i47/n313 ),
    .Y(\i43/i47/n434 ));
 AOI21xp5_ASAP7_75t_SL \i43/i47/i98  (.A1(\i43/i47/n33 ),
    .A2(\i43/i47/n73 ),
    .B(\i43/i47/n511 ),
    .Y(\i43/i47/n433 ));
 INVx1_ASAP7_75t_SL \i43/i47/i99  (.A(\i43/i47/n412 ),
    .Y(\i43/i47/n413 ));
 INVxp67_ASAP7_75t_SL \i43/i470  (.A(net83),
    .Y(\i43/n162 ));
 INVxp67_ASAP7_75t_SL \i43/i471  (.A(net102),
    .Y(\i43/n161 ));
 INVxp67_ASAP7_75t_SL \i43/i472  (.A(net117),
    .Y(\i43/n160 ));
 INVxp67_ASAP7_75t_SL \i43/i473  (.A(net34),
    .Y(\i43/n159 ));
 INVxp67_ASAP7_75t_SL \i43/i474  (.A(net101),
    .Y(\i43/n158 ));
 INVxp67_ASAP7_75t_SL \i43/i475  (.A(net78),
    .Y(\i43/n157 ));
 INVxp67_ASAP7_75t_SL \i43/i476  (.A(net46),
    .Y(\i43/n156 ));
 INVxp67_ASAP7_75t_SL \i43/i477  (.A(net68),
    .Y(\i43/n155 ));
 INVxp67_ASAP7_75t_SL \i43/i478  (.A(net121),
    .Y(\i43/n154 ));
 INVxp67_ASAP7_75t_SL \i43/i479  (.A(net75),
    .Y(\i43/n153 ));
 NOR2x1_ASAP7_75t_SL \i43/i48/i0  (.A(\i43/i48/n479 ),
    .B(\i43/i48/n506 ),
    .Y(\i43/n0 [9]));
 AND3x1_ASAP7_75t_SL \i43/i48/i1  (.A(\i43/i48/n502 ),
    .B(\i43/i48/n504 ),
    .C(\i43/i48/n483 ),
    .Y(\i43/n0 [13]));
 NOR4xp75_ASAP7_75t_SL \i43/i48/i10  (.A(\i43/i48/n492 ),
    .B(\i43/i48/n496 ),
    .C(\i43/i48/n474 ),
    .D(\i43/i48/n489 ),
    .Y(\i43/n0 [10]));
 INVx1_ASAP7_75t_SL \i43/i48/i100  (.A(\i43/i48/n409 ),
    .Y(\i43/i48/n410 ));
 INVx1_ASAP7_75t_SL \i43/i48/i101  (.A(\i43/i48/n407 ),
    .Y(\i43/i48/n408 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i102  (.A(\i43/i48/n356 ),
    .B(\i43/i48/n351 ),
    .Y(\i43/i48/n406 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i103  (.A(\i43/i48/n325 ),
    .B(\i43/i48/n321 ),
    .Y(\i43/i48/n405 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i104  (.A(\i43/i48/n369 ),
    .B(\i43/i48/n324 ),
    .Y(\i43/i48/n404 ));
 NAND3xp33_ASAP7_75t_L \i43/i48/i105  (.A(\i43/i48/n267 ),
    .B(\i43/i48/n273 ),
    .C(\i43/i48/n354 ),
    .Y(\i43/i48/n403 ));
 NAND2xp5_ASAP7_75t_L \i43/i48/i106  (.A(\i43/i48/n337 ),
    .B(\i43/i48/n213 ),
    .Y(\i43/i48/n402 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i107  (.A(\i43/i48/n357 ),
    .B(\i43/i48/n331 ),
    .Y(\i43/i48/n401 ));
 NAND5xp2_ASAP7_75t_SL \i43/i48/i108  (.A(\i43/i48/n296 ),
    .B(\i43/i48/n120 ),
    .C(\i43/i48/n181 ),
    .D(\i43/i48/n123 ),
    .E(\i43/i48/n117 ),
    .Y(\i43/i48/n400 ));
 NOR4xp25_ASAP7_75t_SL \i43/i48/i109  (.A(\i43/i48/n279 ),
    .B(\i43/i48/n196 ),
    .C(\i43/i48/n131 ),
    .D(\i43/i48/n225 ),
    .Y(\i43/i48/n399 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i11  (.A(\i43/i48/n509 ),
    .B(\i43/i48/n491 ),
    .Y(\i43/i48/n504 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i110  (.A(\i43/i48/n347 ),
    .B(\i43/i48/n359 ),
    .Y(\i43/i48/n398 ));
 NAND2xp33_ASAP7_75t_SL \i43/i48/i111  (.A(\i43/i48/n320 ),
    .B(\i43/i48/n303 ),
    .Y(\i43/i48/n397 ));
 AOI221xp5_ASAP7_75t_SL \i43/i48/i112  (.A1(\i43/i48/n109 ),
    .A2(\i43/i48/n95 ),
    .B1(\i43/i48/n115 ),
    .B2(\i43/i48/n47 ),
    .C(\i43/i48/n215 ),
    .Y(\i43/i48/n416 ));
 NAND5xp2_ASAP7_75t_SL \i43/i48/i113  (.A(\i43/i48/n277 ),
    .B(\i43/i48/n205 ),
    .C(\i43/i48/n210 ),
    .D(\i43/i48/n181 ),
    .E(\i43/i48/n122 ),
    .Y(\i43/i48/n396 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i114  (.A(\i43/i48/n293 ),
    .B(\i43/i48/n369 ),
    .Y(\i43/i48/n395 ));
 OAI221xp5_ASAP7_75t_SL \i43/i48/i115  (.A1(\i43/i48/n156 ),
    .A2(\i43/i48/n54 ),
    .B1(\i43/i48/n157 ),
    .B2(\i43/i48/n39 ),
    .C(\i43/i48/n336 ),
    .Y(\i43/i48/n394 ));
 NOR2xp33_ASAP7_75t_L \i43/i48/i116  (.A(\i43/i48/n290 ),
    .B(\i43/i48/n356 ),
    .Y(\i43/i48/n415 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i117  (.A(\i43/i48/n287 ),
    .B(\i43/i48/n319 ),
    .Y(\i43/i48/n414 ));
 NOR3xp33_ASAP7_75t_SL \i43/i48/i118  (.A(\i43/i48/n217 ),
    .B(\i43/i48/n226 ),
    .C(\i43/i48/n195 ),
    .Y(\i43/i48/n412 ));
 NAND3xp33_ASAP7_75t_SL \i43/i48/i119  (.A(\i43/i48/n332 ),
    .B(\i43/i48/n283 ),
    .C(\i43/i48/n238 ),
    .Y(\i43/i48/n411 ));
 NAND3xp33_ASAP7_75t_SL \i43/i48/i12  (.A(\i43/i48/n477 ),
    .B(\i43/i48/n482 ),
    .C(\i43/i48/n416 ),
    .Y(\i43/i48/n503 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i120  (.A(\i43/i48/n214 ),
    .B(\i43/i48/n298 ),
    .Y(\i43/i48/n409 ));
 NOR3xp33_ASAP7_75t_SL \i43/i48/i121  (.A(\i43/i48/n286 ),
    .B(\i43/i48/n231 ),
    .C(\i43/i48/n270 ),
    .Y(\i43/i48/n407 ));
 INVx1_ASAP7_75t_SL \i43/i48/i122  (.A(\i43/i48/n514 ),
    .Y(\i43/i48/n387 ));
 OAI21xp33_ASAP7_75t_SL \i43/i48/i123  (.A1(\i43/i48/n76 ),
    .A2(\i43/i48/n45 ),
    .B(\i43/i48/n367 ),
    .Y(\i43/i48/n386 ));
 NOR3xp33_ASAP7_75t_SL \i43/i48/i124  (.A(\i43/i48/n327 ),
    .B(\i43/i48/n191 ),
    .C(\i43/i48/n231 ),
    .Y(\i43/i48/n385 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i125  (.A1(\i43/i48/n87 ),
    .A2(\i43/i48/n50 ),
    .B(\i43/i48/n354 ),
    .Y(\i43/i48/n393 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i126  (.A1(\i43/i48/n41 ),
    .A2(\i43/i48/n268 ),
    .B(\i43/i48/n263 ),
    .Y(\i43/i48/n384 ));
 NAND4xp25_ASAP7_75t_SL \i43/i48/i127  (.A(\i43/i48/n244 ),
    .B(\i43/i48/n145 ),
    .C(\i43/i48/n96 ),
    .D(\i43/i48/n99 ),
    .Y(\i43/i48/n383 ));
 NAND5xp2_ASAP7_75t_SL \i43/i48/i128  (.A(\i43/i48/n208 ),
    .B(\i43/i48/n120 ),
    .C(\i43/i48/n164 ),
    .D(\i43/i48/n184 ),
    .E(\i43/i48/n140 ),
    .Y(\i43/i48/n382 ));
 AOI211xp5_ASAP7_75t_SL \i43/i48/i129  (.A1(\i43/i48/n41 ),
    .A2(\i43/i48/n62 ),
    .B(\i43/i48/n282 ),
    .C(\i43/i48/n281 ),
    .Y(\i43/i48/n381 ));
 NOR3xp33_ASAP7_75t_SL \i43/i48/i13  (.A(\i43/i48/n508 ),
    .B(\i43/i48/n478 ),
    .C(\i43/i48/n455 ),
    .Y(\i43/i48/n502 ));
 NOR3xp33_ASAP7_75t_SL \i43/i48/i130  (.A(\i43/i48/n292 ),
    .B(\i43/i48/n206 ),
    .C(\i43/i48/n221 ),
    .Y(\i43/i48/n380 ));
 NOR2xp33_ASAP7_75t_L \i43/i48/i131  (.A(\i43/i48/n334 ),
    .B(\i43/i48/n315 ),
    .Y(\i43/i48/n379 ));
 OAI221xp5_ASAP7_75t_SL \i43/i48/i132  (.A1(\i43/i48/n269 ),
    .A2(\i43/i48/n75 ),
    .B1(\i43/i48/n173 ),
    .B2(\i43/i48/n72 ),
    .C(\i43/i48/n89 ),
    .Y(\i43/i48/n378 ));
 NAND5xp2_ASAP7_75t_SL \i43/i48/i133  (.A(\i43/i48/n246 ),
    .B(\i43/i48/n175 ),
    .C(\i43/i48/n105 ),
    .D(\i43/i48/n113 ),
    .E(\i43/i48/n144 ),
    .Y(\i43/i48/n377 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i134  (.A1(\i43/i48/n45 ),
    .A2(\i43/i48/n40 ),
    .B(\i43/i48/n357 ),
    .Y(\i43/i48/n376 ));
 NOR4xp25_ASAP7_75t_SL \i43/i48/i135  (.A(\i43/i48/n333 ),
    .B(\i43/i48/n266 ),
    .C(\i43/i48/n97 ),
    .D(\i43/i48/n98 ),
    .Y(\i43/i48/n375 ));
 OAI211xp5_ASAP7_75t_SL \i43/i48/i136  (.A1(\i43/i48/n40 ),
    .A2(\i43/i48/n259 ),
    .B(\i43/i48/n179 ),
    .C(\i43/i48/n167 ),
    .Y(\i43/i48/n374 ));
 NAND5xp2_ASAP7_75t_SL \i43/i48/i137  (.A(\i43/i48/n257 ),
    .B(\i43/i48/n242 ),
    .C(\i43/i48/n118 ),
    .D(\i43/i48/n180 ),
    .E(\i43/i48/n185 ),
    .Y(\i43/i48/n373 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i138  (.A(\i43/i48/n330 ),
    .B(\i43/i48/n301 ),
    .Y(\i43/i48/n372 ));
 OAI221xp5_ASAP7_75t_SL \i43/i48/i139  (.A1(\i43/i48/n260 ),
    .A2(\i43/i48/n54 ),
    .B1(\i43/i48/n52 ),
    .B2(\i43/i48/n87 ),
    .C(\i43/i48/n222 ),
    .Y(\i43/i48/n371 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i14  (.A(\i43/i48/n493 ),
    .B(\i43/i48/n481 ),
    .Y(\i43/i48/n501 ));
 NOR3xp33_ASAP7_75t_SL \i43/i48/i140  (.A(\i43/i48/n307 ),
    .B(\i43/i48/n274 ),
    .C(\i43/i48/n272 ),
    .Y(\i43/i48/n392 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i141  (.A(\i43/i48/n240 ),
    .B(\i43/i48/n358 ),
    .Y(\i43/i48/n391 ));
 OA211x2_ASAP7_75t_SL \i43/i48/i142  (.A1(\i43/i48/n92 ),
    .A2(\i43/i48/n54 ),
    .B(\i43/i48/n366 ),
    .C(\i43/i48/n146 ),
    .Y(\i43/i48/n390 ));
 NOR2xp33_ASAP7_75t_L \i43/i48/i143  (.A(\i43/i48/n190 ),
    .B(\i43/i48/n316 ),
    .Y(\i43/i48/n389 ));
 NOR2xp33_ASAP7_75t_L \i43/i48/i144  (.A(\i43/i48/n200 ),
    .B(\i43/i48/n362 ),
    .Y(\i43/i48/n388 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i145  (.A(\i43/i48/n364 ),
    .Y(\i43/i48/n365 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i146  (.A(\i43/i48/n362 ),
    .Y(\i43/i48/n363 ));
 INVx1_ASAP7_75t_SL \i43/i48/i147  (.A(\i43/i48/n360 ),
    .Y(\i43/i48/n361 ));
 INVx1_ASAP7_75t_SL \i43/i48/i148  (.A(\i43/i48/n358 ),
    .Y(\i43/i48/n359 ));
 INVx1_ASAP7_75t_SL \i43/i48/i149  (.A(\i43/i48/n512 ),
    .Y(\i43/i48/n352 ));
 NAND3xp33_ASAP7_75t_SL \i43/i48/i15  (.A(\i43/i48/n466 ),
    .B(\i43/i48/n476 ),
    .C(\i43/i48/n454 ),
    .Y(\i43/i48/n500 ));
 NAND2xp33_ASAP7_75t_L \i43/i48/i150  (.A(\i43/i48/n214 ),
    .B(\i43/i48/n271 ),
    .Y(\i43/i48/n351 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i151  (.A(\i43/i48/n130 ),
    .B(\i43/i48/n220 ),
    .Y(\i43/i48/n350 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i152  (.A(\i43/i48/n192 ),
    .B(\i43/i48/n212 ),
    .Y(\i43/i48/n349 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i48/i153  (.A1(\i43/i48/n34 ),
    .A2(\i43/i48/n65 ),
    .B(\i43/i48/n33 ),
    .C(\i43/i48/n227 ),
    .Y(\i43/i48/n348 ));
 OAI31xp33_ASAP7_75t_SL \i43/i48/i154  (.A1(\i43/i48/n65 ),
    .A2(\i43/i48/n41 ),
    .A3(\i43/i48/n55 ),
    .B(\i43/i48/n79 ),
    .Y(\i43/i48/n347 ));
 NAND3xp33_ASAP7_75t_SL \i43/i48/i155  (.A(\i43/i48/n213 ),
    .B(\i43/i48/n183 ),
    .C(\i43/i48/n128 ),
    .Y(\i43/i48/n346 ));
 AOI21xp5_ASAP7_75t_SL \i43/i48/i156  (.A1(\i43/i48/n38 ),
    .A2(\i43/i48/n74 ),
    .B(\i43/i48/n1 ),
    .Y(\i43/i48/n345 ));
 AOI211xp5_ASAP7_75t_SL \i43/i48/i157  (.A1(\i43/i48/n57 ),
    .A2(\i43/i48/n71 ),
    .B(\i43/i48/n182 ),
    .C(\i43/i48/n121 ),
    .Y(\i43/i48/n370 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i158  (.A1(\i43/i48/n94 ),
    .A2(\i43/i48/n58 ),
    .B(\i43/i48/n216 ),
    .Y(\i43/i48/n344 ));
 OAI31xp33_ASAP7_75t_SL \i43/i48/i159  (.A1(\i43/i48/n47 ),
    .A2(\i43/i48/n95 ),
    .A3(\i43/i48/n51 ),
    .B(\i43/i48/n69 ),
    .Y(\i43/i48/n343 ));
 NOR2xp33_ASAP7_75t_L \i43/i48/i16  (.A(\i43/i48/n465 ),
    .B(\i43/i48/n461 ),
    .Y(\i43/i48/n497 ));
 AO21x1_ASAP7_75t_SL \i43/i48/i160  (.A1(\i43/i48/n67 ),
    .A2(\i43/i48/n150 ),
    .B(\i43/i48/n280 ),
    .Y(\i43/i48/n342 ));
 AO21x1_ASAP7_75t_SL \i43/i48/i161  (.A1(\i43/i48/n148 ),
    .A2(\i43/i48/n173 ),
    .B(\i43/i48/n76 ),
    .Y(\i43/i48/n341 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i43/i48/i162  (.A1(\i43/i48/n70 ),
    .A2(\i43/i48/n78 ),
    .B(\i43/i48/n52 ),
    .C(\i43/i48/n197 ),
    .Y(\i43/i48/n340 ));
 AOI21xp5_ASAP7_75t_SL \i43/i48/i163  (.A1(\i43/i48/n44 ),
    .A2(\i43/i48/n67 ),
    .B(\i43/i48/n219 ),
    .Y(\i43/i48/n339 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i43/i48/i164  (.A1(\i43/i48/n42 ),
    .A2(\i43/i48/n35 ),
    .B(\i43/i48/n87 ),
    .C(\i43/i48/n117 ),
    .Y(\i43/i48/n338 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i165  (.A(\i43/i48/n249 ),
    .B(\i43/i48/n236 ),
    .Y(\i43/i48/n337 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i48/i166  (.A1(\i43/i48/n77 ),
    .A2(\i43/i48/n51 ),
    .B(\i43/i48/n33 ),
    .C(\i43/i48/n132 ),
    .Y(\i43/i48/n336 ));
 NAND3xp33_ASAP7_75t_SL \i43/i48/i167  (.A(\i43/i48/n232 ),
    .B(\i43/i48/n172 ),
    .C(\i43/i48/n137 ),
    .Y(\i43/i48/n335 ));
 OAI221xp5_ASAP7_75t_SL \i43/i48/i168  (.A1(\i43/i48/n75 ),
    .A2(\i43/i48/n56 ),
    .B1(\i43/i48/n49 ),
    .B2(\i43/i48/n68 ),
    .C(\i43/i48/n134 ),
    .Y(\i43/i48/n334 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i169  (.A1(\i43/i48/n78 ),
    .A2(\i43/i48/n136 ),
    .B(\i43/i48/n237 ),
    .Y(\i43/i48/n333 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i17  (.A(\i43/i48/n468 ),
    .B(\i43/i48/n476 ),
    .Y(\i43/i48/n496 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i170  (.A(\i43/i48/n233 ),
    .B(\i43/i48/n209 ),
    .Y(\i43/i48/n332 ));
 AOI221xp5_ASAP7_75t_SL \i43/i48/i171  (.A1(\i43/i48/n34 ),
    .A2(\i43/i48/n79 ),
    .B1(\i43/i48/n67 ),
    .B2(\i43/i48/n83 ),
    .C(\i43/i48/n236 ),
    .Y(\i43/i48/n331 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i172  (.A1(\i43/i48/n59 ),
    .A2(\i43/i48/n154 ),
    .B(\i43/i48/n77 ),
    .Y(\i43/i48/n330 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i48/i173  (.A1(\i43/i48/n62 ),
    .A2(\i43/i48/n44 ),
    .B(\i43/i48/n57 ),
    .C(\i43/i48/n125 ),
    .Y(\i43/i48/n329 ));
 OAI221xp5_ASAP7_75t_SL \i43/i48/i174  (.A1(\i43/i48/n46 ),
    .A2(\i43/i48/n87 ),
    .B1(\i43/i48/n52 ),
    .B2(\i43/i48/n80 ),
    .C(\i43/i48/n162 ),
    .Y(\i43/i48/n328 ));
 AOI21xp5_ASAP7_75t_SL \i43/i48/i175  (.A1(\i43/i48/n95 ),
    .A2(\i43/i48/n62 ),
    .B(\i43/i48/n1 ),
    .Y(\i43/i48/n369 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i176  (.A(\i43/i48/n219 ),
    .B(\i43/i48/n251 ),
    .Y(\i43/i48/n368 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i177  (.A(\i43/i48/n253 ),
    .B(\i43/i48/n0 ),
    .Y(\i43/i48/n367 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i178  (.A(\i43/i48/n225 ),
    .B(\i43/i48/n194 ),
    .Y(\i43/i48/n366 ));
 OAI211xp5_ASAP7_75t_SL \i43/i48/i179  (.A1(\i43/i48/n63 ),
    .A2(\i43/i48/n46 ),
    .B(\i43/i48/n176 ),
    .C(\i43/i48/n186 ),
    .Y(\i43/i48/n364 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i18  (.A(\i43/i48/n473 ),
    .B(\i43/i48/n464 ),
    .Y(\i43/i48/n495 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i180  (.A(\i43/i48/n120 ),
    .B(\i43/i48/n245 ),
    .Y(\i43/i48/n362 ));
 AOI222xp33_ASAP7_75t_SL \i43/i48/i181  (.A1(\i43/i48/n85 ),
    .A2(\i43/i48/n41 ),
    .B1(\i43/i48/n59 ),
    .B2(\i43/i48/n38 ),
    .C1(\i43/i48/n69 ),
    .C2(\i43/i48/n47 ),
    .Y(\i43/i48/n360 ));
 OAI221xp5_ASAP7_75t_SL \i43/i48/i182  (.A1(\i43/i48/n45 ),
    .A2(\i43/i48/n35 ),
    .B1(\i43/i48/n37 ),
    .B2(\i43/i48/n52 ),
    .C(\i43/i48/n179 ),
    .Y(\i43/i48/n358 ));
 AOI222xp33_ASAP7_75t_SL \i43/i48/i183  (.A1(\i43/i48/n34 ),
    .A2(\i43/i48/n90 ),
    .B1(\i43/i48/n33 ),
    .B2(\i43/i48/n67 ),
    .C1(\i43/i48/n83 ),
    .C2(\i43/i48/n73 ),
    .Y(\i43/i48/n357 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i184  (.A1(\i43/i48/n39 ),
    .A2(\i43/i48/n91 ),
    .B(\i43/i48/n237 ),
    .Y(\i43/i48/n356 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i185  (.A(\i43/i48/n204 ),
    .B(\i43/i48/n227 ),
    .Y(\i43/i48/n355 ));
 NOR2xp67_ASAP7_75t_SL \i43/i48/i186  (.A(\i43/i48/n255 ),
    .B(\i43/i48/n279 ),
    .Y(\i43/i48/n354 ));
 NOR2x1_ASAP7_75t_SL \i43/i48/i187  (.A(\i43/i48/n141 ),
    .B(\i43/i48/n278 ),
    .Y(\i43/i48/n353 ));
 INVxp33_ASAP7_75t_SL \i43/i48/i188  (.A(\i43/i48/n324 ),
    .Y(\i43/i48/n325 ));
 INVx1_ASAP7_75t_SL \i43/i48/i189  (.A(\i43/i48/n321 ),
    .Y(\i43/i48/n322 ));
 NOR4xp25_ASAP7_75t_SL \i43/i48/i19  (.A(\i43/i48/n429 ),
    .B(\i43/i48/n395 ),
    .C(\i43/i48/n372 ),
    .D(\i43/i48/n371 ),
    .Y(\i43/i48/n494 ));
 INVx1_ASAP7_75t_SL \i43/i48/i190  (.A(\i43/i48/n316 ),
    .Y(\i43/i48/n317 ));
 OAI211xp5_ASAP7_75t_SL \i43/i48/i191  (.A1(\i43/i48/n40 ),
    .A2(\i43/i48/n70 ),
    .B(\i43/i48/n188 ),
    .C(\i43/i48/n187 ),
    .Y(\i43/i48/n315 ));
 AO21x1_ASAP7_75t_SL \i43/i48/i192  (.A1(\i43/i48/n67 ),
    .A2(\i43/i48/n0 ),
    .B(\i43/i48/n224 ),
    .Y(\i43/i48/n314 ));
 OAI221xp5_ASAP7_75t_SL \i43/i48/i193  (.A1(\i43/i48/n72 ),
    .A2(\i43/i48/n70 ),
    .B1(\i43/i48/n42 ),
    .B2(\i43/i48/n63 ),
    .C(\i43/i48/n118 ),
    .Y(\i43/i48/n313 ));
 OA211x2_ASAP7_75t_SL \i43/i48/i194  (.A1(\i43/i48/n37 ),
    .A2(\i43/i48/n136 ),
    .B(\i43/i48/n100 ),
    .C(\i43/i48/n159 ),
    .Y(\i43/i48/n312 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i48/i195  (.A1(\i43/i48/n47 ),
    .A2(\i43/i48/n34 ),
    .B(\i43/i48/n85 ),
    .C(\i43/i48/n241 ),
    .Y(\i43/i48/n311 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i196  (.A(\i43/i48/n265 ),
    .B(\i43/i48/n266 ),
    .Y(\i43/i48/n310 ));
 OAI31xp33_ASAP7_75t_SL \i43/i48/i197  (.A1(\i43/i48/n57 ),
    .A2(\i43/i48/n53 ),
    .A3(\i43/i48/n88 ),
    .B(\i43/i48/n62 ),
    .Y(\i43/i48/n309 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i198  (.A1(\i43/i48/n51 ),
    .A2(\i43/i48/n166 ),
    .B(\i43/i48/n71 ),
    .Y(\i43/i48/n308 ));
 OAI211xp5_ASAP7_75t_SL \i43/i48/i199  (.A1(\i43/i48/n52 ),
    .A2(\i43/i48/n91 ),
    .B(\i43/i48/n138 ),
    .C(\i43/i48/n139 ),
    .Y(\i43/i48/n307 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i2  (.A(\i43/i48/n507 ),
    .B(\i43/i48/n503 ),
    .Y(\i43/n0 [14]));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i20  (.A(\i43/i48/n452 ),
    .B(\i43/i48/n459 ),
    .Y(\i43/i48/n493 ));
 OAI221xp5_ASAP7_75t_SL \i43/i48/i200  (.A1(\i43/i48/n94 ),
    .A2(\i43/i48/n87 ),
    .B1(\i43/i48/n78 ),
    .B2(\i43/i48/n54 ),
    .C(\i43/i48/n137 ),
    .Y(\i43/i48/n306 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i201  (.A1(\i43/i48/n56 ),
    .A2(\i43/i48/n156 ),
    .B1(\i43/i48/n63 ),
    .B2(\i43/i48/n72 ),
    .Y(\i43/i48/n305 ));
 OAI211xp5_ASAP7_75t_SL \i43/i48/i202  (.A1(\i43/i48/n82 ),
    .A2(\i43/i48/n72 ),
    .B(\i43/i48/n264 ),
    .C(\i43/i48/n178 ),
    .Y(\i43/i48/n304 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i48/i203  (.A1(\i43/i48/n51 ),
    .A2(\i43/i48/n53 ),
    .B(\i43/i48/n85 ),
    .C(\i43/i48/n203 ),
    .Y(\i43/i48/n303 ));
 AOI221xp5_ASAP7_75t_SL \i43/i48/i204  (.A1(\i43/i48/n44 ),
    .A2(\i43/i48/n38 ),
    .B1(\i43/i48/n104 ),
    .B2(\i43/i48/n71 ),
    .C(\i43/i48/n161 ),
    .Y(\i43/i48/n302 ));
 NOR3xp33_ASAP7_75t_SL \i43/i48/i205  (.A(\i43/i48/n250 ),
    .B(\i43/i48/n170 ),
    .C(\i43/i48/n101 ),
    .Y(\i43/i48/n301 ));
 AOI21xp5_ASAP7_75t_SL \i43/i48/i206  (.A1(\i43/i48/n150 ),
    .A2(\i43/i48/n73 ),
    .B(\i43/i48/n261 ),
    .Y(\i43/i48/n300 ));
 OAI211xp5_ASAP7_75t_SL \i43/i48/i207  (.A1(\i43/i48/n89 ),
    .A2(\i43/i48/n157 ),
    .B(\i43/i48/n126 ),
    .C(\i43/i48/n135 ),
    .Y(\i43/i48/n299 ));
 AOI222xp33_ASAP7_75t_SL \i43/i48/i208  (.A1(\i43/i48/n112 ),
    .A2(\i43/i48/n67 ),
    .B1(\i43/i48/n65 ),
    .B2(\i43/i48/n79 ),
    .C1(\i43/i48/n59 ),
    .C2(\i43/i48/n48 ),
    .Y(\i43/i48/n298 ));
 NAND4xp25_ASAP7_75t_SL \i43/i48/i209  (.A(\i43/i48/n133 ),
    .B(\i43/i48/n164 ),
    .C(\i43/i48/n171 ),
    .D(\i43/i48/n111 ),
    .Y(\i43/i48/n297 ));
 NAND2x1_ASAP7_75t_SL \i43/i48/i21  (.A(\i43/i48/n458 ),
    .B(\i43/i48/n469 ),
    .Y(\i43/i48/n492 ));
 AOI221xp5_ASAP7_75t_SL \i43/i48/i210  (.A1(\i43/i48/n48 ),
    .A2(\i43/i48/n81 ),
    .B1(\i43/i48/n41 ),
    .B2(\i43/i48/n85 ),
    .C(\i43/i48/n207 ),
    .Y(\i43/i48/n296 ));
 AOI222xp33_ASAP7_75t_SL \i43/i48/i211  (.A1(\i43/i48/n67 ),
    .A2(\i43/i48/n60 ),
    .B1(\i43/i48/n88 ),
    .B2(\i43/i48/n85 ),
    .C1(\i43/i48/n95 ),
    .C2(\i43/i48/n71 ),
    .Y(\i43/i48/n295 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i48/i212  (.A1(\i43/i48/n44 ),
    .A2(\i43/i48/n36 ),
    .B(\i43/i48/n48 ),
    .C(\i43/i48/n215 ),
    .Y(\i43/i48/n294 ));
 AOI22xp33_ASAP7_75t_SL \i43/i48/i213  (.A1(\i43/i48/n65 ),
    .A2(\i43/i48/n0 ),
    .B1(\i43/i48/n33 ),
    .B2(\i43/i48/n106 ),
    .Y(\i43/i48/n293 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i214  (.A1(\i43/i48/n75 ),
    .A2(\i43/i48/n103 ),
    .B1(\i43/i48/n46 ),
    .B2(\i43/i48/n37 ),
    .Y(\i43/i48/n292 ));
 AOI211xp5_ASAP7_75t_SL \i43/i48/i215  (.A1(\i43/i48/n67 ),
    .A2(\i43/i48/n79 ),
    .B(\i43/i48/n254 ),
    .C(\i43/i48/n170 ),
    .Y(\i43/i48/n291 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i216  (.A1(\i43/i48/n87 ),
    .A2(\i43/i48/n114 ),
    .B1(\i43/i48/n76 ),
    .B2(\i43/i48/n37 ),
    .Y(\i43/i48/n290 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i43/i48/i217  (.A1(\i43/i48/n42 ),
    .A2(\i43/i48/n49 ),
    .B(\i43/i48/n80 ),
    .C(\i43/i48/n252 ),
    .Y(\i43/i48/n289 ));
 AOI22xp5_ASAP7_75t_SL \i43/i48/i218  (.A1(\i43/i48/n83 ),
    .A2(\i43/i48/n143 ),
    .B1(\i43/i48/n71 ),
    .B2(\i43/i48/n38 ),
    .Y(\i43/i48/n288 ));
 AOI222xp33_ASAP7_75t_SL \i43/i48/i219  (.A1(\i43/i48/n79 ),
    .A2(\i43/i48/n48 ),
    .B1(\i43/i48/n69 ),
    .B2(\i43/i48/n38 ),
    .C1(\i43/i48/n74 ),
    .C2(\i43/i48/n67 ),
    .Y(\i43/i48/n287 ));
 NAND4xp25_ASAP7_75t_SL \i43/i48/i22  (.A(\i43/i48/n423 ),
    .B(\i43/i48/n427 ),
    .C(\i43/i48/n388 ),
    .D(\i43/i48/n443 ),
    .Y(\i43/i48/n491 ));
 OAI221xp5_ASAP7_75t_SL \i43/i48/i220  (.A1(\i43/i48/n35 ),
    .A2(\i43/i48/n80 ),
    .B1(\i43/i48/n68 ),
    .B2(\i43/i48/n76 ),
    .C(\i43/i48/n116 ),
    .Y(\i43/i48/n286 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i221  (.A(\i43/i48/n281 ),
    .B(\i43/i48/n282 ),
    .Y(\i43/i48/n285 ));
 AO21x1_ASAP7_75t_L \i43/i48/i222  (.A1(\i43/i48/n41 ),
    .A2(\i43/i48/n163 ),
    .B(\i43/i48/n198 ),
    .Y(\i43/i48/n327 ));
 AOI21xp5_ASAP7_75t_SL \i43/i48/i223  (.A1(\i43/i48/n154 ),
    .A2(\i43/i48/n88 ),
    .B(\i43/i48/n202 ),
    .Y(\i43/i48/n326 ));
 OA211x2_ASAP7_75t_SL \i43/i48/i224  (.A1(\i43/i48/n54 ),
    .A2(\i43/i48/n142 ),
    .B(\i43/i48/n128 ),
    .C(\i43/i48/n162 ),
    .Y(\i43/i48/n324 ));
 AOI22xp5_ASAP7_75t_SL \i43/i48/i225  (.A1(\i43/i48/n41 ),
    .A2(\i43/i48/n147 ),
    .B1(\i43/i48/n60 ),
    .B2(\i43/i48/n77 ),
    .Y(\i43/i48/n323 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i226  (.A(\i43/i48/n283 ),
    .B(\i43/i48/n238 ),
    .Y(\i43/i48/n284 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i227  (.A1(\i43/i48/n80 ),
    .A2(\i43/i48/n165 ),
    .B1(\i43/i48/n84 ),
    .B2(\i43/i48/n64 ),
    .Y(\i43/i48/n321 ));
 AOI21xp5_ASAP7_75t_SL \i43/i48/i228  (.A1(\i43/i48/n48 ),
    .A2(\i43/i48/n71 ),
    .B(\i43/i48/n218 ),
    .Y(\i43/i48/n320 ));
 AOI222xp33_ASAP7_75t_SL \i43/i48/i229  (.A1(\i43/i48/n43 ),
    .A2(\i43/i48/n59 ),
    .B1(\i43/i48/n73 ),
    .B2(\i43/i48/n85 ),
    .C1(\i43/i48/n34 ),
    .C2(\i43/i48/n71 ),
    .Y(\i43/i48/n319 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i23  (.A(\i43/i48/n470 ),
    .B(\i43/i48/n474 ),
    .Y(\i43/i48/n490 ));
 O2A1O1Ixp33_ASAP7_75t_L \i43/i48/i230  (.A1(\i43/i48/n41 ),
    .A2(\i43/i48/n48 ),
    .B(\i43/i48/n83 ),
    .C(\i43/i48/n224 ),
    .Y(\i43/i48/n318 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i231  (.A(\i43/i48/n108 ),
    .B(\i43/i48/n273 ),
    .Y(\i43/i48/n316 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i232  (.A(\i43/i48/n275 ),
    .Y(\i43/i48/n276 ));
 INVx1_ASAP7_75t_SL \i43/i48/i233  (.A(\i43/i48/n271 ),
    .Y(\i43/i48/n272 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i234  (.A(\i43/i48/n268 ),
    .Y(\i43/i48/n269 ));
 OAI21xp33_ASAP7_75t_SL \i43/i48/i235  (.A1(\i43/i48/n75 ),
    .A2(\i43/i48/n52 ),
    .B(\i43/i48/n123 ),
    .Y(\i43/i48/n265 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i236  (.A(\i43/i48/n125 ),
    .B(\i43/i48/n152 ),
    .Y(\i43/i48/n264 ));
 NAND2xp33_ASAP7_75t_SL \i43/i48/i237  (.A(\i43/i48/n82 ),
    .B(\i43/i48/n127 ),
    .Y(\i43/i48/n263 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i238  (.A(\i43/i48/n75 ),
    .B(\i43/i48/n157 ),
    .Y(\i43/i48/n262 ));
 NAND2xp33_ASAP7_75t_SL \i43/i48/i239  (.A(\i43/i48/n184 ),
    .B(\i43/i48/n126 ),
    .Y(\i43/i48/n261 ));
 NOR2x1_ASAP7_75t_SL \i43/i48/i24  (.A(\i43/i48/n445 ),
    .B(\i43/i48/n465 ),
    .Y(\i43/i48/n499 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i240  (.A(\i43/i48/n60 ),
    .B(\i43/i48/n147 ),
    .Y(\i43/i48/n260 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i241  (.A(\i43/i48/n55 ),
    .B(\i43/i48/n147 ),
    .Y(\i43/i48/n283 ));
 NOR3xp33_ASAP7_75t_SL \i43/i48/i242  (.A(\i43/i48/n71 ),
    .B(\i43/i48/n33 ),
    .C(\i43/i48/n81 ),
    .Y(\i43/i48/n259 ));
 NAND2xp33_ASAP7_75t_L \i43/i48/i243  (.A(\i43/i48/n149 ),
    .B(\i43/i48/n32 ),
    .Y(\i43/i48/n258 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i244  (.A1(\i43/i48/n79 ),
    .A2(\i43/i48/n33 ),
    .B(\i43/i48/n43 ),
    .Y(\i43/i48/n257 ));
 NAND2xp33_ASAP7_75t_SL \i43/i48/i245  (.A(\i43/i48/n42 ),
    .B(\i43/i48/n134 ),
    .Y(\i43/i48/n256 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i246  (.A1(\i43/i48/n87 ),
    .A2(\i43/i48/n64 ),
    .B(\i43/i48/n172 ),
    .Y(\i43/i48/n255 ));
 OAI21xp33_ASAP7_75t_SL \i43/i48/i247  (.A1(\i43/i48/n35 ),
    .A2(\i43/i48/n87 ),
    .B(\i43/i48/n159 ),
    .Y(\i43/i48/n254 ));
 OAI21xp33_ASAP7_75t_SL \i43/i48/i248  (.A1(\i43/i48/n84 ),
    .A2(\i43/i48/n42 ),
    .B(\i43/i48/n52 ),
    .Y(\i43/i48/n253 ));
 OAI21xp33_ASAP7_75t_SL \i43/i48/i249  (.A1(\i43/i48/n95 ),
    .A2(\i43/i48/n53 ),
    .B(\i43/i48/n163 ),
    .Y(\i43/i48/n252 ));
 NOR3xp33_ASAP7_75t_SL \i43/i48/i25  (.A(\i43/i48/n447 ),
    .B(\i43/i48/n434 ),
    .C(\i43/i48/n393 ),
    .Y(\i43/i48/n498 ));
 OAI21xp33_ASAP7_75t_SL \i43/i48/i250  (.A1(\i43/i48/n66 ),
    .A2(\i43/i48/n80 ),
    .B(\i43/i48/n158 ),
    .Y(\i43/i48/n251 ));
 AOI21xp33_ASAP7_75t_SL \i43/i48/i251  (.A1(\i43/i48/n91 ),
    .A2(\i43/i48/n87 ),
    .B(\i43/i48/n49 ),
    .Y(\i43/i48/n250 ));
 OAI21xp33_ASAP7_75t_SL \i43/i48/i252  (.A1(\i43/i48/n58 ),
    .A2(\i43/i48/n35 ),
    .B(\i43/i48/n180 ),
    .Y(\i43/i48/n249 ));
 OAI21xp33_ASAP7_75t_SL \i43/i48/i253  (.A1(\i43/i48/n82 ),
    .A2(\i43/i48/n35 ),
    .B(\i43/i48/n158 ),
    .Y(\i43/i48/n248 ));
 AOI21xp5_ASAP7_75t_SL \i43/i48/i254  (.A1(\i43/i48/n64 ),
    .A2(\i43/i48/n42 ),
    .B(\i43/i48/n91 ),
    .Y(\i43/i48/n282 ));
 AOI21xp5_ASAP7_75t_SL \i43/i48/i255  (.A1(\i43/i48/n83 ),
    .A2(\i43/i48/n65 ),
    .B(\i43/i48/n129 ),
    .Y(\i43/i48/n247 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i256  (.A1(\i43/i48/n74 ),
    .A2(\i43/i48/n86 ),
    .B(\i43/i48/n55 ),
    .Y(\i43/i48/n246 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i257  (.A1(\i43/i48/n77 ),
    .A2(\i43/i48/n34 ),
    .B(\i43/i48/n79 ),
    .Y(\i43/i48/n245 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i258  (.A1(\i43/i48/n66 ),
    .A2(\i43/i48/n84 ),
    .B(\i43/i48/n178 ),
    .Y(\i43/i48/n281 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i259  (.A1(\i43/i48/n81 ),
    .A2(\i43/i48/n62 ),
    .B(\i43/i48/n65 ),
    .Y(\i43/i48/n244 ));
 NAND3xp33_ASAP7_75t_SL \i43/i48/i26  (.A(\i43/i48/n438 ),
    .B(\i43/i48/n440 ),
    .C(\i43/i48/n439 ),
    .Y(\i43/i48/n489 ));
 NAND3xp33_ASAP7_75t_L \i43/i48/i260  (.A(\i43/i48/n37 ),
    .B(\i43/i48/n87 ),
    .C(\i43/i48/n32 ),
    .Y(\i43/i48/n243 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i261  (.A1(\i43/i48/n90 ),
    .A2(\i43/i48/n69 ),
    .B(\i43/i48/n65 ),
    .Y(\i43/i48/n242 ));
 AOI21xp33_ASAP7_75t_SL \i43/i48/i262  (.A1(\i43/i48/n66 ),
    .A2(\i43/i48/n56 ),
    .B(\i43/i48/n75 ),
    .Y(\i43/i48/n241 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i263  (.A1(\i43/i48/n91 ),
    .A2(\i43/i48/n72 ),
    .B(\i43/i48/n185 ),
    .Y(\i43/i48/n240 ));
 OAI21xp33_ASAP7_75t_SL \i43/i48/i264  (.A1(\i43/i48/n80 ),
    .A2(\i43/i48/n54 ),
    .B(\i43/i48/n160 ),
    .Y(\i43/i48/n239 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i265  (.A1(\i43/i48/n39 ),
    .A2(\i43/i48/n82 ),
    .B(\i43/i48/n133 ),
    .Y(\i43/i48/n280 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i266  (.A1(\i43/i48/n92 ),
    .A2(\i43/i48/n72 ),
    .B(\i43/i48/n135 ),
    .Y(\i43/i48/n279 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i267  (.A1(\i43/i48/n54 ),
    .A2(\i43/i48/n58 ),
    .B1(\i43/i48/n50 ),
    .B2(\i43/i48/n92 ),
    .Y(\i43/i48/n278 ));
 AOI22xp5_ASAP7_75t_SL \i43/i48/i268  (.A1(\i43/i48/n55 ),
    .A2(\i43/i48/n44 ),
    .B1(\i43/i48/n85 ),
    .B2(\i43/i48/n48 ),
    .Y(\i43/i48/n277 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i269  (.A1(\i43/i48/n39 ),
    .A2(\i43/i48/n37 ),
    .B(\i43/i48/n171 ),
    .Y(\i43/i48/n275 ));
 NOR3xp33_ASAP7_75t_SL \i43/i48/i27  (.A(\i43/i48/n449 ),
    .B(\i43/i48/n451 ),
    .C(\i43/i48/n434 ),
    .Y(\i43/i48/n488 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i270  (.A1(\i43/i48/n91 ),
    .A2(\i43/i48/n89 ),
    .B1(\i43/i48/n61 ),
    .B2(\i43/i48/n42 ),
    .Y(\i43/i48/n274 ));
 AOI22xp5_ASAP7_75t_SL \i43/i48/i271  (.A1(\i43/i48/n38 ),
    .A2(\i43/i48/n86 ),
    .B1(\i43/i48/n73 ),
    .B2(\i43/i48/n44 ),
    .Y(\i43/i48/n273 ));
 AOI22xp5_ASAP7_75t_SL \i43/i48/i272  (.A1(\i43/i48/n90 ),
    .A2(\i43/i48/n57 ),
    .B1(\i43/i48/n38 ),
    .B2(\i43/i48/n93 ),
    .Y(\i43/i48/n271 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i273  (.A1(\i43/i48/n80 ),
    .A2(\i43/i48/n89 ),
    .B(\i43/i48/n167 ),
    .Y(\i43/i48/n270 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i274  (.A1(\i43/i48/n89 ),
    .A2(\i43/i48/n45 ),
    .B1(\i43/i48/n40 ),
    .B2(\i43/i48/n68 ),
    .Y(\i43/i48/n1 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i275  (.A(\i43/i48/n46 ),
    .B(\i43/i48/n169 ),
    .Y(\i43/i48/n268 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i276  (.A(\i43/i48/n85 ),
    .B(\i43/i48/n168 ),
    .Y(\i43/i48/n267 ));
 NOR2xp33_ASAP7_75t_L \i43/i48/i277  (.A(\i43/i48/n50 ),
    .B(\i43/i48/n153 ),
    .Y(\i43/i48/n266 ));
 INVx1_ASAP7_75t_SL \i43/i48/i278  (.A(\i43/i48/n234 ),
    .Y(\i43/i48/n235 ));
 INVxp33_ASAP7_75t_SL \i43/i48/i279  (.A(\i43/i48/n232 ),
    .Y(\i43/i48/n233 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i28  (.A(\i43/i48/n472 ),
    .B(\i43/i48/n467 ),
    .Y(\i43/i48/n487 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i280  (.A(\i43/i48/n228 ),
    .Y(\i43/i48/n229 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i281  (.A(\i43/i48/n221 ),
    .Y(\i43/i48/n222 ));
 INVx1_ASAP7_75t_SL \i43/i48/i282  (.A(\i43/i48/n213 ),
    .Y(\i43/i48/n212 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i283  (.A1(\i43/i48/n61 ),
    .A2(\i43/i48/n39 ),
    .B1(\i43/i48/n49 ),
    .B2(\i43/i48/n45 ),
    .Y(\i43/i48/n211 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i284  (.A1(\i43/i48/n53 ),
    .A2(\i43/i48/n34 ),
    .B(\i43/i48/n44 ),
    .Y(\i43/i48/n210 ));
 OAI22xp33_ASAP7_75t_SL \i43/i48/i285  (.A1(\i43/i48/n94 ),
    .A2(\i43/i48/n91 ),
    .B1(\i43/i48/n52 ),
    .B2(\i43/i48/n61 ),
    .Y(\i43/i48/n209 ));
 OAI21xp5_ASAP7_75t_SL \i43/i48/i286  (.A1(\i43/i48/n77 ),
    .A2(\i43/i48/n65 ),
    .B(\i43/i48/n36 ),
    .Y(\i43/i48/n208 ));
 AOI21xp33_ASAP7_75t_SL \i43/i48/i287  (.A1(\i43/i48/n66 ),
    .A2(\i43/i48/n72 ),
    .B(\i43/i48/n70 ),
    .Y(\i43/i48/n207 ));
 AOI21xp33_ASAP7_75t_SL \i43/i48/i288  (.A1(\i43/i48/n45 ),
    .A2(\i43/i48/n70 ),
    .B(\i43/i48/n52 ),
    .Y(\i43/i48/n206 ));
 AOI21xp5_ASAP7_75t_SL \i43/i48/i289  (.A1(\i43/i48/n57 ),
    .A2(\i43/i48/n60 ),
    .B(\i43/i48/n129 ),
    .Y(\i43/i48/n205 ));
 AND5x1_ASAP7_75t_SL \i43/i48/i29  (.A(\i43/i48/n446 ),
    .B(\i43/i48/n421 ),
    .C(\i43/i48/n375 ),
    .D(\i43/i48/n410 ),
    .E(\i43/i48/n412 ),
    .Y(\i43/i48/n486 ));
 OAI22xp33_ASAP7_75t_SL \i43/i48/i290  (.A1(\i43/i48/n84 ),
    .A2(\i43/i48/n39 ),
    .B1(\i43/i48/n75 ),
    .B2(\i43/i48/n76 ),
    .Y(\i43/i48/n204 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i291  (.A1(\i43/i48/n75 ),
    .A2(\i43/i48/n54 ),
    .B1(\i43/i48/n40 ),
    .B2(\i43/i48/n61 ),
    .Y(\i43/i48/n203 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i292  (.A1(\i43/i48/n82 ),
    .A2(\i43/i48/n56 ),
    .B1(\i43/i48/n40 ),
    .B2(\i43/i48/n80 ),
    .Y(\i43/i48/n202 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i293  (.A1(\i43/i48/n63 ),
    .A2(\i43/i48/n49 ),
    .B1(\i43/i48/n84 ),
    .B2(\i43/i48/n46 ),
    .Y(\i43/i48/n201 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i294  (.A1(\i43/i48/n50 ),
    .A2(\i43/i48/n91 ),
    .B1(\i43/i48/n39 ),
    .B2(\i43/i48/n63 ),
    .Y(\i43/i48/n200 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i295  (.A1(\i43/i48/n49 ),
    .A2(\i43/i48/n61 ),
    .B1(\i43/i48/n68 ),
    .B2(\i43/i48/n56 ),
    .Y(\i43/i48/n199 ));
 AOI22xp5_ASAP7_75t_SL \i43/i48/i296  (.A1(\i43/i48/n81 ),
    .A2(\i43/i48/n73 ),
    .B1(\i43/i48/n43 ),
    .B2(\i43/i48/n36 ),
    .Y(\i43/i48/n238 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i297  (.A1(\i43/i48/n82 ),
    .A2(\i43/i48/n89 ),
    .B1(\i43/i48/n75 ),
    .B2(\i43/i48/n46 ),
    .Y(\i43/i48/n198 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i298  (.A1(\i43/i48/n43 ),
    .A2(\i43/i48/n88 ),
    .B1(\i43/i48/n83 ),
    .B2(\i43/i48/n33 ),
    .Y(\i43/i48/n197 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i299  (.A1(\i43/i48/n80 ),
    .A2(\i43/i48/n64 ),
    .B1(\i43/i48/n68 ),
    .B2(\i43/i48/n35 ),
    .Y(\i43/i48/n196 ));
 NOR2x1_ASAP7_75t_SL \i43/i48/i3  (.A(\i43/i48/n500 ),
    .B(\i43/i48/n505 ),
    .Y(\i43/n0 [12]));
 NOR3xp33_ASAP7_75t_SL \i43/i48/i30  (.A(\i43/i48/n462 ),
    .B(\i43/i48/n437 ),
    .C(\i43/i48/n424 ),
    .Y(\i43/i48/n485 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i300  (.A1(\i43/i48/n89 ),
    .A2(\i43/i48/n58 ),
    .B1(\i43/i48/n50 ),
    .B2(\i43/i48/n68 ),
    .Y(\i43/i48/n195 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i301  (.A1(\i43/i48/n32 ),
    .A2(\i43/i48/n89 ),
    .B1(\i43/i48/n52 ),
    .B2(\i43/i48/n58 ),
    .Y(\i43/i48/n194 ));
 AOI22xp5_ASAP7_75t_SL \i43/i48/i302  (.A1(\i43/i48/n53 ),
    .A2(\i43/i48/n79 ),
    .B1(\i43/i48/n95 ),
    .B2(\i43/i48/n44 ),
    .Y(\i43/i48/n237 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i303  (.A1(\i43/i48/n70 ),
    .A2(\i43/i48/n64 ),
    .B1(\i43/i48/n72 ),
    .B2(\i43/i48/n37 ),
    .Y(\i43/i48/n236 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i304  (.A1(\i43/i48/n32 ),
    .A2(\i43/i48/n64 ),
    .B1(\i43/i48/n42 ),
    .B2(\i43/i48/n82 ),
    .Y(\i43/i48/n234 ));
 AOI22xp5_ASAP7_75t_SL \i43/i48/i305  (.A1(\i43/i48/n93 ),
    .A2(\i43/i48/n67 ),
    .B1(\i43/i48/n43 ),
    .B2(\i43/i48/n69 ),
    .Y(\i43/i48/n232 ));
 AO22x1_ASAP7_75t_SL \i43/i48/i306  (.A1(\i43/i48/n33 ),
    .A2(\i43/i48/n34 ),
    .B1(\i43/i48/n57 ),
    .B2(\i43/i48/n81 ),
    .Y(\i43/i48/n231 ));
 AOI22xp5_ASAP7_75t_SL \i43/i48/i307  (.A1(\i43/i48/n73 ),
    .A2(\i43/i48/n79 ),
    .B1(\i43/i48/n53 ),
    .B2(\i43/i48/n69 ),
    .Y(\i43/i48/n230 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i308  (.A1(\i43/i48/n58 ),
    .A2(\i43/i48/n64 ),
    .B1(\i43/i48/n54 ),
    .B2(\i43/i48/n63 ),
    .Y(\i43/i48/n228 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i309  (.A(\i43/i48/n187 ),
    .B(\i43/i48/n188 ),
    .Y(\i43/i48/n193 ));
 NOR3xp33_ASAP7_75t_SL \i43/i48/i31  (.A(\i43/i48/n448 ),
    .B(\i43/i48/n436 ),
    .C(\i43/i48/n428 ),
    .Y(\i43/i48/n484 ));
 NAND2xp33_ASAP7_75t_SL \i43/i48/i310  (.A(\i43/i48/n186 ),
    .B(\i43/i48/n176 ),
    .Y(\i43/i48/n192 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i311  (.A1(\i43/i48/n92 ),
    .A2(\i43/i48/n40 ),
    .B1(\i43/i48/n76 ),
    .B2(\i43/i48/n70 ),
    .Y(\i43/i48/n227 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i312  (.A1(\i43/i48/n35 ),
    .A2(\i43/i48/n63 ),
    .B1(\i43/i48/n72 ),
    .B2(\i43/i48/n68 ),
    .Y(\i43/i48/n226 ));
 OAI22xp33_ASAP7_75t_SL \i43/i48/i313  (.A1(\i43/i48/n92 ),
    .A2(\i43/i48/n89 ),
    .B1(\i43/i48/n37 ),
    .B2(\i43/i48/n49 ),
    .Y(\i43/i48/n225 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i314  (.A1(\i43/i48/n92 ),
    .A2(\i43/i48/n49 ),
    .B1(\i43/i48/n42 ),
    .B2(\i43/i48/n75 ),
    .Y(\i43/i48/n224 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i315  (.A1(\i43/i48/n35 ),
    .A2(\i43/i48/n75 ),
    .B1(\i43/i48/n46 ),
    .B2(\i43/i48/n45 ),
    .Y(\i43/i48/n223 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i316  (.A1(\i43/i48/n80 ),
    .A2(\i43/i48/n39 ),
    .B1(\i43/i48/n54 ),
    .B2(\i43/i48/n68 ),
    .Y(\i43/i48/n221 ));
 AOI22xp5_ASAP7_75t_SL \i43/i48/i317  (.A1(\i43/i48/n33 ),
    .A2(\i43/i48/n57 ),
    .B1(\i43/i48/n41 ),
    .B2(\i43/i48/n36 ),
    .Y(\i43/i48/n220 ));
 OAI22xp33_ASAP7_75t_SL \i43/i48/i318  (.A1(\i43/i48/n87 ),
    .A2(\i43/i48/n89 ),
    .B1(\i43/i48/n78 ),
    .B2(\i43/i48/n42 ),
    .Y(\i43/i48/n219 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i319  (.A1(\i43/i48/n46 ),
    .A2(\i43/i48/n58 ),
    .B1(\i43/i48/n91 ),
    .B2(\i43/i48/n76 ),
    .Y(\i43/i48/n218 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i32  (.A(\i43/i48/n444 ),
    .B(\i43/i48/n474 ),
    .Y(\i43/i48/n483 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i320  (.A1(\i43/i48/n68 ),
    .A2(\i43/i48/n64 ),
    .B1(\i43/i48/n50 ),
    .B2(\i43/i48/n37 ),
    .Y(\i43/i48/n217 ));
 AOI22xp5_ASAP7_75t_SL \i43/i48/i321  (.A1(\i43/i48/n79 ),
    .A2(\i43/i48/n57 ),
    .B1(\i43/i48/n95 ),
    .B2(\i43/i48/n69 ),
    .Y(\i43/i48/n216 ));
 OAI22xp5_ASAP7_75t_SL \i43/i48/i322  (.A1(\i43/i48/n78 ),
    .A2(\i43/i48/n89 ),
    .B1(\i43/i48/n50 ),
    .B2(\i43/i48/n32 ),
    .Y(\i43/i48/n215 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i323  (.A(\i43/i48/n139 ),
    .B(\i43/i48/n138 ),
    .Y(\i43/i48/n191 ));
 AOI22xp5_ASAP7_75t_SL \i43/i48/i324  (.A1(\i43/i48/n93 ),
    .A2(\i43/i48/n34 ),
    .B1(\i43/i48/n77 ),
    .B2(\i43/i48/n62 ),
    .Y(\i43/i48/n214 ));
 OA22x2_ASAP7_75t_SL \i43/i48/i325  (.A1(\i43/i48/n61 ),
    .A2(\i43/i48/n64 ),
    .B1(\i43/i48/n58 ),
    .B2(\i43/i48/n76 ),
    .Y(\i43/i48/n213 ));
 INVx1_ASAP7_75t_SL \i43/i48/i326  (.A(\i43/i48/n189 ),
    .Y(\i43/i48/n190 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i327  (.A(\i43/i48/n182 ),
    .Y(\i43/i48/n183 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i328  (.A(\i43/i48/n176 ),
    .Y(\i43/i48/n177 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i329  (.A(\i43/i48/n174 ),
    .Y(\i43/i48/n175 ));
 NOR5xp2_ASAP7_75t_SL \i43/i48/i33  (.A(\i43/i48/n400 ),
    .B(\i43/i48/n408 ),
    .C(\i43/i48/n305 ),
    .D(\i43/i48/n397 ),
    .E(\i43/i48/n401 ),
    .Y(\i43/i48/n482 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i330  (.A(\i43/i48/n168 ),
    .Y(\i43/i48/n169 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i331  (.A(\i43/i48/n165 ),
    .Y(\i43/i48/n166 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i332  (.A(\i43/i48/n160 ),
    .Y(\i43/i48/n161 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i333  (.A(\i43/i48/n155 ),
    .Y(\i43/i48/n156 ));
 INVx1_ASAP7_75t_SL \i43/i48/i334  (.A(\i43/i48/n153 ),
    .Y(\i43/i48/n154 ));
 INVx1_ASAP7_75t_SL \i43/i48/i335  (.A(\i43/i48/n151 ),
    .Y(\i43/i48/n152 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i336  (.A(\i43/i48/n149 ),
    .Y(\i43/i48/n150 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i337  (.A(\i43/i48/n147 ),
    .Y(\i43/i48/n148 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i338  (.A(\i43/i48/n85 ),
    .B(\i43/i48/n51 ),
    .Y(\i43/i48/n146 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i339  (.A(\i43/i48/n77 ),
    .B(\i43/i48/n81 ),
    .Y(\i43/i48/n189 ));
 NAND5xp2_ASAP7_75t_SL \i43/i48/i34  (.A(\i43/i48/n390 ),
    .B(\i43/i48/n417 ),
    .C(\i43/i48/n352 ),
    .D(\i43/i48/n318 ),
    .E(\i43/i48/n349 ),
    .Y(\i43/i48/n481 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i340  (.A(\i43/i48/n41 ),
    .B(\i43/i48/n90 ),
    .Y(\i43/i48/n145 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i341  (.A(\i43/i48/n90 ),
    .B(\i43/i48/n48 ),
    .Y(\i43/i48/n144 ));
 NAND2xp33_ASAP7_75t_SL \i43/i48/i342  (.A(\i43/i48/n46 ),
    .B(\i43/i48/n64 ),
    .Y(\i43/i48/n143 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i343  (.A(\i43/i48/n36 ),
    .B(\i43/i48/n65 ),
    .Y(\i43/i48/n188 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i344  (.A(\i43/i48/n95 ),
    .B(\i43/i48/n93 ),
    .Y(\i43/i48/n187 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i345  (.A(\i43/i48/n67 ),
    .B(\i43/i48/n59 ),
    .Y(\i43/i48/n186 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i346  (.A(\i43/i48/n85 ),
    .B(\i43/i48/n71 ),
    .Y(\i43/i48/n142 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i347  (.A(\i43/i48/n58 ),
    .B(\i43/i48/n50 ),
    .Y(\i43/i48/n141 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i348  (.A(\i43/i48/n55 ),
    .B(\i43/i48/n83 ),
    .Y(\i43/i48/n185 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i349  (.A(\i43/i48/n69 ),
    .B(\i43/i48/n41 ),
    .Y(\i43/i48/n140 ));
 NOR2xp33_ASAP7_75t_L \i43/i48/i35  (.A(\i43/i48/n455 ),
    .B(\i43/i48/n478 ),
    .Y(\i43/i48/n480 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i350  (.A(\i43/i48/n77 ),
    .B(\i43/i48/n93 ),
    .Y(\i43/i48/n184 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i351  (.A(\i43/i48/n75 ),
    .B(\i43/i48/n40 ),
    .Y(\i43/i48/n182 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i352  (.A(\i43/i48/n69 ),
    .B(\i43/i48/n67 ),
    .Y(\i43/i48/n181 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i353  (.A(\i43/i48/n79 ),
    .B(\i43/i48/n51 ),
    .Y(\i43/i48/n180 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i354  (.A(\i43/i48/n93 ),
    .B(\i43/i48/n65 ),
    .Y(\i43/i48/n179 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i355  (.A(\i43/i48/n79 ),
    .B(\i43/i48/n95 ),
    .Y(\i43/i48/n178 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i356  (.A(\i43/i48/n74 ),
    .B(\i43/i48/n65 ),
    .Y(\i43/i48/n176 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i357  (.A(\i43/i48/n86 ),
    .B(\i43/i48/n77 ),
    .Y(\i43/i48/n174 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i358  (.A(\i43/i48/n85 ),
    .B(\i43/i48/n69 ),
    .Y(\i43/i48/n173 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i359  (.A(\i43/i48/n95 ),
    .B(\i43/i48/n36 ),
    .Y(\i43/i48/n172 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i36  (.A(\i43/i48/n416 ),
    .B(\i43/i48/n477 ),
    .Y(\i43/i48/n479 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i360  (.A(\i43/i48/n44 ),
    .B(\i43/i48/n65 ),
    .Y(\i43/i48/n171 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i361  (.A(\i43/i48/n91 ),
    .B(\i43/i48/n46 ),
    .Y(\i43/i48/n170 ));
 NAND2xp5_ASAP7_75t_L \i43/i48/i362  (.A(\i43/i48/n35 ),
    .B(\i43/i48/n94 ),
    .Y(\i43/i48/n168 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i363  (.A(\i43/i48/n95 ),
    .B(\i43/i48/n33 ),
    .Y(\i43/i48/n167 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i364  (.A(\i43/i48/n95 ),
    .B(\i43/i48/n43 ),
    .Y(\i43/i48/n165 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i365  (.A(\i43/i48/n57 ),
    .B(\i43/i48/n59 ),
    .Y(\i43/i48/n164 ));
 NAND2xp33_ASAP7_75t_SL \i43/i48/i366  (.A(\i43/i48/n61 ),
    .B(\i43/i48/n87 ),
    .Y(\i43/i48/n163 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i367  (.A(\i43/i48/n59 ),
    .B(\i43/i48/n41 ),
    .Y(\i43/i48/n162 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i368  (.A(\i43/i48/n73 ),
    .B(\i43/i48/n59 ),
    .Y(\i43/i48/n160 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i369  (.A(\i43/i48/n77 ),
    .B(\i43/i48/n83 ),
    .Y(\i43/i48/n159 ));
 INVx1_ASAP7_75t_SL \i43/i48/i37  (.A(\i43/i48/n509 ),
    .Y(\i43/i48/n475 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i370  (.A(\i43/i48/n85 ),
    .B(\i43/i48/n57 ),
    .Y(\i43/i48/n158 ));
 NOR2xp33_ASAP7_75t_L \i43/i48/i371  (.A(\i43/i48/n60 ),
    .B(\i43/i48/n69 ),
    .Y(\i43/i48/n157 ));
 NAND2xp5_ASAP7_75t_L \i43/i48/i372  (.A(\i43/i48/n37 ),
    .B(\i43/i48/n68 ),
    .Y(\i43/i48/n155 ));
 NOR2x1_ASAP7_75t_SL \i43/i48/i373  (.A(\i43/i48/n62 ),
    .B(\i43/i48/n71 ),
    .Y(\i43/i48/n153 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i374  (.A(\i43/i48/n88 ),
    .B(\i43/i48/n36 ),
    .Y(\i43/i48/n151 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i375  (.A(\i43/i48/n86 ),
    .B(\i43/i48/n62 ),
    .Y(\i43/i48/n149 ));
 NAND2x1_ASAP7_75t_SL \i43/i48/i376  (.A(\i43/i48/n84 ),
    .B(\i43/i48/n63 ),
    .Y(\i43/i48/n0 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i377  (.A(\i43/i48/n32 ),
    .B(\i43/i48/n91 ),
    .Y(\i43/i48/n147 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i378  (.A(\i43/i48/n130 ),
    .Y(\i43/i48/n131 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i379  (.A(\i43/i48/n121 ),
    .Y(\i43/i48/n122 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i38  (.A(\i43/i48/n453 ),
    .B(\i43/i48/n422 ),
    .Y(\i43/i48/n473 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i380  (.A(\i43/i48/n118 ),
    .Y(\i43/i48/n119 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i381  (.A(\i43/i48/n55 ),
    .B(\i43/i48/n36 ),
    .Y(\i43/i48/n116 ));
 NAND2xp33_ASAP7_75t_SL \i43/i48/i382  (.A(\i43/i48/n70 ),
    .B(\i43/i48/n61 ),
    .Y(\i43/i48/n115 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i383  (.A(\i43/i48/n48 ),
    .B(\i43/i48/n57 ),
    .Y(\i43/i48/n114 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i384  (.A(\i43/i48/n51 ),
    .B(\i43/i48/n83 ),
    .Y(\i43/i48/n113 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i385  (.A(\i43/i48/n57 ),
    .B(\i43/i48/n36 ),
    .Y(\i43/i48/n139 ));
 NAND2xp33_ASAP7_75t_SL \i43/i48/i386  (.A(\i43/i48/n82 ),
    .B(\i43/i48/n45 ),
    .Y(\i43/i48/n112 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i387  (.A(\i43/i48/n71 ),
    .B(\i43/i48/n55 ),
    .Y(\i43/i48/n111 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i388  (.A(\i43/i48/n33 ),
    .B(\i43/i48/n38 ),
    .Y(\i43/i48/n110 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i389  (.A(\i43/i48/n75 ),
    .B(\i43/i48/n82 ),
    .Y(\i43/i48/n109 ));
 NAND2xp33_ASAP7_75t_L \i43/i48/i39  (.A(\i43/i48/n453 ),
    .B(\i43/i48/n433 ),
    .Y(\i43/i48/n472 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i390  (.A(\i43/i48/n93 ),
    .B(\i43/i48/n53 ),
    .Y(\i43/i48/n108 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i391  (.A(\i43/i48/n44 ),
    .B(\i43/i48/n43 ),
    .Y(\i43/i48/n138 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i392  (.A(\i43/i48/n60 ),
    .B(\i43/i48/n34 ),
    .Y(\i43/i48/n107 ));
 NAND2xp33_ASAP7_75t_SL \i43/i48/i393  (.A(\i43/i48/n39 ),
    .B(\i43/i48/n66 ),
    .Y(\i43/i48/n106 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i394  (.A(\i43/i48/n47 ),
    .B(\i43/i48/n33 ),
    .Y(\i43/i48/n105 ));
 NAND2xp5_ASAP7_75t_L \i43/i48/i395  (.A(\i43/i48/n42 ),
    .B(\i43/i48/n66 ),
    .Y(\i43/i48/n104 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i396  (.A(\i43/i48/n38 ),
    .B(\i43/i48/n73 ),
    .Y(\i43/i48/n103 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i397  (.A(\i43/i48/n73 ),
    .B(\i43/i48/n60 ),
    .Y(\i43/i48/n137 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i398  (.A(\i43/i48/n41 ),
    .B(\i43/i48/n73 ),
    .Y(\i43/i48/n136 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i399  (.A(\i43/i48/n74 ),
    .B(\i43/i48/n48 ),
    .Y(\i43/i48/n135 ));
 AND5x1_ASAP7_75t_SL \i43/i48/i4  (.A(\i43/i48/n501 ),
    .B(\i43/i48/n498 ),
    .C(\i43/i48/n477 ),
    .D(\i43/i48/n499 ),
    .E(\i43/i48/n468 ),
    .Y(\i43/n0 [11]));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i40  (.A(\i43/i48/n450 ),
    .B(\i43/i48/n432 ),
    .Y(\i43/i48/n471 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i400  (.A(\i43/i48/n72 ),
    .B(\i43/i48/n45 ),
    .Y(\i43/i48/n102 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i401  (.A(\i43/i48/n67 ),
    .B(\i43/i48/n36 ),
    .Y(\i43/i48/n134 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i402  (.A(\i43/i48/n47 ),
    .B(\i43/i48/n93 ),
    .Y(\i43/i48/n133 ));
 NOR2xp33_ASAP7_75t_L \i43/i48/i403  (.A(\i43/i48/n35 ),
    .B(\i43/i48/n37 ),
    .Y(\i43/i48/n132 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i404  (.A(\i43/i48/n42 ),
    .B(\i43/i48/n75 ),
    .Y(\i43/i48/n101 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i405  (.A(\i43/i48/n71 ),
    .B(\i43/i48/n34 ),
    .Y(\i43/i48/n100 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i406  (.A(\i43/i48/n51 ),
    .B(\i43/i48/n44 ),
    .Y(\i43/i48/n130 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i407  (.A(\i43/i48/n92 ),
    .B(\i43/i48/n42 ),
    .Y(\i43/i48/n129 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i408  (.A(\i43/i48/n47 ),
    .B(\i43/i48/n81 ),
    .Y(\i43/i48/n128 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i409  (.A(\i43/i48/n47 ),
    .B(\i43/i48/n60 ),
    .Y(\i43/i48/n127 ));
 NAND4xp25_ASAP7_75t_SL \i43/i48/i41  (.A(\i43/i48/n415 ),
    .B(\i43/i48/n308 ),
    .C(\i43/i48/n311 ),
    .D(\i43/i48/n343 ),
    .Y(\i43/i48/n470 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i410  (.A(\i43/i48/n74 ),
    .B(\i43/i48/n51 ),
    .Y(\i43/i48/n126 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i411  (.A(\i43/i48/n38 ),
    .B(\i43/i48/n93 ),
    .Y(\i43/i48/n99 ));
 NOR2xp33_ASAP7_75t_L \i43/i48/i412  (.A(\i43/i48/n50 ),
    .B(\i43/i48/n80 ),
    .Y(\i43/i48/n125 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i413  (.A(\i43/i48/n50 ),
    .B(\i43/i48/n92 ),
    .Y(\i43/i48/n98 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i414  (.A(\i43/i48/n61 ),
    .B(\i43/i48/n42 ),
    .Y(\i43/i48/n97 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i415  (.A(\i43/i48/n93 ),
    .B(\i43/i48/n57 ),
    .Y(\i43/i48/n124 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i416  (.A(\i43/i48/n55 ),
    .B(\i43/i48/n44 ),
    .Y(\i43/i48/n96 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i417  (.A(\i43/i48/n79 ),
    .B(\i43/i48/n38 ),
    .Y(\i43/i48/n123 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i418  (.A(\i43/i48/n49 ),
    .B(\i43/i48/n32 ),
    .Y(\i43/i48/n121 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i419  (.A(\i43/i48/n33 ),
    .B(\i43/i48/n53 ),
    .Y(\i43/i48/n120 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i42  (.A(\i43/i48/n433 ),
    .B(\i43/i48/n442 ),
    .Y(\i43/i48/n478 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i420  (.A(\i43/i48/n83 ),
    .B(\i43/i48/n53 ),
    .Y(\i43/i48/n118 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i421  (.A(\i43/i48/n60 ),
    .B(\i43/i48/n51 ),
    .Y(\i43/i48/n117 ));
 INVx1_ASAP7_75t_SL \i43/i48/i422  (.A(\i43/i48/n95 ),
    .Y(\i43/i48/n94 ));
 INVx2_ASAP7_75t_SL \i43/i48/i423  (.A(\i43/i48/n93 ),
    .Y(\i43/i48/n92 ));
 INVx1_ASAP7_75t_SL \i43/i48/i424  (.A(\i43/i48/n91 ),
    .Y(\i43/i48/n90 ));
 INVx2_ASAP7_75t_SL \i43/i48/i425  (.A(\i43/i48/n89 ),
    .Y(\i43/i48/n88 ));
 INVx2_ASAP7_75t_SL \i43/i48/i426  (.A(\i43/i48/n87 ),
    .Y(\i43/i48/n86 ));
 INVx2_ASAP7_75t_SL \i43/i48/i427  (.A(\i43/i48/n85 ),
    .Y(\i43/i48/n84 ));
 INVx3_ASAP7_75t_SL \i43/i48/i428  (.A(\i43/i48/n83 ),
    .Y(\i43/i48/n82 ));
 INVx2_ASAP7_75t_SL \i43/i48/i429  (.A(\i43/i48/n81 ),
    .Y(\i43/i48/n80 ));
 AND4x1_ASAP7_75t_SL \i43/i48/i43  (.A(\i43/i48/n435 ),
    .B(\i43/i48/n415 ),
    .C(\i43/i48/n353 ),
    .D(\i43/i48/n193 ),
    .Y(\i43/i48/n469 ));
 INVx2_ASAP7_75t_SL \i43/i48/i430  (.A(\i43/i48/n79 ),
    .Y(\i43/i48/n78 ));
 INVx2_ASAP7_75t_SL \i43/i48/i431  (.A(\i43/i48/n77 ),
    .Y(\i43/i48/n76 ));
 INVx2_ASAP7_75t_SL \i43/i48/i432  (.A(\i43/i48/n75 ),
    .Y(\i43/i48/n74 ));
 INVx2_ASAP7_75t_SL \i43/i48/i433  (.A(\i43/i48/n73 ),
    .Y(\i43/i48/n72 ));
 INVx2_ASAP7_75t_SL \i43/i48/i434  (.A(\i43/i48/n71 ),
    .Y(\i43/i48/n70 ));
 INVx2_ASAP7_75t_SL \i43/i48/i435  (.A(\i43/i48/n69 ),
    .Y(\i43/i48/n68 ));
 INVx2_ASAP7_75t_SL \i43/i48/i436  (.A(\i43/i48/n67 ),
    .Y(\i43/i48/n66 ));
 INVx2_ASAP7_75t_SL \i43/i48/i437  (.A(\i43/i48/n65 ),
    .Y(\i43/i48/n64 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i438  (.A(\i43/i48/n25 ),
    .B(\i43/i48/n15 ),
    .Y(\i43/i48/n95 ));
 AND2x4_ASAP7_75t_SL \i43/i48/i439  (.A(\i43/i48/n5 ),
    .B(\i43/i48/n6 ),
    .Y(\i43/i48/n93 ));
 AND4x1_ASAP7_75t_SL \i43/i48/i44  (.A(\i43/i48/n380 ),
    .B(\i43/i48/n317 ),
    .C(\i43/i48/n368 ),
    .D(\i43/i48/n189 ),
    .Y(\i43/i48/n477 ));
 OR2x2_ASAP7_75t_SL \i43/i48/i440  (.A(\i43/i48/n27 ),
    .B(\i43/i48/n11 ),
    .Y(\i43/i48/n91 ));
 OR2x2_ASAP7_75t_SL \i43/i48/i441  (.A(\i43/i48/n28 ),
    .B(\i43/i48/n9 ),
    .Y(\i43/i48/n89 ));
 OR2x6_ASAP7_75t_SL \i43/i48/i442  (.A(\i43/i48/n7 ),
    .B(\i43/i48/n11 ),
    .Y(\i43/i48/n87 ));
 AND2x4_ASAP7_75t_SL \i43/i48/i443  (.A(\i43/i48/n4 ),
    .B(\i43/i48/n19 ),
    .Y(\i43/i48/n85 ));
 AND2x4_ASAP7_75t_SL \i43/i48/i444  (.A(\i43/i48/n10 ),
    .B(\i43/i48/n22 ),
    .Y(\i43/i48/n83 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i445  (.A(\i43/i48/n6 ),
    .B(\i43/i48/n19 ),
    .Y(\i43/i48/n81 ));
 AND2x4_ASAP7_75t_SL \i43/i48/i446  (.A(\i43/i48/n5 ),
    .B(\i43/i48/n26 ),
    .Y(\i43/i48/n79 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i447  (.A(\i43/i48/n16 ),
    .B(\i43/i48/n15 ),
    .Y(\i43/i48/n77 ));
 OR2x2_ASAP7_75t_SL \i43/i48/i448  (.A(\i43/i48/n3 ),
    .B(\i43/i48/n31 ),
    .Y(\i43/i48/n75 ));
 AND2x4_ASAP7_75t_SL \i43/i48/i449  (.A(\i43/i48/n25 ),
    .B(\i43/i48/n12 ),
    .Y(\i43/i48/n73 ));
 NOR2x1_ASAP7_75t_SL \i43/i48/i45  (.A(\i43/i48/n306 ),
    .B(\i43/i48/n451 ),
    .Y(\i43/i48/n476 ));
 AND2x4_ASAP7_75t_SL \i43/i48/i450  (.A(\i43/i48/n4 ),
    .B(\i43/i48/n10 ),
    .Y(\i43/i48/n71 ));
 AND2x4_ASAP7_75t_SL \i43/i48/i451  (.A(\i43/i48/n5 ),
    .B(\i43/i48/n4 ),
    .Y(\i43/i48/n69 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i452  (.A(\i43/i48/n16 ),
    .B(\i43/i48/n29 ),
    .Y(\i43/i48/n67 ));
 AND2x4_ASAP7_75t_SL \i43/i48/i453  (.A(\i43/i48/n8 ),
    .B(\i43/i48/n12 ),
    .Y(\i43/i48/n65 ));
 INVx2_ASAP7_75t_SL \i43/i48/i454  (.A(\i43/i48/n63 ),
    .Y(\i43/i48/n62 ));
 INVx3_ASAP7_75t_SL \i43/i48/i455  (.A(\i43/i48/n61 ),
    .Y(\i43/i48/n60 ));
 INVx2_ASAP7_75t_SL \i43/i48/i456  (.A(\i43/i48/n59 ),
    .Y(\i43/i48/n58 ));
 INVx1_ASAP7_75t_SL \i43/i48/i457  (.A(\i43/i48/n57 ),
    .Y(\i43/i48/n56 ));
 INVx2_ASAP7_75t_SL \i43/i48/i458  (.A(\i43/i48/n55 ),
    .Y(\i43/i48/n54 ));
 INVx3_ASAP7_75t_SL \i43/i48/i459  (.A(\i43/i48/n53 ),
    .Y(\i43/i48/n52 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i46  (.A(\i43/i48/n392 ),
    .B(\i43/i48/n426 ),
    .Y(\i43/i48/n474 ));
 INVx2_ASAP7_75t_SL \i43/i48/i460  (.A(\i43/i48/n51 ),
    .Y(\i43/i48/n50 ));
 INVx2_ASAP7_75t_SL \i43/i48/i461  (.A(\i43/i48/n49 ),
    .Y(\i43/i48/n48 ));
 INVx2_ASAP7_75t_SL \i43/i48/i462  (.A(\i43/i48/n47 ),
    .Y(\i43/i48/n46 ));
 INVx4_ASAP7_75t_SL \i43/i48/i463  (.A(\i43/i48/n45 ),
    .Y(\i43/i48/n44 ));
 INVx4_ASAP7_75t_SL \i43/i48/i464  (.A(\i43/i48/n43 ),
    .Y(\i43/i48/n42 ));
 INVx2_ASAP7_75t_SL \i43/i48/i465  (.A(\i43/i48/n41 ),
    .Y(\i43/i48/n40 ));
 INVx2_ASAP7_75t_SL \i43/i48/i466  (.A(\i43/i48/n39 ),
    .Y(\i43/i48/n38 ));
 INVx2_ASAP7_75t_SL \i43/i48/i467  (.A(\i43/i48/n37 ),
    .Y(\i43/i48/n36 ));
 INVx3_ASAP7_75t_SL \i43/i48/i468  (.A(\i43/i48/n35 ),
    .Y(\i43/i48/n34 ));
 INVx2_ASAP7_75t_SL \i43/i48/i469  (.A(\i43/i48/n33 ),
    .Y(\i43/i48/n32 ));
 INVx1_ASAP7_75t_SL \i43/i48/i47  (.A(\i43/i48/n466 ),
    .Y(\i43/i48/n467 ));
 NAND2x1p5_ASAP7_75t_SL \i43/i48/i470  (.A(\i43/i48/n22 ),
    .B(\i43/i48/n5 ),
    .Y(\i43/i48/n63 ));
 OR2x2_ASAP7_75t_SL \i43/i48/i471  (.A(\i43/i48/n27 ),
    .B(\i43/i48/n20 ),
    .Y(\i43/i48/n61 ));
 AND2x4_ASAP7_75t_SL \i43/i48/i472  (.A(\i43/i48/n6 ),
    .B(\i43/i48/n30 ),
    .Y(\i43/i48/n59 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i473  (.A(\i43/i48/n25 ),
    .B(\i43/i48/n18 ),
    .Y(\i43/i48/n57 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i474  (.A(\i43/i48/n8 ),
    .B(\i43/i48/n18 ),
    .Y(\i43/i48/n55 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i475  (.A(\i43/i48/n16 ),
    .B(\i43/i48/n12 ),
    .Y(\i43/i48/n53 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i476  (.A(\i43/i48/n25 ),
    .B(\i43/i48/n29 ),
    .Y(\i43/i48/n51 ));
 OR2x2_ASAP7_75t_SL \i43/i48/i477  (.A(\i43/i48/n17 ),
    .B(\i43/i48/n24 ),
    .Y(\i43/i48/n49 ));
 AND2x4_ASAP7_75t_SL \i43/i48/i478  (.A(\i43/i48/n23 ),
    .B(\i43/i48/n15 ),
    .Y(\i43/i48/n47 ));
 OR2x2_ASAP7_75t_SL \i43/i48/i479  (.A(\i43/i48/n27 ),
    .B(\i43/i48/n31 ),
    .Y(\i43/i48/n45 ));
 NAND2xp5_ASAP7_75t_L \i43/i48/i48  (.A(\i43/i48/n435 ),
    .B(\i43/i48/n419 ),
    .Y(\i43/i48/n464 ));
 AND2x4_ASAP7_75t_SL \i43/i48/i480  (.A(\i43/i48/n23 ),
    .B(\i43/i48/n29 ),
    .Y(\i43/i48/n43 ));
 AND2x4_ASAP7_75t_SL \i43/i48/i481  (.A(\i43/i48/n16 ),
    .B(\i43/i48/n18 ),
    .Y(\i43/i48/n41 ));
 OR2x2_ASAP7_75t_SL \i43/i48/i482  (.A(\i43/i48/n14 ),
    .B(\i43/i48/n9 ),
    .Y(\i43/i48/n39 ));
 OR2x6_ASAP7_75t_SL \i43/i48/i483  (.A(\i43/i48/n20 ),
    .B(\i43/i48/n21 ),
    .Y(\i43/i48/n37 ));
 OR2x6_ASAP7_75t_SL \i43/i48/i484  (.A(\i43/i48/n24 ),
    .B(\i43/i48/n13 ),
    .Y(\i43/i48/n35 ));
 AND2x4_ASAP7_75t_SL \i43/i48/i485  (.A(\i43/i48/n30 ),
    .B(\i43/i48/n22 ),
    .Y(\i43/i48/n33 ));
 INVx2_ASAP7_75t_SL \i43/i48/i486  (.A(\i43/i48/n31 ),
    .Y(\i43/i48/n30 ));
 INVx2_ASAP7_75t_SL \i43/i48/i487  (.A(\i43/i48/n28 ),
    .Y(\i43/i48/n29 ));
 INVxp67_ASAP7_75t_SL \i43/i48/i488  (.A(\i43/i48/n27 ),
    .Y(\i43/i48/n26 ));
 INVx2_ASAP7_75t_SL \i43/i48/i489  (.A(\i43/i48/n24 ),
    .Y(\i43/i48/n23 ));
 AND3x1_ASAP7_75t_SL \i43/i48/i49  (.A(\i43/i48/n420 ),
    .B(\i43/i48/n405 ),
    .C(\i43/i48/n391 ),
    .Y(\i43/i48/n463 ));
 INVx3_ASAP7_75t_SL \i43/i48/i490  (.A(\i43/i48/n21 ),
    .Y(\i43/i48/n22 ));
 INVx2_ASAP7_75t_SL \i43/i48/i491  (.A(\i43/i48/n20 ),
    .Y(\i43/i48/n19 ));
 INVx1_ASAP7_75t_SL \i43/i48/i492  (.A(\i43/i48/n17 ),
    .Y(\i43/i48/n18 ));
 OR2x2_ASAP7_75t_SL \i43/i48/i493  (.A(n79),
    .B(n34[5]),
    .Y(\i43/i48/n31 ));
 OR2x2_ASAP7_75t_SL \i43/i48/i494  (.A(n80),
    .B(n34[0]),
    .Y(\i43/i48/n28 ));
 OR2x2_ASAP7_75t_SL \i43/i48/i495  (.A(n77),
    .B(n34[7]),
    .Y(\i43/i48/n27 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i496  (.A(n34[1]),
    .B(n81),
    .Y(\i43/i48/n25 ));
 NAND2x1_ASAP7_75t_SL \i43/i48/i497  (.A(n34[2]),
    .B(n82),
    .Y(\i43/i48/n24 ));
 OR2x2_ASAP7_75t_SL \i43/i48/i498  (.A(\i43/i48/n2 ),
    .B(n34[6]),
    .Y(\i43/i48/n21 ));
 OR2x2_ASAP7_75t_SL \i43/i48/i499  (.A(n78),
    .B(n34[4]),
    .Y(\i43/i48/n20 ));
 NAND5xp2_ASAP7_75t_SL \i43/i48/i5  (.A(\i43/i48/n466 ),
    .B(\i43/i48/n476 ),
    .C(\i43/i48/n471 ),
    .D(\i43/i48/n460 ),
    .E(\i43/i48/n454 ),
    .Y(\i43/i48/n507 ));
 NAND4xp25_ASAP7_75t_SL \i43/i48/i50  (.A(\i43/i48/n418 ),
    .B(\i43/i48/n384 ),
    .C(\i43/i48/n312 ),
    .D(\i43/i48/n309 ),
    .Y(\i43/i48/n462 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i500  (.A(n34[0]),
    .B(n80),
    .Y(\i43/i48/n17 ));
 INVx1_ASAP7_75t_SL \i43/i48/i501  (.A(\i43/i48/n14 ),
    .Y(\i43/i48/n15 ));
 INVx2_ASAP7_75t_SL \i43/i48/i502  (.A(\i43/i48/n12 ),
    .Y(\i43/i48/n13 ));
 INVx1_ASAP7_75t_SL \i43/i48/i503  (.A(\i43/i48/n11 ),
    .Y(\i43/i48/n10 ));
 INVx1_ASAP7_75t_SL \i43/i48/i504  (.A(\i43/i48/n9 ),
    .Y(\i43/i48/n8 ));
 INVx1_ASAP7_75t_SL \i43/i48/i505  (.A(\i43/i48/n6 ),
    .Y(\i43/i48/n7 ));
 INVx2_ASAP7_75t_SL \i43/i48/i506  (.A(\i43/i48/n3 ),
    .Y(\i43/i48/n4 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i507  (.A(n34[2]),
    .B(n34[1]),
    .Y(\i43/i48/n16 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i508  (.A(n34[3]),
    .B(n34[0]),
    .Y(\i43/i48/n14 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i509  (.A(n80),
    .B(n83),
    .Y(\i43/i48/n12 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i51  (.A(\i43/i48/n247 ),
    .B(\i43/i48/n510 ),
    .Y(\i43/i48/n461 ));
 OR2x2_ASAP7_75t_SL \i43/i48/i510  (.A(n34[5]),
    .B(n34[4]),
    .Y(\i43/i48/n11 ));
 OR2x2_ASAP7_75t_SL \i43/i48/i511  (.A(n34[2]),
    .B(n34[1]),
    .Y(\i43/i48/n9 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i512  (.A(\i43/i48/n2 ),
    .B(n77),
    .Y(\i43/i48/n6 ));
 AND2x2_ASAP7_75t_SL \i43/i48/i513  (.A(n34[5]),
    .B(n34[4]),
    .Y(\i43/i48/n5 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i514  (.A(n34[7]),
    .B(n34[6]),
    .Y(\i43/i48/n3 ));
 INVx1_ASAP7_75t_SL \i43/i48/i515  (.A(n34[7]),
    .Y(\i43/i48/n2 ));
 OR4x1_ASAP7_75t_SL \i43/i48/i516  (.A(\i43/i48/n450 ),
    .B(\i43/i48/n278 ),
    .C(\i43/i48/n248 ),
    .D(\i43/i48/n226 ),
    .Y(\i43/i48/n508 ));
 NAND5xp2_ASAP7_75t_SL \i43/i48/i517  (.A(\i43/i48/n452 ),
    .B(\i43/i48/n288 ),
    .C(\i43/i48/n277 ),
    .D(\i43/i48/n220 ),
    .E(\i43/i48/n414 ),
    .Y(\i43/i48/n509 ));
 AND3x1_ASAP7_75t_SL \i43/i48/i518  (.A(\i43/i48/n326 ),
    .B(\i43/i48/n267 ),
    .C(\i43/i48/n329 ),
    .Y(\i43/i48/n510 ));
 OR3x1_ASAP7_75t_SL \i43/i48/i519  (.A(\i43/i48/n223 ),
    .B(\i43/i48/n132 ),
    .C(\i43/i48/n199 ),
    .Y(\i43/i48/n511 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i52  (.A(\i43/i48/n411 ),
    .B(\i43/i48/n441 ),
    .Y(\i43/i48/n460 ));
 NAND3xp33_ASAP7_75t_SL \i43/i48/i520  (.A(\i43/i48/n230 ),
    .B(\i43/i48/n117 ),
    .C(\i43/i48/n107 ),
    .Y(\i43/i48/n512 ));
 NAND3xp33_ASAP7_75t_SL \i43/i48/i521  (.A(\i43/i48/n513 ),
    .B(\i43/i48/n302 ),
    .C(\i43/i48/n151 ),
    .Y(\i43/i48/n514 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i522  (.A(\i43/i48/n228 ),
    .B(\i43/i48/n124 ),
    .Y(\i43/i48/n513 ));
 NOR3xp33_ASAP7_75t_SL \i43/i48/i53  (.A(\i43/i48/n383 ),
    .B(\i43/i48/n398 ),
    .C(\i43/i48/n304 ),
    .Y(\i43/i48/n459 ));
 AOI211xp5_ASAP7_75t_SL \i43/i48/i54  (.A1(\i43/i48/n378 ),
    .A2(\i43/i48/n4 ),
    .B(\i43/i48/n394 ),
    .C(\i43/i48/n396 ),
    .Y(\i43/i48/n458 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i55  (.A(\i43/i48/n425 ),
    .B(\i43/i48/n431 ),
    .Y(\i43/i48/n457 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i56  (.A(\i43/i48/n393 ),
    .B(\i43/i48/n434 ),
    .Y(\i43/i48/n456 ));
 NOR2xp33_ASAP7_75t_L \i43/i48/i57  (.A(\i43/i48/n411 ),
    .B(\i43/i48/n430 ),
    .Y(\i43/i48/n468 ));
 OA211x2_ASAP7_75t_SL \i43/i48/i58  (.A1(\i43/i48/n91 ),
    .A2(\i43/i48/n66 ),
    .B(\i43/i48/n391 ),
    .C(\i43/i48/n370 ),
    .Y(\i43/i48/n466 ));
 NAND3xp33_ASAP7_75t_SL \i43/i48/i59  (.A(\i43/i48/n353 ),
    .B(\i43/i48/n379 ),
    .C(\i43/i48/n320 ),
    .Y(\i43/i48/n465 ));
 AND4x1_ASAP7_75t_SL \i43/i48/i6  (.A(\i43/i48/n495 ),
    .B(\i43/i48/n499 ),
    .C(\i43/i48/n484 ),
    .D(\i43/i48/n457 ),
    .Y(\i43/n0 [8]));
 INVxp67_ASAP7_75t_SL \i43/i48/i60  (.A(\i43/i48/n510 ),
    .Y(\i43/i48/n449 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i61  (.A(\i43/i48/n407 ),
    .B(\i43/i48/n392 ),
    .Y(\i43/i48/n448 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i62  (.A(\i43/i48/n300 ),
    .B(\i43/i48/n407 ),
    .Y(\i43/i48/n447 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i63  (.A(\i43/i48/n390 ),
    .B(\i43/i48/n387 ),
    .Y(\i43/i48/n455 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i64  (.A(\i43/i48/n511 ),
    .B(\i43/i48/n382 ),
    .Y(\i43/i48/n446 ));
 NAND2xp5_ASAP7_75t_L \i43/i48/i65  (.A(\i43/i48/n388 ),
    .B(\i43/i48/n310 ),
    .Y(\i43/i48/n445 ));
 NOR3xp33_ASAP7_75t_SL \i43/i48/i66  (.A(\i43/i48/n413 ),
    .B(\i43/i48/n342 ),
    .C(\i43/i48/n344 ),
    .Y(\i43/i48/n454 ));
 NAND3xp33_ASAP7_75t_SL \i43/i48/i67  (.A(\i43/i48/n389 ),
    .B(\i43/i48/n341 ),
    .C(\i43/i48/n216 ),
    .Y(\i43/i48/n444 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i68  (.A(\i43/i48/n299 ),
    .B(\i43/i48/n374 ),
    .Y(\i43/i48/n443 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i69  (.A(\i43/i48/n386 ),
    .B(\i43/i48/n512 ),
    .Y(\i43/i48/n442 ));
 AND4x1_ASAP7_75t_L \i43/i48/i7  (.A(\i43/i48/n485 ),
    .B(\i43/i48/n490 ),
    .C(\i43/i48/n498 ),
    .D(\i43/i48/n487 ),
    .Y(\i43/n0 [15]));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i70  (.A(\i43/i48/n353 ),
    .B(\i43/i48/n399 ),
    .Y(\i43/i48/n441 ));
 OA211x2_ASAP7_75t_SL \i43/i48/i71  (.A1(\i43/i48/n66 ),
    .A2(\i43/i48/n87 ),
    .B(\i43/i48/n365 ),
    .C(\i43/i48/n368 ),
    .Y(\i43/i48/n440 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i72  (.A(\i43/i48/n514 ),
    .B(\i43/i48/n403 ),
    .Y(\i43/i48/n439 ));
 AND3x1_ASAP7_75t_SL \i43/i48/i73  (.A(\i43/i48/n352 ),
    .B(\i43/i48/n363 ),
    .C(\i43/i48/n348 ),
    .Y(\i43/i48/n438 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i74  (.A(\i43/i48/n377 ),
    .B(\i43/i48/n364 ),
    .Y(\i43/i48/n453 ));
 NOR3xp33_ASAP7_75t_SL \i43/i48/i75  (.A(\i43/i48/n327 ),
    .B(\i43/i48/n361 ),
    .C(\i43/i48/n201 ),
    .Y(\i43/i48/n452 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i76  (.A(\i43/i48/n323 ),
    .B(\i43/i48/n381 ),
    .Y(\i43/i48/n451 ));
 NAND2xp33_ASAP7_75t_SL \i43/i48/i77  (.A(\i43/i48/n368 ),
    .B(\i43/i48/n389 ),
    .Y(\i43/i48/n437 ));
 NAND3xp33_ASAP7_75t_SL \i43/i48/i78  (.A(\i43/i48/n318 ),
    .B(\i43/i48/n355 ),
    .C(\i43/i48/n295 ),
    .Y(\i43/i48/n450 ));
 NAND2xp33_ASAP7_75t_SL \i43/i48/i79  (.A(\i43/i48/n370 ),
    .B(\i43/i48/n391 ),
    .Y(\i43/i48/n436 ));
 NAND4xp25_ASAP7_75t_SL \i43/i48/i8  (.A(\i43/i48/n486 ),
    .B(\i43/i48/n488 ),
    .C(\i43/i48/n475 ),
    .D(\i43/i48/n463 ),
    .Y(\i43/i48/n506 ));
 NAND2xp33_ASAP7_75t_SL \i43/i48/i80  (.A(\i43/i48/n406 ),
    .B(\i43/i48/n414 ),
    .Y(\i43/i48/n432 ));
 NAND4xp25_ASAP7_75t_SL \i43/i48/i81  (.A(\i43/i48/n323 ),
    .B(\i43/i48/n326 ),
    .C(\i43/i48/n294 ),
    .D(\i43/i48/n360 ),
    .Y(\i43/i48/n431 ));
 NAND3xp33_ASAP7_75t_SL \i43/i48/i82  (.A(\i43/i48/n322 ),
    .B(\i43/i48/n291 ),
    .C(\i43/i48/n276 ),
    .Y(\i43/i48/n430 ));
 NAND2xp5_ASAP7_75t_SL \i43/i48/i83  (.A(\i43/i48/n317 ),
    .B(\i43/i48/n385 ),
    .Y(\i43/i48/n429 ));
 NAND5xp2_ASAP7_75t_SL \i43/i48/i84  (.A(\i43/i48/n355 ),
    .B(\i43/i48/n214 ),
    .C(\i43/i48/n339 ),
    .D(\i43/i48/n235 ),
    .E(\i43/i48/n229 ),
    .Y(\i43/i48/n428 ));
 AOI211xp5_ASAP7_75t_SL \i43/i48/i85  (.A1(\i43/i48/n243 ),
    .A2(\i43/i48/n47 ),
    .B(\i43/i48/n284 ),
    .C(\i43/i48/n275 ),
    .Y(\i43/i48/n427 ));
 NOR2xp33_ASAP7_75t_L \i43/i48/i86  (.A(\i43/i48/n376 ),
    .B(\i43/i48/n409 ),
    .Y(\i43/i48/n426 ));
 NAND5xp2_ASAP7_75t_SL \i43/i48/i87  (.A(\i43/i48/n319 ),
    .B(\i43/i48/n367 ),
    .C(\i43/i48/n230 ),
    .D(\i43/i48/n127 ),
    .E(\i43/i48/n110 ),
    .Y(\i43/i48/n425 ));
 NAND4xp25_ASAP7_75t_SL \i43/i48/i88  (.A(\i43/i48/n352 ),
    .B(\i43/i48/n366 ),
    .C(\i43/i48/n345 ),
    .D(\i43/i48/n285 ),
    .Y(\i43/i48/n424 ));
 NOR2xp33_ASAP7_75t_SL \i43/i48/i89  (.A(\i43/i48/n346 ),
    .B(\i43/i48/n373 ),
    .Y(\i43/i48/n423 ));
 NAND4xp25_ASAP7_75t_SL \i43/i48/i9  (.A(\i43/i48/n480 ),
    .B(\i43/i48/n497 ),
    .C(\i43/i48/n494 ),
    .D(\i43/i48/n456 ),
    .Y(\i43/i48/n505 ));
 NOR5xp2_ASAP7_75t_SL \i43/i48/i90  (.A(\i43/i48/n335 ),
    .B(\i43/i48/n338 ),
    .C(\i43/i48/n119 ),
    .D(\i43/i48/n152 ),
    .E(\i43/i48/n102 ),
    .Y(\i43/i48/n422 ));
 AOI221xp5_ASAP7_75t_SL \i43/i48/i91  (.A1(\i43/i48/n258 ),
    .A2(\i43/i48/n55 ),
    .B1(\i43/i48/n155 ),
    .B2(\i43/i48/n256 ),
    .C(\i43/i48/n211 ),
    .Y(\i43/i48/n421 ));
 NOR5xp2_ASAP7_75t_SL \i43/i48/i92  (.A(\i43/i48/n212 ),
    .B(\i43/i48/n270 ),
    .C(\i43/i48/n239 ),
    .D(\i43/i48/n218 ),
    .E(\i43/i48/n177 ),
    .Y(\i43/i48/n420 ));
 NOR5xp2_ASAP7_75t_SL \i43/i48/i93  (.A(\i43/i48/n314 ),
    .B(\i43/i48/n350 ),
    .C(\i43/i48/n340 ),
    .D(\i43/i48/n217 ),
    .E(\i43/i48/n223 ),
    .Y(\i43/i48/n419 ));
 AOI211xp5_ASAP7_75t_SL \i43/i48/i94  (.A1(\i43/i48/n0 ),
    .A2(\i43/i48/n38 ),
    .B(\i43/i48/n297 ),
    .C(\i43/i48/n289 ),
    .Y(\i43/i48/n418 ));
 NOR5xp2_ASAP7_75t_SL \i43/i48/i95  (.A(\i43/i48/n328 ),
    .B(\i43/i48/n274 ),
    .C(\i43/i48/n280 ),
    .D(\i43/i48/n124 ),
    .E(\i43/i48/n174 ),
    .Y(\i43/i48/n417 ));
 NOR2xp67_ASAP7_75t_SL \i43/i48/i96  (.A(\i43/i48/n402 ),
    .B(\i43/i48/n404 ),
    .Y(\i43/i48/n435 ));
 AO211x2_ASAP7_75t_SL \i43/i48/i97  (.A1(\i43/i48/n88 ),
    .A2(\i43/i48/n262 ),
    .B(\i43/i48/n234 ),
    .C(\i43/i48/n313 ),
    .Y(\i43/i48/n434 ));
 AOI21xp5_ASAP7_75t_SL \i43/i48/i98  (.A1(\i43/i48/n33 ),
    .A2(\i43/i48/n73 ),
    .B(\i43/i48/n511 ),
    .Y(\i43/i48/n433 ));
 INVx1_ASAP7_75t_SL \i43/i48/i99  (.A(\i43/i48/n412 ),
    .Y(\i43/i48/n413 ));
 INVxp67_ASAP7_75t_SL \i43/i480  (.A(net73),
    .Y(\i43/n152 ));
 INVxp67_ASAP7_75t_SL \i43/i481  (.A(net84),
    .Y(\i43/n151 ));
 INVxp67_ASAP7_75t_SL \i43/i482  (.A(net93),
    .Y(\i43/n150 ));
 INVxp67_ASAP7_75t_SL \i43/i483  (.A(net57),
    .Y(\i43/n149 ));
 INVxp67_ASAP7_75t_SL \i43/i484  (.A(net92),
    .Y(\i43/n148 ));
 INVxp67_ASAP7_75t_SL \i43/i485  (.A(net53),
    .Y(\i43/n147 ));
 INVxp67_ASAP7_75t_SL \i43/i486  (.A(net97),
    .Y(\i43/n146 ));
 INVxp67_ASAP7_75t_SL \i43/i487  (.A(net38),
    .Y(\i43/n145 ));
 INVxp67_ASAP7_75t_SL \i43/i488  (.A(net108),
    .Y(\i43/n144 ));
 INVxp67_ASAP7_75t_SL \i43/i489  (.A(net120),
    .Y(\i43/n143 ));
 NOR2x1_ASAP7_75t_SL \i43/i49/i0  (.A(\i43/i49/n479 ),
    .B(\i43/i49/n506 ),
    .Y(\i43/n0 [1]));
 AND3x1_ASAP7_75t_SL \i43/i49/i1  (.A(\i43/i49/n502 ),
    .B(\i43/i49/n504 ),
    .C(\i43/i49/n483 ),
    .Y(\i43/n0 [5]));
 NOR4xp75_ASAP7_75t_SL \i43/i49/i10  (.A(\i43/i49/n492 ),
    .B(\i43/i49/n496 ),
    .C(\i43/i49/n474 ),
    .D(\i43/i49/n489 ),
    .Y(\i43/n0 [2]));
 INVx1_ASAP7_75t_SL \i43/i49/i100  (.A(\i43/i49/n409 ),
    .Y(\i43/i49/n410 ));
 INVx1_ASAP7_75t_SL \i43/i49/i101  (.A(\i43/i49/n407 ),
    .Y(\i43/i49/n408 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i102  (.A(\i43/i49/n356 ),
    .B(\i43/i49/n351 ),
    .Y(\i43/i49/n406 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i103  (.A(\i43/i49/n325 ),
    .B(\i43/i49/n321 ),
    .Y(\i43/i49/n405 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i104  (.A(\i43/i49/n369 ),
    .B(\i43/i49/n324 ),
    .Y(\i43/i49/n404 ));
 NAND3xp33_ASAP7_75t_L \i43/i49/i105  (.A(\i43/i49/n267 ),
    .B(\i43/i49/n273 ),
    .C(\i43/i49/n354 ),
    .Y(\i43/i49/n403 ));
 NAND2xp5_ASAP7_75t_L \i43/i49/i106  (.A(\i43/i49/n337 ),
    .B(\i43/i49/n213 ),
    .Y(\i43/i49/n402 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i107  (.A(\i43/i49/n357 ),
    .B(\i43/i49/n331 ),
    .Y(\i43/i49/n401 ));
 NAND5xp2_ASAP7_75t_SL \i43/i49/i108  (.A(\i43/i49/n296 ),
    .B(\i43/i49/n120 ),
    .C(\i43/i49/n181 ),
    .D(\i43/i49/n123 ),
    .E(\i43/i49/n117 ),
    .Y(\i43/i49/n400 ));
 NOR4xp25_ASAP7_75t_SL \i43/i49/i109  (.A(\i43/i49/n279 ),
    .B(\i43/i49/n196 ),
    .C(\i43/i49/n131 ),
    .D(\i43/i49/n225 ),
    .Y(\i43/i49/n399 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i11  (.A(\i43/i49/n509 ),
    .B(\i43/i49/n491 ),
    .Y(\i43/i49/n504 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i110  (.A(\i43/i49/n347 ),
    .B(\i43/i49/n359 ),
    .Y(\i43/i49/n398 ));
 NAND2xp33_ASAP7_75t_SL \i43/i49/i111  (.A(\i43/i49/n320 ),
    .B(\i43/i49/n303 ),
    .Y(\i43/i49/n397 ));
 AOI221xp5_ASAP7_75t_SL \i43/i49/i112  (.A1(\i43/i49/n109 ),
    .A2(\i43/i49/n95 ),
    .B1(\i43/i49/n115 ),
    .B2(\i43/i49/n47 ),
    .C(\i43/i49/n215 ),
    .Y(\i43/i49/n416 ));
 NAND5xp2_ASAP7_75t_SL \i43/i49/i113  (.A(\i43/i49/n277 ),
    .B(\i43/i49/n205 ),
    .C(\i43/i49/n210 ),
    .D(\i43/i49/n181 ),
    .E(\i43/i49/n122 ),
    .Y(\i43/i49/n396 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i114  (.A(\i43/i49/n293 ),
    .B(\i43/i49/n369 ),
    .Y(\i43/i49/n395 ));
 OAI221xp5_ASAP7_75t_SL \i43/i49/i115  (.A1(\i43/i49/n156 ),
    .A2(\i43/i49/n54 ),
    .B1(\i43/i49/n157 ),
    .B2(\i43/i49/n39 ),
    .C(\i43/i49/n336 ),
    .Y(\i43/i49/n394 ));
 NOR2xp33_ASAP7_75t_L \i43/i49/i116  (.A(\i43/i49/n290 ),
    .B(\i43/i49/n356 ),
    .Y(\i43/i49/n415 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i117  (.A(\i43/i49/n287 ),
    .B(\i43/i49/n319 ),
    .Y(\i43/i49/n414 ));
 NOR3xp33_ASAP7_75t_SL \i43/i49/i118  (.A(\i43/i49/n217 ),
    .B(\i43/i49/n226 ),
    .C(\i43/i49/n195 ),
    .Y(\i43/i49/n412 ));
 NAND3xp33_ASAP7_75t_SL \i43/i49/i119  (.A(\i43/i49/n332 ),
    .B(\i43/i49/n283 ),
    .C(\i43/i49/n238 ),
    .Y(\i43/i49/n411 ));
 NAND3xp33_ASAP7_75t_SL \i43/i49/i12  (.A(\i43/i49/n477 ),
    .B(\i43/i49/n482 ),
    .C(\i43/i49/n416 ),
    .Y(\i43/i49/n503 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i120  (.A(\i43/i49/n214 ),
    .B(\i43/i49/n298 ),
    .Y(\i43/i49/n409 ));
 NOR3xp33_ASAP7_75t_SL \i43/i49/i121  (.A(\i43/i49/n286 ),
    .B(\i43/i49/n231 ),
    .C(\i43/i49/n270 ),
    .Y(\i43/i49/n407 ));
 INVx1_ASAP7_75t_SL \i43/i49/i122  (.A(\i43/i49/n514 ),
    .Y(\i43/i49/n387 ));
 OAI21xp33_ASAP7_75t_SL \i43/i49/i123  (.A1(\i43/i49/n76 ),
    .A2(\i43/i49/n45 ),
    .B(\i43/i49/n367 ),
    .Y(\i43/i49/n386 ));
 NOR3xp33_ASAP7_75t_SL \i43/i49/i124  (.A(\i43/i49/n327 ),
    .B(\i43/i49/n191 ),
    .C(\i43/i49/n231 ),
    .Y(\i43/i49/n385 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i125  (.A1(\i43/i49/n87 ),
    .A2(\i43/i49/n50 ),
    .B(\i43/i49/n354 ),
    .Y(\i43/i49/n393 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i126  (.A1(\i43/i49/n41 ),
    .A2(\i43/i49/n268 ),
    .B(\i43/i49/n263 ),
    .Y(\i43/i49/n384 ));
 NAND4xp25_ASAP7_75t_SL \i43/i49/i127  (.A(\i43/i49/n244 ),
    .B(\i43/i49/n145 ),
    .C(\i43/i49/n96 ),
    .D(\i43/i49/n99 ),
    .Y(\i43/i49/n383 ));
 NAND5xp2_ASAP7_75t_SL \i43/i49/i128  (.A(\i43/i49/n208 ),
    .B(\i43/i49/n120 ),
    .C(\i43/i49/n164 ),
    .D(\i43/i49/n184 ),
    .E(\i43/i49/n140 ),
    .Y(\i43/i49/n382 ));
 AOI211xp5_ASAP7_75t_SL \i43/i49/i129  (.A1(\i43/i49/n41 ),
    .A2(\i43/i49/n62 ),
    .B(\i43/i49/n282 ),
    .C(\i43/i49/n281 ),
    .Y(\i43/i49/n381 ));
 NOR3xp33_ASAP7_75t_SL \i43/i49/i13  (.A(\i43/i49/n508 ),
    .B(\i43/i49/n478 ),
    .C(\i43/i49/n455 ),
    .Y(\i43/i49/n502 ));
 NOR3xp33_ASAP7_75t_SL \i43/i49/i130  (.A(\i43/i49/n292 ),
    .B(\i43/i49/n206 ),
    .C(\i43/i49/n221 ),
    .Y(\i43/i49/n380 ));
 NOR2xp33_ASAP7_75t_L \i43/i49/i131  (.A(\i43/i49/n334 ),
    .B(\i43/i49/n315 ),
    .Y(\i43/i49/n379 ));
 OAI221xp5_ASAP7_75t_SL \i43/i49/i132  (.A1(\i43/i49/n269 ),
    .A2(\i43/i49/n75 ),
    .B1(\i43/i49/n173 ),
    .B2(\i43/i49/n72 ),
    .C(\i43/i49/n89 ),
    .Y(\i43/i49/n378 ));
 NAND5xp2_ASAP7_75t_SL \i43/i49/i133  (.A(\i43/i49/n246 ),
    .B(\i43/i49/n175 ),
    .C(\i43/i49/n105 ),
    .D(\i43/i49/n113 ),
    .E(\i43/i49/n144 ),
    .Y(\i43/i49/n377 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i134  (.A1(\i43/i49/n45 ),
    .A2(\i43/i49/n40 ),
    .B(\i43/i49/n357 ),
    .Y(\i43/i49/n376 ));
 NOR4xp25_ASAP7_75t_SL \i43/i49/i135  (.A(\i43/i49/n333 ),
    .B(\i43/i49/n266 ),
    .C(\i43/i49/n97 ),
    .D(\i43/i49/n98 ),
    .Y(\i43/i49/n375 ));
 OAI211xp5_ASAP7_75t_SL \i43/i49/i136  (.A1(\i43/i49/n40 ),
    .A2(\i43/i49/n259 ),
    .B(\i43/i49/n179 ),
    .C(\i43/i49/n167 ),
    .Y(\i43/i49/n374 ));
 NAND5xp2_ASAP7_75t_SL \i43/i49/i137  (.A(\i43/i49/n257 ),
    .B(\i43/i49/n242 ),
    .C(\i43/i49/n118 ),
    .D(\i43/i49/n180 ),
    .E(\i43/i49/n185 ),
    .Y(\i43/i49/n373 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i138  (.A(\i43/i49/n330 ),
    .B(\i43/i49/n301 ),
    .Y(\i43/i49/n372 ));
 OAI221xp5_ASAP7_75t_SL \i43/i49/i139  (.A1(\i43/i49/n260 ),
    .A2(\i43/i49/n54 ),
    .B1(\i43/i49/n52 ),
    .B2(\i43/i49/n87 ),
    .C(\i43/i49/n222 ),
    .Y(\i43/i49/n371 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i14  (.A(\i43/i49/n493 ),
    .B(\i43/i49/n481 ),
    .Y(\i43/i49/n501 ));
 NOR3xp33_ASAP7_75t_SL \i43/i49/i140  (.A(\i43/i49/n307 ),
    .B(\i43/i49/n274 ),
    .C(\i43/i49/n272 ),
    .Y(\i43/i49/n392 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i141  (.A(\i43/i49/n240 ),
    .B(\i43/i49/n358 ),
    .Y(\i43/i49/n391 ));
 OA211x2_ASAP7_75t_SL \i43/i49/i142  (.A1(\i43/i49/n92 ),
    .A2(\i43/i49/n54 ),
    .B(\i43/i49/n366 ),
    .C(\i43/i49/n146 ),
    .Y(\i43/i49/n390 ));
 NOR2xp33_ASAP7_75t_L \i43/i49/i143  (.A(\i43/i49/n190 ),
    .B(\i43/i49/n316 ),
    .Y(\i43/i49/n389 ));
 NOR2xp33_ASAP7_75t_L \i43/i49/i144  (.A(\i43/i49/n200 ),
    .B(\i43/i49/n362 ),
    .Y(\i43/i49/n388 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i145  (.A(\i43/i49/n364 ),
    .Y(\i43/i49/n365 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i146  (.A(\i43/i49/n362 ),
    .Y(\i43/i49/n363 ));
 INVx1_ASAP7_75t_SL \i43/i49/i147  (.A(\i43/i49/n360 ),
    .Y(\i43/i49/n361 ));
 INVx1_ASAP7_75t_SL \i43/i49/i148  (.A(\i43/i49/n358 ),
    .Y(\i43/i49/n359 ));
 INVx1_ASAP7_75t_SL \i43/i49/i149  (.A(\i43/i49/n512 ),
    .Y(\i43/i49/n352 ));
 NAND3xp33_ASAP7_75t_SL \i43/i49/i15  (.A(\i43/i49/n466 ),
    .B(\i43/i49/n476 ),
    .C(\i43/i49/n454 ),
    .Y(\i43/i49/n500 ));
 NAND2xp33_ASAP7_75t_L \i43/i49/i150  (.A(\i43/i49/n214 ),
    .B(\i43/i49/n271 ),
    .Y(\i43/i49/n351 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i151  (.A(\i43/i49/n130 ),
    .B(\i43/i49/n220 ),
    .Y(\i43/i49/n350 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i152  (.A(\i43/i49/n192 ),
    .B(\i43/i49/n212 ),
    .Y(\i43/i49/n349 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i49/i153  (.A1(\i43/i49/n34 ),
    .A2(\i43/i49/n65 ),
    .B(\i43/i49/n33 ),
    .C(\i43/i49/n227 ),
    .Y(\i43/i49/n348 ));
 OAI31xp33_ASAP7_75t_SL \i43/i49/i154  (.A1(\i43/i49/n65 ),
    .A2(\i43/i49/n41 ),
    .A3(\i43/i49/n55 ),
    .B(\i43/i49/n79 ),
    .Y(\i43/i49/n347 ));
 NAND3xp33_ASAP7_75t_SL \i43/i49/i155  (.A(\i43/i49/n213 ),
    .B(\i43/i49/n183 ),
    .C(\i43/i49/n128 ),
    .Y(\i43/i49/n346 ));
 AOI21xp5_ASAP7_75t_SL \i43/i49/i156  (.A1(\i43/i49/n38 ),
    .A2(\i43/i49/n74 ),
    .B(\i43/i49/n1 ),
    .Y(\i43/i49/n345 ));
 AOI211xp5_ASAP7_75t_SL \i43/i49/i157  (.A1(\i43/i49/n57 ),
    .A2(\i43/i49/n71 ),
    .B(\i43/i49/n182 ),
    .C(\i43/i49/n121 ),
    .Y(\i43/i49/n370 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i158  (.A1(\i43/i49/n94 ),
    .A2(\i43/i49/n58 ),
    .B(\i43/i49/n216 ),
    .Y(\i43/i49/n344 ));
 OAI31xp33_ASAP7_75t_SL \i43/i49/i159  (.A1(\i43/i49/n47 ),
    .A2(\i43/i49/n95 ),
    .A3(\i43/i49/n51 ),
    .B(\i43/i49/n69 ),
    .Y(\i43/i49/n343 ));
 NOR2xp33_ASAP7_75t_L \i43/i49/i16  (.A(\i43/i49/n465 ),
    .B(\i43/i49/n461 ),
    .Y(\i43/i49/n497 ));
 AO21x1_ASAP7_75t_SL \i43/i49/i160  (.A1(\i43/i49/n67 ),
    .A2(\i43/i49/n150 ),
    .B(\i43/i49/n280 ),
    .Y(\i43/i49/n342 ));
 AO21x1_ASAP7_75t_SL \i43/i49/i161  (.A1(\i43/i49/n148 ),
    .A2(\i43/i49/n173 ),
    .B(\i43/i49/n76 ),
    .Y(\i43/i49/n341 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i43/i49/i162  (.A1(\i43/i49/n70 ),
    .A2(\i43/i49/n78 ),
    .B(\i43/i49/n52 ),
    .C(\i43/i49/n197 ),
    .Y(\i43/i49/n340 ));
 AOI21xp5_ASAP7_75t_SL \i43/i49/i163  (.A1(\i43/i49/n44 ),
    .A2(\i43/i49/n67 ),
    .B(\i43/i49/n219 ),
    .Y(\i43/i49/n339 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i43/i49/i164  (.A1(\i43/i49/n42 ),
    .A2(\i43/i49/n35 ),
    .B(\i43/i49/n87 ),
    .C(\i43/i49/n117 ),
    .Y(\i43/i49/n338 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i165  (.A(\i43/i49/n249 ),
    .B(\i43/i49/n236 ),
    .Y(\i43/i49/n337 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i49/i166  (.A1(\i43/i49/n77 ),
    .A2(\i43/i49/n51 ),
    .B(\i43/i49/n33 ),
    .C(\i43/i49/n132 ),
    .Y(\i43/i49/n336 ));
 NAND3xp33_ASAP7_75t_SL \i43/i49/i167  (.A(\i43/i49/n232 ),
    .B(\i43/i49/n172 ),
    .C(\i43/i49/n137 ),
    .Y(\i43/i49/n335 ));
 OAI221xp5_ASAP7_75t_SL \i43/i49/i168  (.A1(\i43/i49/n75 ),
    .A2(\i43/i49/n56 ),
    .B1(\i43/i49/n49 ),
    .B2(\i43/i49/n68 ),
    .C(\i43/i49/n134 ),
    .Y(\i43/i49/n334 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i169  (.A1(\i43/i49/n78 ),
    .A2(\i43/i49/n136 ),
    .B(\i43/i49/n237 ),
    .Y(\i43/i49/n333 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i17  (.A(\i43/i49/n468 ),
    .B(\i43/i49/n476 ),
    .Y(\i43/i49/n496 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i170  (.A(\i43/i49/n233 ),
    .B(\i43/i49/n209 ),
    .Y(\i43/i49/n332 ));
 AOI221xp5_ASAP7_75t_SL \i43/i49/i171  (.A1(\i43/i49/n34 ),
    .A2(\i43/i49/n79 ),
    .B1(\i43/i49/n67 ),
    .B2(\i43/i49/n83 ),
    .C(\i43/i49/n236 ),
    .Y(\i43/i49/n331 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i172  (.A1(\i43/i49/n59 ),
    .A2(\i43/i49/n154 ),
    .B(\i43/i49/n77 ),
    .Y(\i43/i49/n330 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i49/i173  (.A1(\i43/i49/n62 ),
    .A2(\i43/i49/n44 ),
    .B(\i43/i49/n57 ),
    .C(\i43/i49/n125 ),
    .Y(\i43/i49/n329 ));
 OAI221xp5_ASAP7_75t_SL \i43/i49/i174  (.A1(\i43/i49/n46 ),
    .A2(\i43/i49/n87 ),
    .B1(\i43/i49/n52 ),
    .B2(\i43/i49/n80 ),
    .C(\i43/i49/n162 ),
    .Y(\i43/i49/n328 ));
 AOI21xp5_ASAP7_75t_SL \i43/i49/i175  (.A1(\i43/i49/n95 ),
    .A2(\i43/i49/n62 ),
    .B(\i43/i49/n1 ),
    .Y(\i43/i49/n369 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i176  (.A(\i43/i49/n219 ),
    .B(\i43/i49/n251 ),
    .Y(\i43/i49/n368 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i177  (.A(\i43/i49/n253 ),
    .B(\i43/i49/n0 ),
    .Y(\i43/i49/n367 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i178  (.A(\i43/i49/n225 ),
    .B(\i43/i49/n194 ),
    .Y(\i43/i49/n366 ));
 OAI211xp5_ASAP7_75t_SL \i43/i49/i179  (.A1(\i43/i49/n63 ),
    .A2(\i43/i49/n46 ),
    .B(\i43/i49/n176 ),
    .C(\i43/i49/n186 ),
    .Y(\i43/i49/n364 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i18  (.A(\i43/i49/n473 ),
    .B(\i43/i49/n464 ),
    .Y(\i43/i49/n495 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i180  (.A(\i43/i49/n120 ),
    .B(\i43/i49/n245 ),
    .Y(\i43/i49/n362 ));
 AOI222xp33_ASAP7_75t_SL \i43/i49/i181  (.A1(\i43/i49/n85 ),
    .A2(\i43/i49/n41 ),
    .B1(\i43/i49/n59 ),
    .B2(\i43/i49/n38 ),
    .C1(\i43/i49/n69 ),
    .C2(\i43/i49/n47 ),
    .Y(\i43/i49/n360 ));
 OAI221xp5_ASAP7_75t_SL \i43/i49/i182  (.A1(\i43/i49/n45 ),
    .A2(\i43/i49/n35 ),
    .B1(\i43/i49/n37 ),
    .B2(\i43/i49/n52 ),
    .C(\i43/i49/n179 ),
    .Y(\i43/i49/n358 ));
 AOI222xp33_ASAP7_75t_SL \i43/i49/i183  (.A1(\i43/i49/n34 ),
    .A2(\i43/i49/n90 ),
    .B1(\i43/i49/n33 ),
    .B2(\i43/i49/n67 ),
    .C1(\i43/i49/n83 ),
    .C2(\i43/i49/n73 ),
    .Y(\i43/i49/n357 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i184  (.A1(\i43/i49/n39 ),
    .A2(\i43/i49/n91 ),
    .B(\i43/i49/n237 ),
    .Y(\i43/i49/n356 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i185  (.A(\i43/i49/n204 ),
    .B(\i43/i49/n227 ),
    .Y(\i43/i49/n355 ));
 NOR2xp67_ASAP7_75t_SL \i43/i49/i186  (.A(\i43/i49/n255 ),
    .B(\i43/i49/n279 ),
    .Y(\i43/i49/n354 ));
 NOR2x1_ASAP7_75t_SL \i43/i49/i187  (.A(\i43/i49/n141 ),
    .B(\i43/i49/n278 ),
    .Y(\i43/i49/n353 ));
 INVxp33_ASAP7_75t_SL \i43/i49/i188  (.A(\i43/i49/n324 ),
    .Y(\i43/i49/n325 ));
 INVx1_ASAP7_75t_SL \i43/i49/i189  (.A(\i43/i49/n321 ),
    .Y(\i43/i49/n322 ));
 NOR4xp25_ASAP7_75t_SL \i43/i49/i19  (.A(\i43/i49/n429 ),
    .B(\i43/i49/n395 ),
    .C(\i43/i49/n372 ),
    .D(\i43/i49/n371 ),
    .Y(\i43/i49/n494 ));
 INVx1_ASAP7_75t_SL \i43/i49/i190  (.A(\i43/i49/n316 ),
    .Y(\i43/i49/n317 ));
 OAI211xp5_ASAP7_75t_SL \i43/i49/i191  (.A1(\i43/i49/n40 ),
    .A2(\i43/i49/n70 ),
    .B(\i43/i49/n188 ),
    .C(\i43/i49/n187 ),
    .Y(\i43/i49/n315 ));
 AO21x1_ASAP7_75t_SL \i43/i49/i192  (.A1(\i43/i49/n67 ),
    .A2(\i43/i49/n0 ),
    .B(\i43/i49/n224 ),
    .Y(\i43/i49/n314 ));
 OAI221xp5_ASAP7_75t_SL \i43/i49/i193  (.A1(\i43/i49/n72 ),
    .A2(\i43/i49/n70 ),
    .B1(\i43/i49/n42 ),
    .B2(\i43/i49/n63 ),
    .C(\i43/i49/n118 ),
    .Y(\i43/i49/n313 ));
 OA211x2_ASAP7_75t_SL \i43/i49/i194  (.A1(\i43/i49/n37 ),
    .A2(\i43/i49/n136 ),
    .B(\i43/i49/n100 ),
    .C(\i43/i49/n159 ),
    .Y(\i43/i49/n312 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i49/i195  (.A1(\i43/i49/n47 ),
    .A2(\i43/i49/n34 ),
    .B(\i43/i49/n85 ),
    .C(\i43/i49/n241 ),
    .Y(\i43/i49/n311 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i196  (.A(\i43/i49/n265 ),
    .B(\i43/i49/n266 ),
    .Y(\i43/i49/n310 ));
 OAI31xp33_ASAP7_75t_SL \i43/i49/i197  (.A1(\i43/i49/n57 ),
    .A2(\i43/i49/n53 ),
    .A3(\i43/i49/n88 ),
    .B(\i43/i49/n62 ),
    .Y(\i43/i49/n309 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i198  (.A1(\i43/i49/n51 ),
    .A2(\i43/i49/n166 ),
    .B(\i43/i49/n71 ),
    .Y(\i43/i49/n308 ));
 OAI211xp5_ASAP7_75t_SL \i43/i49/i199  (.A1(\i43/i49/n52 ),
    .A2(\i43/i49/n91 ),
    .B(\i43/i49/n138 ),
    .C(\i43/i49/n139 ),
    .Y(\i43/i49/n307 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i2  (.A(\i43/i49/n507 ),
    .B(\i43/i49/n503 ),
    .Y(\i43/n0 [6]));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i20  (.A(\i43/i49/n452 ),
    .B(\i43/i49/n459 ),
    .Y(\i43/i49/n493 ));
 OAI221xp5_ASAP7_75t_SL \i43/i49/i200  (.A1(\i43/i49/n94 ),
    .A2(\i43/i49/n87 ),
    .B1(\i43/i49/n78 ),
    .B2(\i43/i49/n54 ),
    .C(\i43/i49/n137 ),
    .Y(\i43/i49/n306 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i201  (.A1(\i43/i49/n56 ),
    .A2(\i43/i49/n156 ),
    .B1(\i43/i49/n63 ),
    .B2(\i43/i49/n72 ),
    .Y(\i43/i49/n305 ));
 OAI211xp5_ASAP7_75t_SL \i43/i49/i202  (.A1(\i43/i49/n82 ),
    .A2(\i43/i49/n72 ),
    .B(\i43/i49/n264 ),
    .C(\i43/i49/n178 ),
    .Y(\i43/i49/n304 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i49/i203  (.A1(\i43/i49/n51 ),
    .A2(\i43/i49/n53 ),
    .B(\i43/i49/n85 ),
    .C(\i43/i49/n203 ),
    .Y(\i43/i49/n303 ));
 AOI221xp5_ASAP7_75t_SL \i43/i49/i204  (.A1(\i43/i49/n44 ),
    .A2(\i43/i49/n38 ),
    .B1(\i43/i49/n104 ),
    .B2(\i43/i49/n71 ),
    .C(\i43/i49/n161 ),
    .Y(\i43/i49/n302 ));
 NOR3xp33_ASAP7_75t_SL \i43/i49/i205  (.A(\i43/i49/n250 ),
    .B(\i43/i49/n170 ),
    .C(\i43/i49/n101 ),
    .Y(\i43/i49/n301 ));
 AOI21xp5_ASAP7_75t_SL \i43/i49/i206  (.A1(\i43/i49/n150 ),
    .A2(\i43/i49/n73 ),
    .B(\i43/i49/n261 ),
    .Y(\i43/i49/n300 ));
 OAI211xp5_ASAP7_75t_SL \i43/i49/i207  (.A1(\i43/i49/n89 ),
    .A2(\i43/i49/n157 ),
    .B(\i43/i49/n126 ),
    .C(\i43/i49/n135 ),
    .Y(\i43/i49/n299 ));
 AOI222xp33_ASAP7_75t_SL \i43/i49/i208  (.A1(\i43/i49/n112 ),
    .A2(\i43/i49/n67 ),
    .B1(\i43/i49/n65 ),
    .B2(\i43/i49/n79 ),
    .C1(\i43/i49/n59 ),
    .C2(\i43/i49/n48 ),
    .Y(\i43/i49/n298 ));
 NAND4xp25_ASAP7_75t_SL \i43/i49/i209  (.A(\i43/i49/n133 ),
    .B(\i43/i49/n164 ),
    .C(\i43/i49/n171 ),
    .D(\i43/i49/n111 ),
    .Y(\i43/i49/n297 ));
 NAND2x1_ASAP7_75t_SL \i43/i49/i21  (.A(\i43/i49/n458 ),
    .B(\i43/i49/n469 ),
    .Y(\i43/i49/n492 ));
 AOI221xp5_ASAP7_75t_SL \i43/i49/i210  (.A1(\i43/i49/n48 ),
    .A2(\i43/i49/n81 ),
    .B1(\i43/i49/n41 ),
    .B2(\i43/i49/n85 ),
    .C(\i43/i49/n207 ),
    .Y(\i43/i49/n296 ));
 AOI222xp33_ASAP7_75t_SL \i43/i49/i211  (.A1(\i43/i49/n67 ),
    .A2(\i43/i49/n60 ),
    .B1(\i43/i49/n88 ),
    .B2(\i43/i49/n85 ),
    .C1(\i43/i49/n95 ),
    .C2(\i43/i49/n71 ),
    .Y(\i43/i49/n295 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i43/i49/i212  (.A1(\i43/i49/n44 ),
    .A2(\i43/i49/n36 ),
    .B(\i43/i49/n48 ),
    .C(\i43/i49/n215 ),
    .Y(\i43/i49/n294 ));
 AOI22xp33_ASAP7_75t_SL \i43/i49/i213  (.A1(\i43/i49/n65 ),
    .A2(\i43/i49/n0 ),
    .B1(\i43/i49/n33 ),
    .B2(\i43/i49/n106 ),
    .Y(\i43/i49/n293 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i214  (.A1(\i43/i49/n75 ),
    .A2(\i43/i49/n103 ),
    .B1(\i43/i49/n46 ),
    .B2(\i43/i49/n37 ),
    .Y(\i43/i49/n292 ));
 AOI211xp5_ASAP7_75t_SL \i43/i49/i215  (.A1(\i43/i49/n67 ),
    .A2(\i43/i49/n79 ),
    .B(\i43/i49/n254 ),
    .C(\i43/i49/n170 ),
    .Y(\i43/i49/n291 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i216  (.A1(\i43/i49/n87 ),
    .A2(\i43/i49/n114 ),
    .B1(\i43/i49/n76 ),
    .B2(\i43/i49/n37 ),
    .Y(\i43/i49/n290 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i43/i49/i217  (.A1(\i43/i49/n42 ),
    .A2(\i43/i49/n49 ),
    .B(\i43/i49/n80 ),
    .C(\i43/i49/n252 ),
    .Y(\i43/i49/n289 ));
 AOI22xp5_ASAP7_75t_SL \i43/i49/i218  (.A1(\i43/i49/n83 ),
    .A2(\i43/i49/n143 ),
    .B1(\i43/i49/n71 ),
    .B2(\i43/i49/n38 ),
    .Y(\i43/i49/n288 ));
 AOI222xp33_ASAP7_75t_SL \i43/i49/i219  (.A1(\i43/i49/n79 ),
    .A2(\i43/i49/n48 ),
    .B1(\i43/i49/n69 ),
    .B2(\i43/i49/n38 ),
    .C1(\i43/i49/n74 ),
    .C2(\i43/i49/n67 ),
    .Y(\i43/i49/n287 ));
 NAND4xp25_ASAP7_75t_SL \i43/i49/i22  (.A(\i43/i49/n423 ),
    .B(\i43/i49/n427 ),
    .C(\i43/i49/n388 ),
    .D(\i43/i49/n443 ),
    .Y(\i43/i49/n491 ));
 OAI221xp5_ASAP7_75t_SL \i43/i49/i220  (.A1(\i43/i49/n35 ),
    .A2(\i43/i49/n80 ),
    .B1(\i43/i49/n68 ),
    .B2(\i43/i49/n76 ),
    .C(\i43/i49/n116 ),
    .Y(\i43/i49/n286 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i221  (.A(\i43/i49/n281 ),
    .B(\i43/i49/n282 ),
    .Y(\i43/i49/n285 ));
 AO21x1_ASAP7_75t_L \i43/i49/i222  (.A1(\i43/i49/n41 ),
    .A2(\i43/i49/n163 ),
    .B(\i43/i49/n198 ),
    .Y(\i43/i49/n327 ));
 AOI21xp5_ASAP7_75t_SL \i43/i49/i223  (.A1(\i43/i49/n154 ),
    .A2(\i43/i49/n88 ),
    .B(\i43/i49/n202 ),
    .Y(\i43/i49/n326 ));
 OA211x2_ASAP7_75t_SL \i43/i49/i224  (.A1(\i43/i49/n54 ),
    .A2(\i43/i49/n142 ),
    .B(\i43/i49/n128 ),
    .C(\i43/i49/n162 ),
    .Y(\i43/i49/n324 ));
 AOI22xp5_ASAP7_75t_SL \i43/i49/i225  (.A1(\i43/i49/n41 ),
    .A2(\i43/i49/n147 ),
    .B1(\i43/i49/n60 ),
    .B2(\i43/i49/n77 ),
    .Y(\i43/i49/n323 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i226  (.A(\i43/i49/n283 ),
    .B(\i43/i49/n238 ),
    .Y(\i43/i49/n284 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i227  (.A1(\i43/i49/n80 ),
    .A2(\i43/i49/n165 ),
    .B1(\i43/i49/n84 ),
    .B2(\i43/i49/n64 ),
    .Y(\i43/i49/n321 ));
 AOI21xp5_ASAP7_75t_SL \i43/i49/i228  (.A1(\i43/i49/n48 ),
    .A2(\i43/i49/n71 ),
    .B(\i43/i49/n218 ),
    .Y(\i43/i49/n320 ));
 AOI222xp33_ASAP7_75t_SL \i43/i49/i229  (.A1(\i43/i49/n43 ),
    .A2(\i43/i49/n59 ),
    .B1(\i43/i49/n73 ),
    .B2(\i43/i49/n85 ),
    .C1(\i43/i49/n34 ),
    .C2(\i43/i49/n71 ),
    .Y(\i43/i49/n319 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i23  (.A(\i43/i49/n470 ),
    .B(\i43/i49/n474 ),
    .Y(\i43/i49/n490 ));
 O2A1O1Ixp33_ASAP7_75t_L \i43/i49/i230  (.A1(\i43/i49/n41 ),
    .A2(\i43/i49/n48 ),
    .B(\i43/i49/n83 ),
    .C(\i43/i49/n224 ),
    .Y(\i43/i49/n318 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i231  (.A(\i43/i49/n108 ),
    .B(\i43/i49/n273 ),
    .Y(\i43/i49/n316 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i232  (.A(\i43/i49/n275 ),
    .Y(\i43/i49/n276 ));
 INVx1_ASAP7_75t_SL \i43/i49/i233  (.A(\i43/i49/n271 ),
    .Y(\i43/i49/n272 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i234  (.A(\i43/i49/n268 ),
    .Y(\i43/i49/n269 ));
 OAI21xp33_ASAP7_75t_SL \i43/i49/i235  (.A1(\i43/i49/n75 ),
    .A2(\i43/i49/n52 ),
    .B(\i43/i49/n123 ),
    .Y(\i43/i49/n265 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i236  (.A(\i43/i49/n125 ),
    .B(\i43/i49/n152 ),
    .Y(\i43/i49/n264 ));
 NAND2xp33_ASAP7_75t_SL \i43/i49/i237  (.A(\i43/i49/n82 ),
    .B(\i43/i49/n127 ),
    .Y(\i43/i49/n263 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i238  (.A(\i43/i49/n75 ),
    .B(\i43/i49/n157 ),
    .Y(\i43/i49/n262 ));
 NAND2xp33_ASAP7_75t_SL \i43/i49/i239  (.A(\i43/i49/n184 ),
    .B(\i43/i49/n126 ),
    .Y(\i43/i49/n261 ));
 NOR2x1_ASAP7_75t_SL \i43/i49/i24  (.A(\i43/i49/n445 ),
    .B(\i43/i49/n465 ),
    .Y(\i43/i49/n499 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i240  (.A(\i43/i49/n60 ),
    .B(\i43/i49/n147 ),
    .Y(\i43/i49/n260 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i241  (.A(\i43/i49/n55 ),
    .B(\i43/i49/n147 ),
    .Y(\i43/i49/n283 ));
 NOR3xp33_ASAP7_75t_SL \i43/i49/i242  (.A(\i43/i49/n71 ),
    .B(\i43/i49/n33 ),
    .C(\i43/i49/n81 ),
    .Y(\i43/i49/n259 ));
 NAND2xp33_ASAP7_75t_L \i43/i49/i243  (.A(\i43/i49/n149 ),
    .B(\i43/i49/n32 ),
    .Y(\i43/i49/n258 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i244  (.A1(\i43/i49/n79 ),
    .A2(\i43/i49/n33 ),
    .B(\i43/i49/n43 ),
    .Y(\i43/i49/n257 ));
 NAND2xp33_ASAP7_75t_SL \i43/i49/i245  (.A(\i43/i49/n42 ),
    .B(\i43/i49/n134 ),
    .Y(\i43/i49/n256 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i246  (.A1(\i43/i49/n87 ),
    .A2(\i43/i49/n64 ),
    .B(\i43/i49/n172 ),
    .Y(\i43/i49/n255 ));
 OAI21xp33_ASAP7_75t_SL \i43/i49/i247  (.A1(\i43/i49/n35 ),
    .A2(\i43/i49/n87 ),
    .B(\i43/i49/n159 ),
    .Y(\i43/i49/n254 ));
 OAI21xp33_ASAP7_75t_SL \i43/i49/i248  (.A1(\i43/i49/n84 ),
    .A2(\i43/i49/n42 ),
    .B(\i43/i49/n52 ),
    .Y(\i43/i49/n253 ));
 OAI21xp33_ASAP7_75t_SL \i43/i49/i249  (.A1(\i43/i49/n95 ),
    .A2(\i43/i49/n53 ),
    .B(\i43/i49/n163 ),
    .Y(\i43/i49/n252 ));
 NOR3xp33_ASAP7_75t_SL \i43/i49/i25  (.A(\i43/i49/n447 ),
    .B(\i43/i49/n434 ),
    .C(\i43/i49/n393 ),
    .Y(\i43/i49/n498 ));
 OAI21xp33_ASAP7_75t_SL \i43/i49/i250  (.A1(\i43/i49/n66 ),
    .A2(\i43/i49/n80 ),
    .B(\i43/i49/n158 ),
    .Y(\i43/i49/n251 ));
 AOI21xp33_ASAP7_75t_SL \i43/i49/i251  (.A1(\i43/i49/n91 ),
    .A2(\i43/i49/n87 ),
    .B(\i43/i49/n49 ),
    .Y(\i43/i49/n250 ));
 OAI21xp33_ASAP7_75t_SL \i43/i49/i252  (.A1(\i43/i49/n58 ),
    .A2(\i43/i49/n35 ),
    .B(\i43/i49/n180 ),
    .Y(\i43/i49/n249 ));
 OAI21xp33_ASAP7_75t_SL \i43/i49/i253  (.A1(\i43/i49/n82 ),
    .A2(\i43/i49/n35 ),
    .B(\i43/i49/n158 ),
    .Y(\i43/i49/n248 ));
 AOI21xp5_ASAP7_75t_SL \i43/i49/i254  (.A1(\i43/i49/n64 ),
    .A2(\i43/i49/n42 ),
    .B(\i43/i49/n91 ),
    .Y(\i43/i49/n282 ));
 AOI21xp5_ASAP7_75t_SL \i43/i49/i255  (.A1(\i43/i49/n83 ),
    .A2(\i43/i49/n65 ),
    .B(\i43/i49/n129 ),
    .Y(\i43/i49/n247 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i256  (.A1(\i43/i49/n74 ),
    .A2(\i43/i49/n86 ),
    .B(\i43/i49/n55 ),
    .Y(\i43/i49/n246 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i257  (.A1(\i43/i49/n77 ),
    .A2(\i43/i49/n34 ),
    .B(\i43/i49/n79 ),
    .Y(\i43/i49/n245 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i258  (.A1(\i43/i49/n66 ),
    .A2(\i43/i49/n84 ),
    .B(\i43/i49/n178 ),
    .Y(\i43/i49/n281 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i259  (.A1(\i43/i49/n81 ),
    .A2(\i43/i49/n62 ),
    .B(\i43/i49/n65 ),
    .Y(\i43/i49/n244 ));
 NAND3xp33_ASAP7_75t_SL \i43/i49/i26  (.A(\i43/i49/n438 ),
    .B(\i43/i49/n440 ),
    .C(\i43/i49/n439 ),
    .Y(\i43/i49/n489 ));
 NAND3xp33_ASAP7_75t_L \i43/i49/i260  (.A(\i43/i49/n37 ),
    .B(\i43/i49/n87 ),
    .C(\i43/i49/n32 ),
    .Y(\i43/i49/n243 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i261  (.A1(\i43/i49/n90 ),
    .A2(\i43/i49/n69 ),
    .B(\i43/i49/n65 ),
    .Y(\i43/i49/n242 ));
 AOI21xp33_ASAP7_75t_SL \i43/i49/i262  (.A1(\i43/i49/n66 ),
    .A2(\i43/i49/n56 ),
    .B(\i43/i49/n75 ),
    .Y(\i43/i49/n241 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i263  (.A1(\i43/i49/n91 ),
    .A2(\i43/i49/n72 ),
    .B(\i43/i49/n185 ),
    .Y(\i43/i49/n240 ));
 OAI21xp33_ASAP7_75t_SL \i43/i49/i264  (.A1(\i43/i49/n80 ),
    .A2(\i43/i49/n54 ),
    .B(\i43/i49/n160 ),
    .Y(\i43/i49/n239 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i265  (.A1(\i43/i49/n39 ),
    .A2(\i43/i49/n82 ),
    .B(\i43/i49/n133 ),
    .Y(\i43/i49/n280 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i266  (.A1(\i43/i49/n92 ),
    .A2(\i43/i49/n72 ),
    .B(\i43/i49/n135 ),
    .Y(\i43/i49/n279 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i267  (.A1(\i43/i49/n54 ),
    .A2(\i43/i49/n58 ),
    .B1(\i43/i49/n50 ),
    .B2(\i43/i49/n92 ),
    .Y(\i43/i49/n278 ));
 AOI22xp5_ASAP7_75t_SL \i43/i49/i268  (.A1(\i43/i49/n55 ),
    .A2(\i43/i49/n44 ),
    .B1(\i43/i49/n85 ),
    .B2(\i43/i49/n48 ),
    .Y(\i43/i49/n277 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i269  (.A1(\i43/i49/n39 ),
    .A2(\i43/i49/n37 ),
    .B(\i43/i49/n171 ),
    .Y(\i43/i49/n275 ));
 NOR3xp33_ASAP7_75t_SL \i43/i49/i27  (.A(\i43/i49/n449 ),
    .B(\i43/i49/n451 ),
    .C(\i43/i49/n434 ),
    .Y(\i43/i49/n488 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i270  (.A1(\i43/i49/n91 ),
    .A2(\i43/i49/n89 ),
    .B1(\i43/i49/n61 ),
    .B2(\i43/i49/n42 ),
    .Y(\i43/i49/n274 ));
 AOI22xp5_ASAP7_75t_SL \i43/i49/i271  (.A1(\i43/i49/n38 ),
    .A2(\i43/i49/n86 ),
    .B1(\i43/i49/n73 ),
    .B2(\i43/i49/n44 ),
    .Y(\i43/i49/n273 ));
 AOI22xp5_ASAP7_75t_SL \i43/i49/i272  (.A1(\i43/i49/n90 ),
    .A2(\i43/i49/n57 ),
    .B1(\i43/i49/n38 ),
    .B2(\i43/i49/n93 ),
    .Y(\i43/i49/n271 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i273  (.A1(\i43/i49/n80 ),
    .A2(\i43/i49/n89 ),
    .B(\i43/i49/n167 ),
    .Y(\i43/i49/n270 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i274  (.A1(\i43/i49/n89 ),
    .A2(\i43/i49/n45 ),
    .B1(\i43/i49/n40 ),
    .B2(\i43/i49/n68 ),
    .Y(\i43/i49/n1 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i275  (.A(\i43/i49/n46 ),
    .B(\i43/i49/n169 ),
    .Y(\i43/i49/n268 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i276  (.A(\i43/i49/n85 ),
    .B(\i43/i49/n168 ),
    .Y(\i43/i49/n267 ));
 NOR2xp33_ASAP7_75t_L \i43/i49/i277  (.A(\i43/i49/n50 ),
    .B(\i43/i49/n153 ),
    .Y(\i43/i49/n266 ));
 INVx1_ASAP7_75t_SL \i43/i49/i278  (.A(\i43/i49/n234 ),
    .Y(\i43/i49/n235 ));
 INVxp33_ASAP7_75t_SL \i43/i49/i279  (.A(\i43/i49/n232 ),
    .Y(\i43/i49/n233 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i28  (.A(\i43/i49/n472 ),
    .B(\i43/i49/n467 ),
    .Y(\i43/i49/n487 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i280  (.A(\i43/i49/n228 ),
    .Y(\i43/i49/n229 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i281  (.A(\i43/i49/n221 ),
    .Y(\i43/i49/n222 ));
 INVx1_ASAP7_75t_SL \i43/i49/i282  (.A(\i43/i49/n213 ),
    .Y(\i43/i49/n212 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i283  (.A1(\i43/i49/n61 ),
    .A2(\i43/i49/n39 ),
    .B1(\i43/i49/n49 ),
    .B2(\i43/i49/n45 ),
    .Y(\i43/i49/n211 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i284  (.A1(\i43/i49/n53 ),
    .A2(\i43/i49/n34 ),
    .B(\i43/i49/n44 ),
    .Y(\i43/i49/n210 ));
 OAI22xp33_ASAP7_75t_SL \i43/i49/i285  (.A1(\i43/i49/n94 ),
    .A2(\i43/i49/n91 ),
    .B1(\i43/i49/n52 ),
    .B2(\i43/i49/n61 ),
    .Y(\i43/i49/n209 ));
 OAI21xp5_ASAP7_75t_SL \i43/i49/i286  (.A1(\i43/i49/n77 ),
    .A2(\i43/i49/n65 ),
    .B(\i43/i49/n36 ),
    .Y(\i43/i49/n208 ));
 AOI21xp33_ASAP7_75t_SL \i43/i49/i287  (.A1(\i43/i49/n66 ),
    .A2(\i43/i49/n72 ),
    .B(\i43/i49/n70 ),
    .Y(\i43/i49/n207 ));
 AOI21xp33_ASAP7_75t_SL \i43/i49/i288  (.A1(\i43/i49/n45 ),
    .A2(\i43/i49/n70 ),
    .B(\i43/i49/n52 ),
    .Y(\i43/i49/n206 ));
 AOI21xp5_ASAP7_75t_SL \i43/i49/i289  (.A1(\i43/i49/n57 ),
    .A2(\i43/i49/n60 ),
    .B(\i43/i49/n129 ),
    .Y(\i43/i49/n205 ));
 AND5x1_ASAP7_75t_SL \i43/i49/i29  (.A(\i43/i49/n446 ),
    .B(\i43/i49/n421 ),
    .C(\i43/i49/n375 ),
    .D(\i43/i49/n410 ),
    .E(\i43/i49/n412 ),
    .Y(\i43/i49/n486 ));
 OAI22xp33_ASAP7_75t_SL \i43/i49/i290  (.A1(\i43/i49/n84 ),
    .A2(\i43/i49/n39 ),
    .B1(\i43/i49/n75 ),
    .B2(\i43/i49/n76 ),
    .Y(\i43/i49/n204 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i291  (.A1(\i43/i49/n75 ),
    .A2(\i43/i49/n54 ),
    .B1(\i43/i49/n40 ),
    .B2(\i43/i49/n61 ),
    .Y(\i43/i49/n203 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i292  (.A1(\i43/i49/n82 ),
    .A2(\i43/i49/n56 ),
    .B1(\i43/i49/n40 ),
    .B2(\i43/i49/n80 ),
    .Y(\i43/i49/n202 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i293  (.A1(\i43/i49/n63 ),
    .A2(\i43/i49/n49 ),
    .B1(\i43/i49/n84 ),
    .B2(\i43/i49/n46 ),
    .Y(\i43/i49/n201 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i294  (.A1(\i43/i49/n50 ),
    .A2(\i43/i49/n91 ),
    .B1(\i43/i49/n39 ),
    .B2(\i43/i49/n63 ),
    .Y(\i43/i49/n200 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i295  (.A1(\i43/i49/n49 ),
    .A2(\i43/i49/n61 ),
    .B1(\i43/i49/n68 ),
    .B2(\i43/i49/n56 ),
    .Y(\i43/i49/n199 ));
 AOI22xp5_ASAP7_75t_SL \i43/i49/i296  (.A1(\i43/i49/n81 ),
    .A2(\i43/i49/n73 ),
    .B1(\i43/i49/n43 ),
    .B2(\i43/i49/n36 ),
    .Y(\i43/i49/n238 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i297  (.A1(\i43/i49/n82 ),
    .A2(\i43/i49/n89 ),
    .B1(\i43/i49/n75 ),
    .B2(\i43/i49/n46 ),
    .Y(\i43/i49/n198 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i298  (.A1(\i43/i49/n43 ),
    .A2(\i43/i49/n88 ),
    .B1(\i43/i49/n83 ),
    .B2(\i43/i49/n33 ),
    .Y(\i43/i49/n197 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i299  (.A1(\i43/i49/n80 ),
    .A2(\i43/i49/n64 ),
    .B1(\i43/i49/n68 ),
    .B2(\i43/i49/n35 ),
    .Y(\i43/i49/n196 ));
 NOR2x1_ASAP7_75t_SL \i43/i49/i3  (.A(\i43/i49/n500 ),
    .B(\i43/i49/n505 ),
    .Y(\i43/n0 [4]));
 NOR3xp33_ASAP7_75t_SL \i43/i49/i30  (.A(\i43/i49/n462 ),
    .B(\i43/i49/n437 ),
    .C(\i43/i49/n424 ),
    .Y(\i43/i49/n485 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i300  (.A1(\i43/i49/n89 ),
    .A2(\i43/i49/n58 ),
    .B1(\i43/i49/n50 ),
    .B2(\i43/i49/n68 ),
    .Y(\i43/i49/n195 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i301  (.A1(\i43/i49/n32 ),
    .A2(\i43/i49/n89 ),
    .B1(\i43/i49/n52 ),
    .B2(\i43/i49/n58 ),
    .Y(\i43/i49/n194 ));
 AOI22xp5_ASAP7_75t_SL \i43/i49/i302  (.A1(\i43/i49/n53 ),
    .A2(\i43/i49/n79 ),
    .B1(\i43/i49/n95 ),
    .B2(\i43/i49/n44 ),
    .Y(\i43/i49/n237 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i303  (.A1(\i43/i49/n70 ),
    .A2(\i43/i49/n64 ),
    .B1(\i43/i49/n72 ),
    .B2(\i43/i49/n37 ),
    .Y(\i43/i49/n236 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i304  (.A1(\i43/i49/n32 ),
    .A2(\i43/i49/n64 ),
    .B1(\i43/i49/n42 ),
    .B2(\i43/i49/n82 ),
    .Y(\i43/i49/n234 ));
 AOI22xp5_ASAP7_75t_SL \i43/i49/i305  (.A1(\i43/i49/n93 ),
    .A2(\i43/i49/n67 ),
    .B1(\i43/i49/n43 ),
    .B2(\i43/i49/n69 ),
    .Y(\i43/i49/n232 ));
 AO22x1_ASAP7_75t_SL \i43/i49/i306  (.A1(\i43/i49/n33 ),
    .A2(\i43/i49/n34 ),
    .B1(\i43/i49/n57 ),
    .B2(\i43/i49/n81 ),
    .Y(\i43/i49/n231 ));
 AOI22xp5_ASAP7_75t_SL \i43/i49/i307  (.A1(\i43/i49/n73 ),
    .A2(\i43/i49/n79 ),
    .B1(\i43/i49/n53 ),
    .B2(\i43/i49/n69 ),
    .Y(\i43/i49/n230 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i308  (.A1(\i43/i49/n58 ),
    .A2(\i43/i49/n64 ),
    .B1(\i43/i49/n54 ),
    .B2(\i43/i49/n63 ),
    .Y(\i43/i49/n228 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i309  (.A(\i43/i49/n187 ),
    .B(\i43/i49/n188 ),
    .Y(\i43/i49/n193 ));
 NOR3xp33_ASAP7_75t_SL \i43/i49/i31  (.A(\i43/i49/n448 ),
    .B(\i43/i49/n436 ),
    .C(\i43/i49/n428 ),
    .Y(\i43/i49/n484 ));
 NAND2xp33_ASAP7_75t_SL \i43/i49/i310  (.A(\i43/i49/n186 ),
    .B(\i43/i49/n176 ),
    .Y(\i43/i49/n192 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i311  (.A1(\i43/i49/n92 ),
    .A2(\i43/i49/n40 ),
    .B1(\i43/i49/n76 ),
    .B2(\i43/i49/n70 ),
    .Y(\i43/i49/n227 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i312  (.A1(\i43/i49/n35 ),
    .A2(\i43/i49/n63 ),
    .B1(\i43/i49/n72 ),
    .B2(\i43/i49/n68 ),
    .Y(\i43/i49/n226 ));
 OAI22xp33_ASAP7_75t_SL \i43/i49/i313  (.A1(\i43/i49/n92 ),
    .A2(\i43/i49/n89 ),
    .B1(\i43/i49/n37 ),
    .B2(\i43/i49/n49 ),
    .Y(\i43/i49/n225 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i314  (.A1(\i43/i49/n92 ),
    .A2(\i43/i49/n49 ),
    .B1(\i43/i49/n42 ),
    .B2(\i43/i49/n75 ),
    .Y(\i43/i49/n224 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i315  (.A1(\i43/i49/n35 ),
    .A2(\i43/i49/n75 ),
    .B1(\i43/i49/n46 ),
    .B2(\i43/i49/n45 ),
    .Y(\i43/i49/n223 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i316  (.A1(\i43/i49/n80 ),
    .A2(\i43/i49/n39 ),
    .B1(\i43/i49/n54 ),
    .B2(\i43/i49/n68 ),
    .Y(\i43/i49/n221 ));
 AOI22xp5_ASAP7_75t_SL \i43/i49/i317  (.A1(\i43/i49/n33 ),
    .A2(\i43/i49/n57 ),
    .B1(\i43/i49/n41 ),
    .B2(\i43/i49/n36 ),
    .Y(\i43/i49/n220 ));
 OAI22xp33_ASAP7_75t_SL \i43/i49/i318  (.A1(\i43/i49/n87 ),
    .A2(\i43/i49/n89 ),
    .B1(\i43/i49/n78 ),
    .B2(\i43/i49/n42 ),
    .Y(\i43/i49/n219 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i319  (.A1(\i43/i49/n46 ),
    .A2(\i43/i49/n58 ),
    .B1(\i43/i49/n91 ),
    .B2(\i43/i49/n76 ),
    .Y(\i43/i49/n218 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i32  (.A(\i43/i49/n444 ),
    .B(\i43/i49/n474 ),
    .Y(\i43/i49/n483 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i320  (.A1(\i43/i49/n68 ),
    .A2(\i43/i49/n64 ),
    .B1(\i43/i49/n50 ),
    .B2(\i43/i49/n37 ),
    .Y(\i43/i49/n217 ));
 AOI22xp5_ASAP7_75t_SL \i43/i49/i321  (.A1(\i43/i49/n79 ),
    .A2(\i43/i49/n57 ),
    .B1(\i43/i49/n95 ),
    .B2(\i43/i49/n69 ),
    .Y(\i43/i49/n216 ));
 OAI22xp5_ASAP7_75t_SL \i43/i49/i322  (.A1(\i43/i49/n78 ),
    .A2(\i43/i49/n89 ),
    .B1(\i43/i49/n50 ),
    .B2(\i43/i49/n32 ),
    .Y(\i43/i49/n215 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i323  (.A(\i43/i49/n139 ),
    .B(\i43/i49/n138 ),
    .Y(\i43/i49/n191 ));
 AOI22xp5_ASAP7_75t_SL \i43/i49/i324  (.A1(\i43/i49/n93 ),
    .A2(\i43/i49/n34 ),
    .B1(\i43/i49/n77 ),
    .B2(\i43/i49/n62 ),
    .Y(\i43/i49/n214 ));
 OA22x2_ASAP7_75t_SL \i43/i49/i325  (.A1(\i43/i49/n61 ),
    .A2(\i43/i49/n64 ),
    .B1(\i43/i49/n58 ),
    .B2(\i43/i49/n76 ),
    .Y(\i43/i49/n213 ));
 INVx1_ASAP7_75t_SL \i43/i49/i326  (.A(\i43/i49/n189 ),
    .Y(\i43/i49/n190 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i327  (.A(\i43/i49/n182 ),
    .Y(\i43/i49/n183 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i328  (.A(\i43/i49/n176 ),
    .Y(\i43/i49/n177 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i329  (.A(\i43/i49/n174 ),
    .Y(\i43/i49/n175 ));
 NOR5xp2_ASAP7_75t_SL \i43/i49/i33  (.A(\i43/i49/n400 ),
    .B(\i43/i49/n408 ),
    .C(\i43/i49/n305 ),
    .D(\i43/i49/n397 ),
    .E(\i43/i49/n401 ),
    .Y(\i43/i49/n482 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i330  (.A(\i43/i49/n168 ),
    .Y(\i43/i49/n169 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i331  (.A(\i43/i49/n165 ),
    .Y(\i43/i49/n166 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i332  (.A(\i43/i49/n160 ),
    .Y(\i43/i49/n161 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i333  (.A(\i43/i49/n155 ),
    .Y(\i43/i49/n156 ));
 INVx1_ASAP7_75t_SL \i43/i49/i334  (.A(\i43/i49/n153 ),
    .Y(\i43/i49/n154 ));
 INVx1_ASAP7_75t_SL \i43/i49/i335  (.A(\i43/i49/n151 ),
    .Y(\i43/i49/n152 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i336  (.A(\i43/i49/n149 ),
    .Y(\i43/i49/n150 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i337  (.A(\i43/i49/n147 ),
    .Y(\i43/i49/n148 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i338  (.A(\i43/i49/n85 ),
    .B(\i43/i49/n51 ),
    .Y(\i43/i49/n146 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i339  (.A(\i43/i49/n77 ),
    .B(\i43/i49/n81 ),
    .Y(\i43/i49/n189 ));
 NAND5xp2_ASAP7_75t_SL \i43/i49/i34  (.A(\i43/i49/n390 ),
    .B(\i43/i49/n417 ),
    .C(\i43/i49/n352 ),
    .D(\i43/i49/n318 ),
    .E(\i43/i49/n349 ),
    .Y(\i43/i49/n481 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i340  (.A(\i43/i49/n41 ),
    .B(\i43/i49/n90 ),
    .Y(\i43/i49/n145 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i341  (.A(\i43/i49/n90 ),
    .B(\i43/i49/n48 ),
    .Y(\i43/i49/n144 ));
 NAND2xp33_ASAP7_75t_SL \i43/i49/i342  (.A(\i43/i49/n46 ),
    .B(\i43/i49/n64 ),
    .Y(\i43/i49/n143 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i343  (.A(\i43/i49/n36 ),
    .B(\i43/i49/n65 ),
    .Y(\i43/i49/n188 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i344  (.A(\i43/i49/n95 ),
    .B(\i43/i49/n93 ),
    .Y(\i43/i49/n187 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i345  (.A(\i43/i49/n67 ),
    .B(\i43/i49/n59 ),
    .Y(\i43/i49/n186 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i346  (.A(\i43/i49/n85 ),
    .B(\i43/i49/n71 ),
    .Y(\i43/i49/n142 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i347  (.A(\i43/i49/n58 ),
    .B(\i43/i49/n50 ),
    .Y(\i43/i49/n141 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i348  (.A(\i43/i49/n55 ),
    .B(\i43/i49/n83 ),
    .Y(\i43/i49/n185 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i349  (.A(\i43/i49/n69 ),
    .B(\i43/i49/n41 ),
    .Y(\i43/i49/n140 ));
 NOR2xp33_ASAP7_75t_L \i43/i49/i35  (.A(\i43/i49/n455 ),
    .B(\i43/i49/n478 ),
    .Y(\i43/i49/n480 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i350  (.A(\i43/i49/n77 ),
    .B(\i43/i49/n93 ),
    .Y(\i43/i49/n184 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i351  (.A(\i43/i49/n75 ),
    .B(\i43/i49/n40 ),
    .Y(\i43/i49/n182 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i352  (.A(\i43/i49/n69 ),
    .B(\i43/i49/n67 ),
    .Y(\i43/i49/n181 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i353  (.A(\i43/i49/n79 ),
    .B(\i43/i49/n51 ),
    .Y(\i43/i49/n180 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i354  (.A(\i43/i49/n93 ),
    .B(\i43/i49/n65 ),
    .Y(\i43/i49/n179 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i355  (.A(\i43/i49/n79 ),
    .B(\i43/i49/n95 ),
    .Y(\i43/i49/n178 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i356  (.A(\i43/i49/n74 ),
    .B(\i43/i49/n65 ),
    .Y(\i43/i49/n176 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i357  (.A(\i43/i49/n86 ),
    .B(\i43/i49/n77 ),
    .Y(\i43/i49/n174 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i358  (.A(\i43/i49/n85 ),
    .B(\i43/i49/n69 ),
    .Y(\i43/i49/n173 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i359  (.A(\i43/i49/n95 ),
    .B(\i43/i49/n36 ),
    .Y(\i43/i49/n172 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i36  (.A(\i43/i49/n416 ),
    .B(\i43/i49/n477 ),
    .Y(\i43/i49/n479 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i360  (.A(\i43/i49/n44 ),
    .B(\i43/i49/n65 ),
    .Y(\i43/i49/n171 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i361  (.A(\i43/i49/n91 ),
    .B(\i43/i49/n46 ),
    .Y(\i43/i49/n170 ));
 NAND2xp5_ASAP7_75t_L \i43/i49/i362  (.A(\i43/i49/n35 ),
    .B(\i43/i49/n94 ),
    .Y(\i43/i49/n168 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i363  (.A(\i43/i49/n95 ),
    .B(\i43/i49/n33 ),
    .Y(\i43/i49/n167 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i364  (.A(\i43/i49/n95 ),
    .B(\i43/i49/n43 ),
    .Y(\i43/i49/n165 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i365  (.A(\i43/i49/n57 ),
    .B(\i43/i49/n59 ),
    .Y(\i43/i49/n164 ));
 NAND2xp33_ASAP7_75t_SL \i43/i49/i366  (.A(\i43/i49/n61 ),
    .B(\i43/i49/n87 ),
    .Y(\i43/i49/n163 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i367  (.A(\i43/i49/n59 ),
    .B(\i43/i49/n41 ),
    .Y(\i43/i49/n162 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i368  (.A(\i43/i49/n73 ),
    .B(\i43/i49/n59 ),
    .Y(\i43/i49/n160 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i369  (.A(\i43/i49/n77 ),
    .B(\i43/i49/n83 ),
    .Y(\i43/i49/n159 ));
 INVx1_ASAP7_75t_SL \i43/i49/i37  (.A(\i43/i49/n509 ),
    .Y(\i43/i49/n475 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i370  (.A(\i43/i49/n85 ),
    .B(\i43/i49/n57 ),
    .Y(\i43/i49/n158 ));
 NOR2xp33_ASAP7_75t_L \i43/i49/i371  (.A(\i43/i49/n60 ),
    .B(\i43/i49/n69 ),
    .Y(\i43/i49/n157 ));
 NAND2xp5_ASAP7_75t_L \i43/i49/i372  (.A(\i43/i49/n37 ),
    .B(\i43/i49/n68 ),
    .Y(\i43/i49/n155 ));
 NOR2x1_ASAP7_75t_SL \i43/i49/i373  (.A(\i43/i49/n62 ),
    .B(\i43/i49/n71 ),
    .Y(\i43/i49/n153 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i374  (.A(\i43/i49/n88 ),
    .B(\i43/i49/n36 ),
    .Y(\i43/i49/n151 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i375  (.A(\i43/i49/n86 ),
    .B(\i43/i49/n62 ),
    .Y(\i43/i49/n149 ));
 NAND2x1_ASAP7_75t_SL \i43/i49/i376  (.A(\i43/i49/n84 ),
    .B(\i43/i49/n63 ),
    .Y(\i43/i49/n0 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i377  (.A(\i43/i49/n32 ),
    .B(\i43/i49/n91 ),
    .Y(\i43/i49/n147 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i378  (.A(\i43/i49/n130 ),
    .Y(\i43/i49/n131 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i379  (.A(\i43/i49/n121 ),
    .Y(\i43/i49/n122 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i38  (.A(\i43/i49/n453 ),
    .B(\i43/i49/n422 ),
    .Y(\i43/i49/n473 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i380  (.A(\i43/i49/n118 ),
    .Y(\i43/i49/n119 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i381  (.A(\i43/i49/n55 ),
    .B(\i43/i49/n36 ),
    .Y(\i43/i49/n116 ));
 NAND2xp33_ASAP7_75t_SL \i43/i49/i382  (.A(\i43/i49/n70 ),
    .B(\i43/i49/n61 ),
    .Y(\i43/i49/n115 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i383  (.A(\i43/i49/n48 ),
    .B(\i43/i49/n57 ),
    .Y(\i43/i49/n114 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i384  (.A(\i43/i49/n51 ),
    .B(\i43/i49/n83 ),
    .Y(\i43/i49/n113 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i385  (.A(\i43/i49/n57 ),
    .B(\i43/i49/n36 ),
    .Y(\i43/i49/n139 ));
 NAND2xp33_ASAP7_75t_SL \i43/i49/i386  (.A(\i43/i49/n82 ),
    .B(\i43/i49/n45 ),
    .Y(\i43/i49/n112 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i387  (.A(\i43/i49/n71 ),
    .B(\i43/i49/n55 ),
    .Y(\i43/i49/n111 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i388  (.A(\i43/i49/n33 ),
    .B(\i43/i49/n38 ),
    .Y(\i43/i49/n110 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i389  (.A(\i43/i49/n75 ),
    .B(\i43/i49/n82 ),
    .Y(\i43/i49/n109 ));
 NAND2xp33_ASAP7_75t_L \i43/i49/i39  (.A(\i43/i49/n453 ),
    .B(\i43/i49/n433 ),
    .Y(\i43/i49/n472 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i390  (.A(\i43/i49/n93 ),
    .B(\i43/i49/n53 ),
    .Y(\i43/i49/n108 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i391  (.A(\i43/i49/n44 ),
    .B(\i43/i49/n43 ),
    .Y(\i43/i49/n138 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i392  (.A(\i43/i49/n60 ),
    .B(\i43/i49/n34 ),
    .Y(\i43/i49/n107 ));
 NAND2xp33_ASAP7_75t_SL \i43/i49/i393  (.A(\i43/i49/n39 ),
    .B(\i43/i49/n66 ),
    .Y(\i43/i49/n106 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i394  (.A(\i43/i49/n47 ),
    .B(\i43/i49/n33 ),
    .Y(\i43/i49/n105 ));
 NAND2xp5_ASAP7_75t_L \i43/i49/i395  (.A(\i43/i49/n42 ),
    .B(\i43/i49/n66 ),
    .Y(\i43/i49/n104 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i396  (.A(\i43/i49/n38 ),
    .B(\i43/i49/n73 ),
    .Y(\i43/i49/n103 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i397  (.A(\i43/i49/n73 ),
    .B(\i43/i49/n60 ),
    .Y(\i43/i49/n137 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i398  (.A(\i43/i49/n41 ),
    .B(\i43/i49/n73 ),
    .Y(\i43/i49/n136 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i399  (.A(\i43/i49/n74 ),
    .B(\i43/i49/n48 ),
    .Y(\i43/i49/n135 ));
 AND5x1_ASAP7_75t_SL \i43/i49/i4  (.A(\i43/i49/n501 ),
    .B(\i43/i49/n498 ),
    .C(\i43/i49/n477 ),
    .D(\i43/i49/n499 ),
    .E(\i43/i49/n468 ),
    .Y(\i43/n0 [3]));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i40  (.A(\i43/i49/n450 ),
    .B(\i43/i49/n432 ),
    .Y(\i43/i49/n471 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i400  (.A(\i43/i49/n72 ),
    .B(\i43/i49/n45 ),
    .Y(\i43/i49/n102 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i401  (.A(\i43/i49/n67 ),
    .B(\i43/i49/n36 ),
    .Y(\i43/i49/n134 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i402  (.A(\i43/i49/n47 ),
    .B(\i43/i49/n93 ),
    .Y(\i43/i49/n133 ));
 NOR2xp33_ASAP7_75t_L \i43/i49/i403  (.A(\i43/i49/n35 ),
    .B(\i43/i49/n37 ),
    .Y(\i43/i49/n132 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i404  (.A(\i43/i49/n42 ),
    .B(\i43/i49/n75 ),
    .Y(\i43/i49/n101 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i405  (.A(\i43/i49/n71 ),
    .B(\i43/i49/n34 ),
    .Y(\i43/i49/n100 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i406  (.A(\i43/i49/n51 ),
    .B(\i43/i49/n44 ),
    .Y(\i43/i49/n130 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i407  (.A(\i43/i49/n92 ),
    .B(\i43/i49/n42 ),
    .Y(\i43/i49/n129 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i408  (.A(\i43/i49/n47 ),
    .B(\i43/i49/n81 ),
    .Y(\i43/i49/n128 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i409  (.A(\i43/i49/n47 ),
    .B(\i43/i49/n60 ),
    .Y(\i43/i49/n127 ));
 NAND4xp25_ASAP7_75t_SL \i43/i49/i41  (.A(\i43/i49/n415 ),
    .B(\i43/i49/n308 ),
    .C(\i43/i49/n311 ),
    .D(\i43/i49/n343 ),
    .Y(\i43/i49/n470 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i410  (.A(\i43/i49/n74 ),
    .B(\i43/i49/n51 ),
    .Y(\i43/i49/n126 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i411  (.A(\i43/i49/n38 ),
    .B(\i43/i49/n93 ),
    .Y(\i43/i49/n99 ));
 NOR2xp33_ASAP7_75t_L \i43/i49/i412  (.A(\i43/i49/n50 ),
    .B(\i43/i49/n80 ),
    .Y(\i43/i49/n125 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i413  (.A(\i43/i49/n50 ),
    .B(\i43/i49/n92 ),
    .Y(\i43/i49/n98 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i414  (.A(\i43/i49/n61 ),
    .B(\i43/i49/n42 ),
    .Y(\i43/i49/n97 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i415  (.A(\i43/i49/n93 ),
    .B(\i43/i49/n57 ),
    .Y(\i43/i49/n124 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i416  (.A(\i43/i49/n55 ),
    .B(\i43/i49/n44 ),
    .Y(\i43/i49/n96 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i417  (.A(\i43/i49/n79 ),
    .B(\i43/i49/n38 ),
    .Y(\i43/i49/n123 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i418  (.A(\i43/i49/n49 ),
    .B(\i43/i49/n32 ),
    .Y(\i43/i49/n121 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i419  (.A(\i43/i49/n33 ),
    .B(\i43/i49/n53 ),
    .Y(\i43/i49/n120 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i42  (.A(\i43/i49/n433 ),
    .B(\i43/i49/n442 ),
    .Y(\i43/i49/n478 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i420  (.A(\i43/i49/n83 ),
    .B(\i43/i49/n53 ),
    .Y(\i43/i49/n118 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i421  (.A(\i43/i49/n60 ),
    .B(\i43/i49/n51 ),
    .Y(\i43/i49/n117 ));
 INVx1_ASAP7_75t_SL \i43/i49/i422  (.A(\i43/i49/n95 ),
    .Y(\i43/i49/n94 ));
 INVx2_ASAP7_75t_SL \i43/i49/i423  (.A(\i43/i49/n93 ),
    .Y(\i43/i49/n92 ));
 INVx1_ASAP7_75t_SL \i43/i49/i424  (.A(\i43/i49/n91 ),
    .Y(\i43/i49/n90 ));
 INVx2_ASAP7_75t_SL \i43/i49/i425  (.A(\i43/i49/n89 ),
    .Y(\i43/i49/n88 ));
 INVx2_ASAP7_75t_SL \i43/i49/i426  (.A(\i43/i49/n87 ),
    .Y(\i43/i49/n86 ));
 INVx2_ASAP7_75t_SL \i43/i49/i427  (.A(\i43/i49/n85 ),
    .Y(\i43/i49/n84 ));
 INVx3_ASAP7_75t_SL \i43/i49/i428  (.A(\i43/i49/n83 ),
    .Y(\i43/i49/n82 ));
 INVx2_ASAP7_75t_SL \i43/i49/i429  (.A(\i43/i49/n81 ),
    .Y(\i43/i49/n80 ));
 AND4x1_ASAP7_75t_SL \i43/i49/i43  (.A(\i43/i49/n435 ),
    .B(\i43/i49/n415 ),
    .C(\i43/i49/n353 ),
    .D(\i43/i49/n193 ),
    .Y(\i43/i49/n469 ));
 INVx2_ASAP7_75t_SL \i43/i49/i430  (.A(\i43/i49/n79 ),
    .Y(\i43/i49/n78 ));
 INVx2_ASAP7_75t_SL \i43/i49/i431  (.A(\i43/i49/n77 ),
    .Y(\i43/i49/n76 ));
 INVx2_ASAP7_75t_SL \i43/i49/i432  (.A(\i43/i49/n75 ),
    .Y(\i43/i49/n74 ));
 INVx2_ASAP7_75t_SL \i43/i49/i433  (.A(\i43/i49/n73 ),
    .Y(\i43/i49/n72 ));
 INVx2_ASAP7_75t_SL \i43/i49/i434  (.A(\i43/i49/n71 ),
    .Y(\i43/i49/n70 ));
 INVx2_ASAP7_75t_SL \i43/i49/i435  (.A(\i43/i49/n69 ),
    .Y(\i43/i49/n68 ));
 INVx2_ASAP7_75t_SL \i43/i49/i436  (.A(\i43/i49/n67 ),
    .Y(\i43/i49/n66 ));
 INVx2_ASAP7_75t_SL \i43/i49/i437  (.A(\i43/i49/n65 ),
    .Y(\i43/i49/n64 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i438  (.A(\i43/i49/n25 ),
    .B(\i43/i49/n15 ),
    .Y(\i43/i49/n95 ));
 AND2x4_ASAP7_75t_SL \i43/i49/i439  (.A(\i43/i49/n5 ),
    .B(\i43/i49/n6 ),
    .Y(\i43/i49/n93 ));
 AND4x1_ASAP7_75t_SL \i43/i49/i44  (.A(\i43/i49/n380 ),
    .B(\i43/i49/n317 ),
    .C(\i43/i49/n368 ),
    .D(\i43/i49/n189 ),
    .Y(\i43/i49/n477 ));
 OR2x2_ASAP7_75t_SL \i43/i49/i440  (.A(\i43/i49/n27 ),
    .B(\i43/i49/n11 ),
    .Y(\i43/i49/n91 ));
 OR2x2_ASAP7_75t_SL \i43/i49/i441  (.A(\i43/i49/n28 ),
    .B(\i43/i49/n9 ),
    .Y(\i43/i49/n89 ));
 OR2x6_ASAP7_75t_SL \i43/i49/i442  (.A(\i43/i49/n7 ),
    .B(\i43/i49/n11 ),
    .Y(\i43/i49/n87 ));
 AND2x4_ASAP7_75t_SL \i43/i49/i443  (.A(\i43/i49/n4 ),
    .B(\i43/i49/n19 ),
    .Y(\i43/i49/n85 ));
 AND2x4_ASAP7_75t_SL \i43/i49/i444  (.A(\i43/i49/n10 ),
    .B(\i43/i49/n22 ),
    .Y(\i43/i49/n83 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i445  (.A(\i43/i49/n6 ),
    .B(\i43/i49/n19 ),
    .Y(\i43/i49/n81 ));
 AND2x4_ASAP7_75t_SL \i43/i49/i446  (.A(\i43/i49/n5 ),
    .B(\i43/i49/n26 ),
    .Y(\i43/i49/n79 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i447  (.A(\i43/i49/n16 ),
    .B(\i43/i49/n15 ),
    .Y(\i43/i49/n77 ));
 OR2x2_ASAP7_75t_SL \i43/i49/i448  (.A(\i43/i49/n3 ),
    .B(\i43/i49/n31 ),
    .Y(\i43/i49/n75 ));
 AND2x4_ASAP7_75t_SL \i43/i49/i449  (.A(\i43/i49/n25 ),
    .B(\i43/i49/n12 ),
    .Y(\i43/i49/n73 ));
 NOR2x1_ASAP7_75t_SL \i43/i49/i45  (.A(\i43/i49/n306 ),
    .B(\i43/i49/n451 ),
    .Y(\i43/i49/n476 ));
 AND2x4_ASAP7_75t_SL \i43/i49/i450  (.A(\i43/i49/n4 ),
    .B(\i43/i49/n10 ),
    .Y(\i43/i49/n71 ));
 AND2x4_ASAP7_75t_SL \i43/i49/i451  (.A(\i43/i49/n5 ),
    .B(\i43/i49/n4 ),
    .Y(\i43/i49/n69 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i452  (.A(\i43/i49/n16 ),
    .B(\i43/i49/n29 ),
    .Y(\i43/i49/n67 ));
 AND2x4_ASAP7_75t_SL \i43/i49/i453  (.A(\i43/i49/n8 ),
    .B(\i43/i49/n12 ),
    .Y(\i43/i49/n65 ));
 INVx2_ASAP7_75t_SL \i43/i49/i454  (.A(\i43/i49/n63 ),
    .Y(\i43/i49/n62 ));
 INVx3_ASAP7_75t_SL \i43/i49/i455  (.A(\i43/i49/n61 ),
    .Y(\i43/i49/n60 ));
 INVx2_ASAP7_75t_SL \i43/i49/i456  (.A(\i43/i49/n59 ),
    .Y(\i43/i49/n58 ));
 INVx1_ASAP7_75t_SL \i43/i49/i457  (.A(\i43/i49/n57 ),
    .Y(\i43/i49/n56 ));
 INVx2_ASAP7_75t_SL \i43/i49/i458  (.A(\i43/i49/n55 ),
    .Y(\i43/i49/n54 ));
 INVx4_ASAP7_75t_SL \i43/i49/i459  (.A(\i43/i49/n53 ),
    .Y(\i43/i49/n52 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i46  (.A(\i43/i49/n392 ),
    .B(\i43/i49/n426 ),
    .Y(\i43/i49/n474 ));
 INVx2_ASAP7_75t_SL \i43/i49/i460  (.A(\i43/i49/n51 ),
    .Y(\i43/i49/n50 ));
 INVx2_ASAP7_75t_SL \i43/i49/i461  (.A(\i43/i49/n49 ),
    .Y(\i43/i49/n48 ));
 INVx2_ASAP7_75t_SL \i43/i49/i462  (.A(\i43/i49/n47 ),
    .Y(\i43/i49/n46 ));
 INVx4_ASAP7_75t_SL \i43/i49/i463  (.A(\i43/i49/n45 ),
    .Y(\i43/i49/n44 ));
 INVx4_ASAP7_75t_SL \i43/i49/i464  (.A(\i43/i49/n43 ),
    .Y(\i43/i49/n42 ));
 INVx2_ASAP7_75t_SL \i43/i49/i465  (.A(\i43/i49/n41 ),
    .Y(\i43/i49/n40 ));
 INVx2_ASAP7_75t_SL \i43/i49/i466  (.A(\i43/i49/n39 ),
    .Y(\i43/i49/n38 ));
 INVx2_ASAP7_75t_SL \i43/i49/i467  (.A(\i43/i49/n37 ),
    .Y(\i43/i49/n36 ));
 INVx3_ASAP7_75t_SL \i43/i49/i468  (.A(\i43/i49/n35 ),
    .Y(\i43/i49/n34 ));
 INVx2_ASAP7_75t_SL \i43/i49/i469  (.A(\i43/i49/n33 ),
    .Y(\i43/i49/n32 ));
 INVx1_ASAP7_75t_SL \i43/i49/i47  (.A(\i43/i49/n466 ),
    .Y(\i43/i49/n467 ));
 NAND2x1p5_ASAP7_75t_SL \i43/i49/i470  (.A(\i43/i49/n22 ),
    .B(\i43/i49/n5 ),
    .Y(\i43/i49/n63 ));
 OR2x2_ASAP7_75t_SL \i43/i49/i471  (.A(\i43/i49/n27 ),
    .B(\i43/i49/n20 ),
    .Y(\i43/i49/n61 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i472  (.A(\i43/i49/n6 ),
    .B(\i43/i49/n30 ),
    .Y(\i43/i49/n59 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i473  (.A(\i43/i49/n25 ),
    .B(\i43/i49/n18 ),
    .Y(\i43/i49/n57 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i474  (.A(\i43/i49/n8 ),
    .B(\i43/i49/n18 ),
    .Y(\i43/i49/n55 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i475  (.A(\i43/i49/n16 ),
    .B(\i43/i49/n12 ),
    .Y(\i43/i49/n53 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i476  (.A(\i43/i49/n25 ),
    .B(\i43/i49/n29 ),
    .Y(\i43/i49/n51 ));
 OR2x2_ASAP7_75t_SL \i43/i49/i477  (.A(\i43/i49/n17 ),
    .B(\i43/i49/n24 ),
    .Y(\i43/i49/n49 ));
 AND2x4_ASAP7_75t_SL \i43/i49/i478  (.A(\i43/i49/n23 ),
    .B(\i43/i49/n15 ),
    .Y(\i43/i49/n47 ));
 OR2x2_ASAP7_75t_SL \i43/i49/i479  (.A(\i43/i49/n27 ),
    .B(\i43/i49/n31 ),
    .Y(\i43/i49/n45 ));
 NAND2xp5_ASAP7_75t_L \i43/i49/i48  (.A(\i43/i49/n435 ),
    .B(\i43/i49/n419 ),
    .Y(\i43/i49/n464 ));
 AND2x4_ASAP7_75t_SL \i43/i49/i480  (.A(\i43/i49/n23 ),
    .B(\i43/i49/n29 ),
    .Y(\i43/i49/n43 ));
 AND2x4_ASAP7_75t_SL \i43/i49/i481  (.A(\i43/i49/n16 ),
    .B(\i43/i49/n18 ),
    .Y(\i43/i49/n41 ));
 OR2x2_ASAP7_75t_SL \i43/i49/i482  (.A(\i43/i49/n14 ),
    .B(\i43/i49/n9 ),
    .Y(\i43/i49/n39 ));
 OR2x6_ASAP7_75t_SL \i43/i49/i483  (.A(\i43/i49/n20 ),
    .B(\i43/i49/n21 ),
    .Y(\i43/i49/n37 ));
 OR2x6_ASAP7_75t_SL \i43/i49/i484  (.A(\i43/i49/n24 ),
    .B(\i43/i49/n13 ),
    .Y(\i43/i49/n35 ));
 AND2x4_ASAP7_75t_SL \i43/i49/i485  (.A(\i43/i49/n30 ),
    .B(\i43/i49/n22 ),
    .Y(\i43/i49/n33 ));
 INVx2_ASAP7_75t_SL \i43/i49/i486  (.A(\i43/i49/n31 ),
    .Y(\i43/i49/n30 ));
 INVx2_ASAP7_75t_SL \i43/i49/i487  (.A(\i43/i49/n28 ),
    .Y(\i43/i49/n29 ));
 INVxp67_ASAP7_75t_SL \i43/i49/i488  (.A(\i43/i49/n27 ),
    .Y(\i43/i49/n26 ));
 INVx2_ASAP7_75t_SL \i43/i49/i489  (.A(\i43/i49/n24 ),
    .Y(\i43/i49/n23 ));
 AND3x1_ASAP7_75t_SL \i43/i49/i49  (.A(\i43/i49/n420 ),
    .B(\i43/i49/n405 ),
    .C(\i43/i49/n391 ),
    .Y(\i43/i49/n463 ));
 INVx3_ASAP7_75t_SL \i43/i49/i490  (.A(\i43/i49/n21 ),
    .Y(\i43/i49/n22 ));
 INVx2_ASAP7_75t_SL \i43/i49/i491  (.A(\i43/i49/n20 ),
    .Y(\i43/i49/n19 ));
 INVx1_ASAP7_75t_SL \i43/i49/i492  (.A(\i43/i49/n17 ),
    .Y(\i43/i49/n18 ));
 OR2x2_ASAP7_75t_SL \i43/i49/i493  (.A(n58),
    .B(n34[29]),
    .Y(\i43/i49/n31 ));
 OR2x2_ASAP7_75t_SL \i43/i49/i494  (.A(n59),
    .B(n34[24]),
    .Y(\i43/i49/n28 ));
 OR2x2_ASAP7_75t_SL \i43/i49/i495  (.A(n56),
    .B(n34[31]),
    .Y(\i43/i49/n27 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i496  (.A(n34[25]),
    .B(n60),
    .Y(\i43/i49/n25 ));
 NAND2x1_ASAP7_75t_SL \i43/i49/i497  (.A(n34[26]),
    .B(n61),
    .Y(\i43/i49/n24 ));
 OR2x2_ASAP7_75t_SL \i43/i49/i498  (.A(\i43/i49/n2 ),
    .B(n34[30]),
    .Y(\i43/i49/n21 ));
 OR2x2_ASAP7_75t_SL \i43/i49/i499  (.A(n57),
    .B(n34[28]),
    .Y(\i43/i49/n20 ));
 NAND5xp2_ASAP7_75t_SL \i43/i49/i5  (.A(\i43/i49/n466 ),
    .B(\i43/i49/n476 ),
    .C(\i43/i49/n471 ),
    .D(\i43/i49/n460 ),
    .E(\i43/i49/n454 ),
    .Y(\i43/i49/n507 ));
 NAND4xp25_ASAP7_75t_SL \i43/i49/i50  (.A(\i43/i49/n418 ),
    .B(\i43/i49/n384 ),
    .C(\i43/i49/n312 ),
    .D(\i43/i49/n309 ),
    .Y(\i43/i49/n462 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i500  (.A(n34[24]),
    .B(n59),
    .Y(\i43/i49/n17 ));
 INVx1_ASAP7_75t_SL \i43/i49/i501  (.A(\i43/i49/n14 ),
    .Y(\i43/i49/n15 ));
 INVx2_ASAP7_75t_SL \i43/i49/i502  (.A(\i43/i49/n12 ),
    .Y(\i43/i49/n13 ));
 INVx1_ASAP7_75t_SL \i43/i49/i503  (.A(\i43/i49/n11 ),
    .Y(\i43/i49/n10 ));
 INVx1_ASAP7_75t_SL \i43/i49/i504  (.A(\i43/i49/n9 ),
    .Y(\i43/i49/n8 ));
 INVx1_ASAP7_75t_SL \i43/i49/i505  (.A(\i43/i49/n6 ),
    .Y(\i43/i49/n7 ));
 INVx2_ASAP7_75t_SL \i43/i49/i506  (.A(\i43/i49/n3 ),
    .Y(\i43/i49/n4 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i507  (.A(n34[26]),
    .B(n34[25]),
    .Y(\i43/i49/n16 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i508  (.A(n34[27]),
    .B(n34[24]),
    .Y(\i43/i49/n14 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i509  (.A(n59),
    .B(n62),
    .Y(\i43/i49/n12 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i51  (.A(\i43/i49/n247 ),
    .B(\i43/i49/n510 ),
    .Y(\i43/i49/n461 ));
 OR2x2_ASAP7_75t_SL \i43/i49/i510  (.A(n34[29]),
    .B(n34[28]),
    .Y(\i43/i49/n11 ));
 OR2x2_ASAP7_75t_SL \i43/i49/i511  (.A(n34[26]),
    .B(n34[25]),
    .Y(\i43/i49/n9 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i512  (.A(\i43/i49/n2 ),
    .B(n56),
    .Y(\i43/i49/n6 ));
 AND2x2_ASAP7_75t_SL \i43/i49/i513  (.A(n34[29]),
    .B(n34[28]),
    .Y(\i43/i49/n5 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i514  (.A(n34[31]),
    .B(n34[30]),
    .Y(\i43/i49/n3 ));
 INVx1_ASAP7_75t_SL \i43/i49/i515  (.A(n34[31]),
    .Y(\i43/i49/n2 ));
 OR4x1_ASAP7_75t_SL \i43/i49/i516  (.A(\i43/i49/n450 ),
    .B(\i43/i49/n278 ),
    .C(\i43/i49/n248 ),
    .D(\i43/i49/n226 ),
    .Y(\i43/i49/n508 ));
 NAND5xp2_ASAP7_75t_SL \i43/i49/i517  (.A(\i43/i49/n452 ),
    .B(\i43/i49/n288 ),
    .C(\i43/i49/n277 ),
    .D(\i43/i49/n220 ),
    .E(\i43/i49/n414 ),
    .Y(\i43/i49/n509 ));
 AND3x1_ASAP7_75t_SL \i43/i49/i518  (.A(\i43/i49/n326 ),
    .B(\i43/i49/n267 ),
    .C(\i43/i49/n329 ),
    .Y(\i43/i49/n510 ));
 OR3x1_ASAP7_75t_SL \i43/i49/i519  (.A(\i43/i49/n223 ),
    .B(\i43/i49/n132 ),
    .C(\i43/i49/n199 ),
    .Y(\i43/i49/n511 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i52  (.A(\i43/i49/n411 ),
    .B(\i43/i49/n441 ),
    .Y(\i43/i49/n460 ));
 NAND3xp33_ASAP7_75t_SL \i43/i49/i520  (.A(\i43/i49/n230 ),
    .B(\i43/i49/n117 ),
    .C(\i43/i49/n107 ),
    .Y(\i43/i49/n512 ));
 NAND3xp33_ASAP7_75t_SL \i43/i49/i521  (.A(\i43/i49/n513 ),
    .B(\i43/i49/n302 ),
    .C(\i43/i49/n151 ),
    .Y(\i43/i49/n514 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i522  (.A(\i43/i49/n228 ),
    .B(\i43/i49/n124 ),
    .Y(\i43/i49/n513 ));
 NOR3xp33_ASAP7_75t_SL \i43/i49/i53  (.A(\i43/i49/n383 ),
    .B(\i43/i49/n398 ),
    .C(\i43/i49/n304 ),
    .Y(\i43/i49/n459 ));
 AOI211xp5_ASAP7_75t_SL \i43/i49/i54  (.A1(\i43/i49/n378 ),
    .A2(\i43/i49/n4 ),
    .B(\i43/i49/n394 ),
    .C(\i43/i49/n396 ),
    .Y(\i43/i49/n458 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i55  (.A(\i43/i49/n425 ),
    .B(\i43/i49/n431 ),
    .Y(\i43/i49/n457 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i56  (.A(\i43/i49/n393 ),
    .B(\i43/i49/n434 ),
    .Y(\i43/i49/n456 ));
 NOR2xp33_ASAP7_75t_L \i43/i49/i57  (.A(\i43/i49/n411 ),
    .B(\i43/i49/n430 ),
    .Y(\i43/i49/n468 ));
 OA211x2_ASAP7_75t_SL \i43/i49/i58  (.A1(\i43/i49/n91 ),
    .A2(\i43/i49/n66 ),
    .B(\i43/i49/n391 ),
    .C(\i43/i49/n370 ),
    .Y(\i43/i49/n466 ));
 NAND3xp33_ASAP7_75t_SL \i43/i49/i59  (.A(\i43/i49/n353 ),
    .B(\i43/i49/n379 ),
    .C(\i43/i49/n320 ),
    .Y(\i43/i49/n465 ));
 AND4x1_ASAP7_75t_SL \i43/i49/i6  (.A(\i43/i49/n495 ),
    .B(\i43/i49/n499 ),
    .C(\i43/i49/n484 ),
    .D(\i43/i49/n457 ),
    .Y(\i43/n0 [0]));
 INVxp67_ASAP7_75t_SL \i43/i49/i60  (.A(\i43/i49/n510 ),
    .Y(\i43/i49/n449 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i61  (.A(\i43/i49/n407 ),
    .B(\i43/i49/n392 ),
    .Y(\i43/i49/n448 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i62  (.A(\i43/i49/n300 ),
    .B(\i43/i49/n407 ),
    .Y(\i43/i49/n447 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i63  (.A(\i43/i49/n390 ),
    .B(\i43/i49/n387 ),
    .Y(\i43/i49/n455 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i64  (.A(\i43/i49/n511 ),
    .B(\i43/i49/n382 ),
    .Y(\i43/i49/n446 ));
 NAND2xp5_ASAP7_75t_L \i43/i49/i65  (.A(\i43/i49/n388 ),
    .B(\i43/i49/n310 ),
    .Y(\i43/i49/n445 ));
 NOR3xp33_ASAP7_75t_SL \i43/i49/i66  (.A(\i43/i49/n413 ),
    .B(\i43/i49/n342 ),
    .C(\i43/i49/n344 ),
    .Y(\i43/i49/n454 ));
 NAND3xp33_ASAP7_75t_SL \i43/i49/i67  (.A(\i43/i49/n389 ),
    .B(\i43/i49/n341 ),
    .C(\i43/i49/n216 ),
    .Y(\i43/i49/n444 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i68  (.A(\i43/i49/n299 ),
    .B(\i43/i49/n374 ),
    .Y(\i43/i49/n443 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i69  (.A(\i43/i49/n386 ),
    .B(\i43/i49/n512 ),
    .Y(\i43/i49/n442 ));
 AND4x1_ASAP7_75t_L \i43/i49/i7  (.A(\i43/i49/n485 ),
    .B(\i43/i49/n490 ),
    .C(\i43/i49/n498 ),
    .D(\i43/i49/n487 ),
    .Y(\i43/n0 [7]));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i70  (.A(\i43/i49/n353 ),
    .B(\i43/i49/n399 ),
    .Y(\i43/i49/n441 ));
 OA211x2_ASAP7_75t_SL \i43/i49/i71  (.A1(\i43/i49/n66 ),
    .A2(\i43/i49/n87 ),
    .B(\i43/i49/n365 ),
    .C(\i43/i49/n368 ),
    .Y(\i43/i49/n440 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i72  (.A(\i43/i49/n514 ),
    .B(\i43/i49/n403 ),
    .Y(\i43/i49/n439 ));
 AND3x1_ASAP7_75t_SL \i43/i49/i73  (.A(\i43/i49/n352 ),
    .B(\i43/i49/n363 ),
    .C(\i43/i49/n348 ),
    .Y(\i43/i49/n438 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i74  (.A(\i43/i49/n377 ),
    .B(\i43/i49/n364 ),
    .Y(\i43/i49/n453 ));
 NOR3xp33_ASAP7_75t_SL \i43/i49/i75  (.A(\i43/i49/n327 ),
    .B(\i43/i49/n361 ),
    .C(\i43/i49/n201 ),
    .Y(\i43/i49/n452 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i76  (.A(\i43/i49/n323 ),
    .B(\i43/i49/n381 ),
    .Y(\i43/i49/n451 ));
 NAND2xp33_ASAP7_75t_SL \i43/i49/i77  (.A(\i43/i49/n368 ),
    .B(\i43/i49/n389 ),
    .Y(\i43/i49/n437 ));
 NAND3xp33_ASAP7_75t_SL \i43/i49/i78  (.A(\i43/i49/n318 ),
    .B(\i43/i49/n355 ),
    .C(\i43/i49/n295 ),
    .Y(\i43/i49/n450 ));
 NAND2xp33_ASAP7_75t_SL \i43/i49/i79  (.A(\i43/i49/n370 ),
    .B(\i43/i49/n391 ),
    .Y(\i43/i49/n436 ));
 NAND4xp25_ASAP7_75t_SL \i43/i49/i8  (.A(\i43/i49/n486 ),
    .B(\i43/i49/n488 ),
    .C(\i43/i49/n475 ),
    .D(\i43/i49/n463 ),
    .Y(\i43/i49/n506 ));
 NAND2xp33_ASAP7_75t_SL \i43/i49/i80  (.A(\i43/i49/n406 ),
    .B(\i43/i49/n414 ),
    .Y(\i43/i49/n432 ));
 NAND4xp25_ASAP7_75t_SL \i43/i49/i81  (.A(\i43/i49/n323 ),
    .B(\i43/i49/n326 ),
    .C(\i43/i49/n294 ),
    .D(\i43/i49/n360 ),
    .Y(\i43/i49/n431 ));
 NAND3xp33_ASAP7_75t_SL \i43/i49/i82  (.A(\i43/i49/n322 ),
    .B(\i43/i49/n291 ),
    .C(\i43/i49/n276 ),
    .Y(\i43/i49/n430 ));
 NAND2xp5_ASAP7_75t_SL \i43/i49/i83  (.A(\i43/i49/n317 ),
    .B(\i43/i49/n385 ),
    .Y(\i43/i49/n429 ));
 NAND5xp2_ASAP7_75t_SL \i43/i49/i84  (.A(\i43/i49/n355 ),
    .B(\i43/i49/n214 ),
    .C(\i43/i49/n339 ),
    .D(\i43/i49/n235 ),
    .E(\i43/i49/n229 ),
    .Y(\i43/i49/n428 ));
 AOI211xp5_ASAP7_75t_SL \i43/i49/i85  (.A1(\i43/i49/n243 ),
    .A2(\i43/i49/n47 ),
    .B(\i43/i49/n284 ),
    .C(\i43/i49/n275 ),
    .Y(\i43/i49/n427 ));
 NOR2xp33_ASAP7_75t_L \i43/i49/i86  (.A(\i43/i49/n376 ),
    .B(\i43/i49/n409 ),
    .Y(\i43/i49/n426 ));
 NAND5xp2_ASAP7_75t_SL \i43/i49/i87  (.A(\i43/i49/n319 ),
    .B(\i43/i49/n367 ),
    .C(\i43/i49/n230 ),
    .D(\i43/i49/n127 ),
    .E(\i43/i49/n110 ),
    .Y(\i43/i49/n425 ));
 NAND4xp25_ASAP7_75t_SL \i43/i49/i88  (.A(\i43/i49/n352 ),
    .B(\i43/i49/n366 ),
    .C(\i43/i49/n345 ),
    .D(\i43/i49/n285 ),
    .Y(\i43/i49/n424 ));
 NOR2xp33_ASAP7_75t_SL \i43/i49/i89  (.A(\i43/i49/n346 ),
    .B(\i43/i49/n373 ),
    .Y(\i43/i49/n423 ));
 NAND4xp25_ASAP7_75t_SL \i43/i49/i9  (.A(\i43/i49/n480 ),
    .B(\i43/i49/n497 ),
    .C(\i43/i49/n494 ),
    .D(\i43/i49/n456 ),
    .Y(\i43/i49/n505 ));
 NOR5xp2_ASAP7_75t_SL \i43/i49/i90  (.A(\i43/i49/n335 ),
    .B(\i43/i49/n338 ),
    .C(\i43/i49/n119 ),
    .D(\i43/i49/n152 ),
    .E(\i43/i49/n102 ),
    .Y(\i43/i49/n422 ));
 AOI221xp5_ASAP7_75t_SL \i43/i49/i91  (.A1(\i43/i49/n258 ),
    .A2(\i43/i49/n55 ),
    .B1(\i43/i49/n155 ),
    .B2(\i43/i49/n256 ),
    .C(\i43/i49/n211 ),
    .Y(\i43/i49/n421 ));
 NOR5xp2_ASAP7_75t_SL \i43/i49/i92  (.A(\i43/i49/n212 ),
    .B(\i43/i49/n270 ),
    .C(\i43/i49/n239 ),
    .D(\i43/i49/n218 ),
    .E(\i43/i49/n177 ),
    .Y(\i43/i49/n420 ));
 NOR5xp2_ASAP7_75t_SL \i43/i49/i93  (.A(\i43/i49/n314 ),
    .B(\i43/i49/n350 ),
    .C(\i43/i49/n340 ),
    .D(\i43/i49/n217 ),
    .E(\i43/i49/n223 ),
    .Y(\i43/i49/n419 ));
 AOI211xp5_ASAP7_75t_SL \i43/i49/i94  (.A1(\i43/i49/n0 ),
    .A2(\i43/i49/n38 ),
    .B(\i43/i49/n297 ),
    .C(\i43/i49/n289 ),
    .Y(\i43/i49/n418 ));
 NOR5xp2_ASAP7_75t_SL \i43/i49/i95  (.A(\i43/i49/n328 ),
    .B(\i43/i49/n274 ),
    .C(\i43/i49/n280 ),
    .D(\i43/i49/n124 ),
    .E(\i43/i49/n174 ),
    .Y(\i43/i49/n417 ));
 NOR2xp67_ASAP7_75t_SL \i43/i49/i96  (.A(\i43/i49/n402 ),
    .B(\i43/i49/n404 ),
    .Y(\i43/i49/n435 ));
 AO211x2_ASAP7_75t_SL \i43/i49/i97  (.A1(\i43/i49/n88 ),
    .A2(\i43/i49/n262 ),
    .B(\i43/i49/n234 ),
    .C(\i43/i49/n313 ),
    .Y(\i43/i49/n434 ));
 AOI21xp5_ASAP7_75t_SL \i43/i49/i98  (.A1(\i43/i49/n33 ),
    .A2(\i43/i49/n73 ),
    .B(\i43/i49/n511 ),
    .Y(\i43/i49/n433 ));
 INVx1_ASAP7_75t_SL \i43/i49/i99  (.A(\i43/i49/n412 ),
    .Y(\i43/i49/n413 ));
 INVxp67_ASAP7_75t_SL \i43/i490  (.A(net55),
    .Y(\i43/n142 ));
 INVxp67_ASAP7_75t_SL \i43/i491  (.A(net80),
    .Y(\i43/n141 ));
 INVxp67_ASAP7_75t_SL \i43/i492  (.A(net44),
    .Y(\i43/n140 ));
 INVxp67_ASAP7_75t_SL \i43/i493  (.A(net45),
    .Y(\i43/n139 ));
 INVxp67_ASAP7_75t_SL \i43/i494  (.A(net86),
    .Y(\i43/n138 ));
 INVxp67_ASAP7_75t_SL \i43/i495  (.A(net70),
    .Y(\i43/n137 ));
 INVxp67_ASAP7_75t_SL \i43/i496  (.A(net114),
    .Y(\i43/n136 ));
 INVxp67_ASAP7_75t_SL \i43/i497  (.A(net48),
    .Y(\i43/n135 ));
 INVxp67_ASAP7_75t_SL \i43/i498  (.A(net32),
    .Y(\i43/n134 ));
 INVxp67_ASAP7_75t_SL \i43/i499  (.A(net127),
    .Y(\i43/n133 ));
 INVx1_ASAP7_75t_SL \i43/i5  (.A(n37[25]),
    .Y(n44));
 DFFHQNx1_ASAP7_75t_L \i43/i50  (.CLK(clk),
    .D(\i43/n361 ),
    .QN(n37[0]));
 INVxp67_ASAP7_75t_SL \i43/i500  (.A(net76),
    .Y(\i43/n132 ));
 INVxp67_ASAP7_75t_SL \i43/i501  (.A(net52),
    .Y(\i43/n131 ));
 INVxp67_ASAP7_75t_SL \i43/i502  (.A(net65),
    .Y(\i43/n130 ));
 INVxp67_ASAP7_75t_SL \i43/i503  (.A(net50),
    .Y(\i43/n129 ));
 INVxp67_ASAP7_75t_SL \i43/i504  (.A(net105),
    .Y(\i43/n128 ));
 INVxp67_ASAP7_75t_SL \i43/i505  (.A(net62),
    .Y(\i43/n127 ));
 INVxp67_ASAP7_75t_SL \i43/i506  (.A(net122),
    .Y(\i43/n126 ));
 INVxp67_ASAP7_75t_SL \i43/i507  (.A(net90),
    .Y(\i43/n125 ));
 INVxp67_ASAP7_75t_SL \i43/i508  (.A(net67),
    .Y(\i43/n124 ));
 INVxp67_ASAP7_75t_SL \i43/i509  (.A(net18),
    .Y(\i43/n123 ));
 DFFHQNx1_ASAP7_75t_SL \i43/i51  (.CLK(clk),
    .D(\i43/n384 ),
    .QN(n37[1]));
 INVxp67_ASAP7_75t_SL \i43/i510  (.A(net69),
    .Y(\i43/n122 ));
 INVxp67_ASAP7_75t_SL \i43/i511  (.A(net51),
    .Y(\i43/n121 ));
 INVxp67_ASAP7_75t_SL \i43/i512  (.A(net95),
    .Y(\i43/n120 ));
 INVxp67_ASAP7_75t_SL \i43/i513  (.A(net123),
    .Y(\i43/n119 ));
 INVxp67_ASAP7_75t_SL \i43/i514  (.A(net1),
    .Y(\i43/n118 ));
 INVxp67_ASAP7_75t_SL \i43/i515  (.A(net66),
    .Y(\i43/n117 ));
 INVxp67_ASAP7_75t_SL \i43/i516  (.A(net59),
    .Y(\i43/n116 ));
 INVxp67_ASAP7_75t_SL \i43/i517  (.A(net112),
    .Y(\i43/n115 ));
 INVxp67_ASAP7_75t_SL \i43/i518  (.A(net106),
    .Y(\i43/n114 ));
 INVx1_ASAP7_75t_SL \i43/i519  (.A(net26),
    .Y(\i43/n113 ));
 DFFHQNx1_ASAP7_75t_SL \i43/i52  (.CLK(clk),
    .D(\i43/n383 ),
    .QN(n37[2]));
 INVxp67_ASAP7_75t_SL \i43/i520  (.A(net118),
    .Y(\i43/n112 ));
 INVxp67_ASAP7_75t_SL \i43/i521  (.A(net49),
    .Y(\i43/n111 ));
 INVxp67_ASAP7_75t_SL \i43/i522  (.A(net74),
    .Y(\i43/n110 ));
 INVxp67_ASAP7_75t_SL \i43/i523  (.A(net119),
    .Y(\i43/n109 ));
 INVxp67_ASAP7_75t_SL \i43/i524  (.A(net37),
    .Y(\i43/n108 ));
 INVxp67_ASAP7_75t_SL \i43/i525  (.A(net9),
    .Y(\i43/n107 ));
 INVxp67_ASAP7_75t_SL \i43/i526  (.A(net113),
    .Y(\i43/n106 ));
 INVxp67_ASAP7_75t_SL \i43/i527  (.A(net94),
    .Y(\i43/n105 ));
 INVxp67_ASAP7_75t_SL \i43/i528  (.A(net33),
    .Y(\i43/n104 ));
 INVxp67_ASAP7_75t_SL \i43/i529  (.A(net36),
    .Y(\i43/n103 ));
 SDFHx1_ASAP7_75t_SL \i43/i53  (.CLK(clk),
    .QN(n37[3]),
    .D(\i43/n133 ),
    .SE(n38),
    .SI(\i43/n252 ));
 INVxp67_ASAP7_75t_SL \i43/i530  (.A(net56),
    .Y(\i43/n102 ));
 INVxp67_ASAP7_75t_SL \i43/i531  (.A(net60),
    .Y(\i43/n101 ));
 INVxp67_ASAP7_75t_SL \i43/i532  (.A(net58),
    .Y(\i43/n100 ));
 INVxp67_ASAP7_75t_SL \i43/i533  (.A(net40),
    .Y(\i43/n99 ));
 INVxp67_ASAP7_75t_SL \i43/i534  (.A(net96),
    .Y(\i43/n98 ));
 INVxp67_ASAP7_75t_SL \i43/i535  (.A(net103),
    .Y(\i43/n97 ));
 INVxp67_ASAP7_75t_SL \i43/i536  (.A(net77),
    .Y(\i43/n96 ));
 INVxp67_ASAP7_75t_SL \i43/i537  (.A(net110),
    .Y(\i43/n95 ));
 INVxp67_ASAP7_75t_SL \i43/i538  (.A(net104),
    .Y(\i43/n94 ));
 INVxp67_ASAP7_75t_SL \i43/i539  (.A(net61),
    .Y(\i43/n93 ));
 DFFHQNx1_ASAP7_75t_SL \i43/i54  (.CLK(clk),
    .D(\i43/n382 ),
    .QN(n37[4]));
 INVxp67_ASAP7_75t_SL \i43/i540  (.A(net42),
    .Y(\i43/n92 ));
 INVxp67_ASAP7_75t_SL \i43/i541  (.A(net23),
    .Y(\i43/n91 ));
 INVx2_ASAP7_75t_SL \i43/i542  (.A(\i43/n0 [29]),
    .Y(\i43/n90 ));
 INVx1_ASAP7_75t_SL \i43/i543  (.A(\i43/n2 [27]),
    .Y(\i43/n89 ));
 INVx1_ASAP7_75t_SL \i43/i544  (.A(\i43/n2 [28]),
    .Y(\i43/n88 ));
 INVx1_ASAP7_75t_SL \i43/i545  (.A(\i43/n0 [10]),
    .Y(\i43/n87 ));
 INVx2_ASAP7_75t_SL \i43/i546  (.A(\i43/n0 [27]),
    .Y(\i43/n86 ));
 INVx1_ASAP7_75t_SL \i43/i547  (.A(\i43/n2 [25]),
    .Y(\i43/n85 ));
 INVxp67_ASAP7_75t_SL \i43/i548  (.A(\i43/n0 [12]),
    .Y(\i43/n84 ));
 INVx1_ASAP7_75t_SL \i43/i549  (.A(\i43/n0 [18]),
    .Y(\i43/n83 ));
 DFFHQNx1_ASAP7_75t_SL \i43/i55  (.CLK(clk),
    .D(\i43/n381 ),
    .QN(n37[5]));
 INVx1_ASAP7_75t_SL \i43/i550  (.A(\i43/n2 [29]),
    .Y(\i43/n82 ));
 INVx1_ASAP7_75t_SL \i43/i551  (.A(\i43/n0 [28]),
    .Y(\i43/n81 ));
 INVx1_ASAP7_75t_SL \i43/i552  (.A(\i43/n2 [30]),
    .Y(\i43/n80 ));
 INVx1_ASAP7_75t_SL \i43/i553  (.A(\i43/n2 [26]),
    .Y(\i43/n79 ));
 INVxp67_ASAP7_75t_SL \i43/i554  (.A(\i43/n0 [20]),
    .Y(\i43/n78 ));
 INVx1_ASAP7_75t_SL \i43/i555  (.A(\i43/n0 [30]),
    .Y(\i43/n77 ));
 INVx1_ASAP7_75t_SL \i43/i556  (.A(\i43/n0 [26]),
    .Y(\i43/n76 ));
 INVx1_ASAP7_75t_SL \i43/i557  (.A(\i43/n0 [21]),
    .Y(\i43/n75 ));
 INVx1_ASAP7_75t_SL \i43/i558  (.A(\i43/n0 [2]),
    .Y(\i43/n74 ));
 INVx1_ASAP7_75t_SL \i43/i559  (.A(\i43/n0 [25]),
    .Y(\i43/n73 ));
 DFFHQNx1_ASAP7_75t_SL \i43/i56  (.CLK(clk),
    .D(\i43/n380 ),
    .QN(n37[6]));
 XNOR2xp5_ASAP7_75t_SL \i43/i560  (.A(\i43/n288 ),
    .B(\i43/n0 [23]),
    .Y(\i43/n67 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i561  (.A(\i43/n287 ),
    .B(\i43/n0 [22]),
    .Y(\i43/n66 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i562  (.A(\i43/n283 ),
    .B(\i43/n0 [14]),
    .Y(\i43/n65 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i563  (.A(\i43/n281 ),
    .B(\i43/n0 [15]),
    .Y(\i43/n64 ));
 XNOR2xp5_ASAP7_75t_SL \i43/i564  (.A(\i43/n271 ),
    .B(\i43/n0 [7]),
    .Y(\i43/n63 ));
 XOR2xp5_ASAP7_75t_SL \i43/i565  (.A(\i43/n262 ),
    .B(\i43/n41 ),
    .Y(\i43/n62 ));
 XOR2xp5_ASAP7_75t_SL \i43/i566  (.A(\i43/n256 ),
    .B(\i43/n194 ),
    .Y(\i43/n61 ));
 XOR2xp5_ASAP7_75t_SL \i43/i567  (.A(\i43/n254 ),
    .B(n36[10]),
    .Y(\i43/n60 ));
 XOR2xp5_ASAP7_75t_SL \i43/i568  (.A(\i43/n217 ),
    .B(\i43/n253 ),
    .Y(\i43/n59 ));
 XOR2xp5_ASAP7_75t_SL \i43/i569  (.A(\i43/n251 ),
    .B(n36[2]),
    .Y(\i43/n58 ));
 DFFHQNx1_ASAP7_75t_SL \i43/i57  (.CLK(clk),
    .D(\i43/n379 ),
    .QN(n37[7]));
 XNOR2xp5_ASAP7_75t_SL \i43/i570  (.A(\i43/n224 ),
    .B(\i43/n0 [6]),
    .Y(\i43/n57 ));
 XOR2xp5_ASAP7_75t_SL \i43/i571  (.A(\i43/n211 ),
    .B(\i43/n204 ),
    .Y(\i43/n56 ));
 XOR2xp5_ASAP7_75t_SL \i43/i572  (.A(\i43/n208 ),
    .B(\i43/n201 ),
    .Y(\i43/n55 ));
 XOR2xp5_ASAP7_75t_SL \i43/i573  (.A(\i43/n202 ),
    .B(n36[18]),
    .Y(\i43/n54 ));
 XOR2xp5_ASAP7_75t_SL \i43/i574  (.A(n37[17]),
    .B(\i43/n0 [17]),
    .Y(\i43/n53 ));
 XOR2xp5_ASAP7_75t_SL \i43/i575  (.A(n37[23]),
    .B(\i43/n0 [23]),
    .Y(\i43/n52 ));
 XOR2xp5_ASAP7_75t_SL \i43/i576  (.A(n37[15]),
    .B(\i43/n0 [15]),
    .Y(\i43/n51 ));
 XOR2xp5_ASAP7_75t_SL \i43/i577  (.A(n37[4]),
    .B(\i43/n0 [4]),
    .Y(\i43/n50 ));
 XOR2xp5_ASAP7_75t_SL \i43/i578  (.A(n37[7]),
    .B(\i43/n0 [7]),
    .Y(\i43/n49 ));
 XOR2xp5_ASAP7_75t_SL \i43/i579  (.A(n37[11]),
    .B(\i43/n0 [11]),
    .Y(\i43/n48 ));
 DFFHQNx1_ASAP7_75t_L \i43/i58  (.CLK(clk),
    .D(\i43/n378 ),
    .QN(n37[8]));
 XOR2xp5_ASAP7_75t_SL \i43/i580  (.A(n37[14]),
    .B(\i43/n0 [14]),
    .Y(\i43/n47 ));
 XOR2xp5_ASAP7_75t_SL \i43/i581  (.A(n37[19]),
    .B(\i43/n0 [19]),
    .Y(\i43/n46 ));
 XOR2xp5_ASAP7_75t_SL \i43/i582  (.A(n37[9]),
    .B(\i43/n0 [9]),
    .Y(\i43/n45 ));
 XOR2xp5_ASAP7_75t_SL \i43/i583  (.A(n37[3]),
    .B(\i43/n0 [3]),
    .Y(\i43/n44 ));
 XOR2xp5_ASAP7_75t_SL \i43/i584  (.A(n37[22]),
    .B(\i43/n0 [22]),
    .Y(\i43/n43 ));
 XOR2xp5_ASAP7_75t_SL \i43/i585  (.A(n37[1]),
    .B(\i43/n0 [1]),
    .Y(\i43/n42 ));
 XOR2x2_ASAP7_75t_SL \i43/i586  (.A(\i43/n2 [31]),
    .B(\i43/n0 [31]),
    .Y(\i43/n41 ));
 XOR2xp5_ASAP7_75t_SL \i43/i587  (.A(\i43/n255 ),
    .B(\i43/n189 ),
    .Y(\i43/n450 ));
 FAx1_ASAP7_75t_SL \i43/i588  (.SN(\i43/n451 ),
    .A(\i43/n246 ),
    .B(\i43/n2 [29]),
    .CI(\i43/n238 ),
    .CON(\i43/n27 ));
 FAx1_ASAP7_75t_SL \i43/i589  (.SN(\i43/n452 ),
    .A(\i43/n244 ),
    .B(\i43/n2 [31]),
    .CI(\i43/n236 ),
    .CON(\i43/n28 ));
 DFFHQNx1_ASAP7_75t_SL \i43/i59  (.CLK(clk),
    .D(\i43/n377 ),
    .QN(n37[9]));
 FAx1_ASAP7_75t_SL \i43/i590  (.SN(\i43/n453 ),
    .A(\i43/n289 ),
    .B(\i43/n0 [1]),
    .CI(\i43/n206 ),
    .CON(\i43/n29 ));
 FAx1_ASAP7_75t_SL \i43/i591  (.SN(\i43/n454 ),
    .A(\i43/n272 ),
    .B(\i43/n0 [3]),
    .CI(\i43/n220 ),
    .CON(\i43/n30 ));
 FAx1_ASAP7_75t_SL \i43/i592  (.SN(\i43/n455 ),
    .A(\i43/n228 ),
    .B(\i43/n0 [4]),
    .CI(\i43/n218 ),
    .CON(\i43/n31 ));
 FAx1_ASAP7_75t_SL \i43/i593  (.SN(\i43/n456 ),
    .A(\i43/n275 ),
    .B(\i43/n0 [9]),
    .CI(\i43/n209 ),
    .CON(\i43/n32 ));
 FAx1_ASAP7_75t_SL \i43/i594  (.SN(\i43/n457 ),
    .A(\i43/n276 ),
    .B(\i43/n0 [11]),
    .CI(\i43/n223 ),
    .CON(\i43/n33 ));
 FAx1_ASAP7_75t_SL \i43/i595  (.SN(\i43/n458 ),
    .A(\i43/n225 ),
    .B(\i43/n0 [12]),
    .CI(\i43/n205 ),
    .CON(\i43/n34 ));
 FAx1_ASAP7_75t_SL \i43/i596  (.SN(\i43/n459 ),
    .A(\i43/n282 ),
    .B(\i43/n0 [17]),
    .CI(\i43/n210 ),
    .CON(\i43/n35 ));
 FAx1_ASAP7_75t_SL \i43/i597  (.SN(\i43/n460 ),
    .A(\i43/n284 ),
    .B(\i43/n0 [19]),
    .CI(\i43/n216 ),
    .CON(\i43/n36 ));
 FAx1_ASAP7_75t_SL \i43/i598  (.SN(\i43/n461 ),
    .A(\i43/n235 ),
    .B(\i43/n0 [20]),
    .CI(\i43/n221 ),
    .CON(\i43/n37 ));
 FAx1_ASAP7_75t_SL \i43/i599  (.SN(\i43/n462 ),
    .A(\i43/n2 [26]),
    .B(n35[26]),
    .CI(n43),
    .CON(\i43/n38 ));
 INVx1_ASAP7_75t_SL \i43/i6  (.A(n37[21]),
    .Y(n45));
 DFFHQNx1_ASAP7_75t_SL \i43/i60  (.CLK(clk),
    .D(\i43/n376 ),
    .QN(n37[10]));
 FAx1_ASAP7_75t_SL \i43/i600  (.SN(\i43/n463 ),
    .A(\i43/n165 ),
    .B(n35[27]),
    .CI(\i43/n2 [27]),
    .CON(\i43/n39 ));
 FAx1_ASAP7_75t_SL \i43/i601  (.SN(\i43/n464 ),
    .A(n37[28]),
    .B(n35[28]),
    .CI(\i43/n2 [28]),
    .CON(\i43/n40 ));
 SDFHx1_ASAP7_75t_SL \i43/i61  (.CLK(clk),
    .QN(n37[11]),
    .D(\i43/n107 ),
    .SE(n38),
    .SI(\i43/n200 ));
 DFFHQNx1_ASAP7_75t_SL \i43/i62  (.CLK(clk),
    .D(\i43/n372 ),
    .QN(n37[12]));
 DFFHQNx1_ASAP7_75t_SL \i43/i63  (.CLK(clk),
    .D(\i43/n375 ),
    .QN(n37[13]));
 DFFHQNx1_ASAP7_75t_SL \i43/i64  (.CLK(clk),
    .D(\i43/n374 ),
    .QN(n37[14]));
 DFFHQNx1_ASAP7_75t_SL \i43/i65  (.CLK(clk),
    .D(\i43/n373 ),
    .QN(n37[15]));
 DFFHQNx1_ASAP7_75t_L \i43/i66  (.CLK(clk),
    .D(\i43/n371 ),
    .QN(n37[16]));
 DFFHQNx1_ASAP7_75t_SL \i43/i67  (.CLK(clk),
    .D(\i43/n369 ),
    .QN(n37[17]));
 DFFHQNx1_ASAP7_75t_SL \i43/i68  (.CLK(clk),
    .D(\i43/n370 ),
    .QN(n37[18]));
 SDFHx1_ASAP7_75t_SL \i43/i69  (.CLK(clk),
    .QN(n37[19]),
    .D(\i43/n123 ),
    .SE(n38),
    .SI(\i43/n203 ));
 INVx1_ASAP7_75t_SL \i43/i7  (.A(n37[20]),
    .Y(n46));
 DFFHQNx1_ASAP7_75t_SL \i43/i70  (.CLK(clk),
    .D(\i43/n368 ),
    .QN(n37[20]));
 DFFHQNx1_ASAP7_75t_SL \i43/i71  (.CLK(clk),
    .D(\i43/n367 ),
    .QN(n37[21]));
 DFFHQNx1_ASAP7_75t_SL \i43/i72  (.CLK(clk),
    .D(\i43/n366 ),
    .QN(n37[22]));
 DFFHQNx1_ASAP7_75t_SL \i43/i73  (.CLK(clk),
    .D(\i43/n365 ),
    .QN(n37[23]));
 DFFHQNx1_ASAP7_75t_SL \i43/i74  (.CLK(clk),
    .D(\i43/n421 ),
    .QN(n37[24]));
 DFFHQNx2_ASAP7_75t_SL \i43/i75  (.CLK(clk),
    .D(\i43/n426 ),
    .QN(n37[25]));
 SDFHx1_ASAP7_75t_L \i43/i76  (.CLK(clk),
    .QN(n37[26]),
    .D(\i43/n113 ),
    .SE(n38),
    .SI(\i43/n320 ));
 DFFHQNx1_ASAP7_75t_L \i43/i77  (.CLK(clk),
    .D(\i43/n427 ),
    .QN(n37[27]));
 DFFHQNx2_ASAP7_75t_SL \i43/i78  (.CLK(clk),
    .D(\i43/n425 ),
    .QN(n37[28]));
 DFFHQNx1_ASAP7_75t_L \i43/i79  (.CLK(clk),
    .D(\i43/n413 ),
    .QN(n37[29]));
 INVx1_ASAP7_75t_SL \i43/i8  (.A(n37[18]),
    .Y(n47));
 DFFHQNx1_ASAP7_75t_L \i43/i80  (.CLK(clk),
    .D(\i43/n436 ),
    .QN(n37[30]));
 DFFHQNx1_ASAP7_75t_L \i43/i81  (.CLK(clk),
    .D(\i43/n435 ),
    .QN(n37[31]));
 DFFHQNx1_ASAP7_75t_SL \i43/i82  (.CLK(clk),
    .D(\i43/n434 ),
    .QN(n36[0]));
 SDFHx1_ASAP7_75t_SL \i43/i83  (.CLK(clk),
    .QN(n36[1]),
    .D(\i43/n125 ),
    .SE(n38),
    .SI(\i43/n362 ));
 DFFHQNx1_ASAP7_75t_L \i43/i84  (.CLK(clk),
    .D(\i43/n433 ),
    .QN(n36[2]));
 SDFHx1_ASAP7_75t_SL \i43/i85  (.CLK(clk),
    .QN(n36[3]),
    .D(\i43/n148 ),
    .SE(n38),
    .SI(\i43/n360 ));
 SDFHx1_ASAP7_75t_SL \i43/i86  (.CLK(clk),
    .QN(n36[4]),
    .D(\i43/n150 ),
    .SE(n38),
    .SI(\i43/n359 ));
 SDFHx1_ASAP7_75t_SL \i43/i87  (.CLK(clk),
    .QN(n36[5]),
    .D(\i43/n105 ),
    .SE(n38),
    .SI(\i43/n358 ));
 SDFHx1_ASAP7_75t_SL \i43/i88  (.CLK(clk),
    .QN(n36[6]),
    .D(\i43/n98 ),
    .SE(n38),
    .SI(\i43/n357 ));
 SDFHx1_ASAP7_75t_SL \i43/i89  (.CLK(clk),
    .QN(n36[7]),
    .D(\i43/n146 ),
    .SE(n38),
    .SI(\i43/n356 ));
 INVx1_ASAP7_75t_SL \i43/i9  (.A(n37[13]),
    .Y(n48));
 DFFHQNx1_ASAP7_75t_SL \i43/i90  (.CLK(clk),
    .D(\i43/n432 ),
    .QN(n36[8]));
 SDFHx1_ASAP7_75t_SL \i43/i91  (.CLK(clk),
    .QN(n36[9]),
    .D(\i43/n173 ),
    .SE(n38),
    .SI(\i43/n355 ));
 DFFHQNx1_ASAP7_75t_L \i43/i92  (.CLK(clk),
    .D(\i43/n431 ),
    .QN(n36[10]));
 SDFHx1_ASAP7_75t_SL \i43/i93  (.CLK(clk),
    .QN(n36[11]),
    .D(\i43/n158 ),
    .SE(n38),
    .SI(\i43/n354 ));
 SDFHx1_ASAP7_75t_SL \i43/i94  (.CLK(clk),
    .QN(n36[12]),
    .D(\i43/n161 ),
    .SE(n38),
    .SI(\i43/n353 ));
 SDFHx1_ASAP7_75t_SL \i43/i95  (.CLK(clk),
    .QN(n36[13]),
    .D(\i43/n97 ),
    .SE(n38),
    .SI(\i43/n351 ));
 SDFHx1_ASAP7_75t_SL \i43/i96  (.CLK(clk),
    .QN(n36[14]),
    .D(\i43/n94 ),
    .SE(n38),
    .SI(\i43/n350 ));
 SDFHx1_ASAP7_75t_SL \i43/i97  (.CLK(clk),
    .QN(n36[15]),
    .D(\i43/n128 ),
    .SE(n38),
    .SI(\i43/n349 ));
 DFFHQNx1_ASAP7_75t_SL \i43/i98  (.CLK(clk),
    .D(\i43/n430 ),
    .QN(n36[16]));
 SDFHx1_ASAP7_75t_SL \i43/i99  (.CLK(clk),
    .QN(n36[17]),
    .D(\i43/n144 ),
    .SE(n38),
    .SI(\i43/n308 ));
 XNOR2xp5_ASAP7_75t_SL i430 (.A(n811),
    .B(n935),
    .Y(n1042));
 XNOR2xp5_ASAP7_75t_SL i431 (.A(n481),
    .B(n934),
    .Y(n1041));
 XOR2xp5_ASAP7_75t_SL i432 (.A(n887),
    .B(n933),
    .Y(n1040));
 XOR2xp5_ASAP7_75t_SL i433 (.A(n886),
    .B(n927),
    .Y(n1039));
 XNOR2xp5_ASAP7_75t_SL i434 (.A(n925),
    .B(n907),
    .Y(n1038));
 XOR2xp5_ASAP7_75t_SL i435 (.A(n772),
    .B(n926),
    .Y(n1037));
 XNOR2xp5_ASAP7_75t_SL i436 (.A(n475),
    .B(n998),
    .Y(n1036));
 XOR2xp5_ASAP7_75t_SL i437 (.A(n124),
    .B(n989),
    .Y(n1035));
 XOR2xp5_ASAP7_75t_SL i438 (.A(n124),
    .B(n986),
    .Y(n1034));
 XOR2xp5_ASAP7_75t_SL i439 (.A(n1163),
    .B(n974),
    .Y(n1033));
 INVxp67_ASAP7_75t_SL \i44/i0  (.A(n33[4]),
    .Y(\i44/n0 ));
 INVx2_ASAP7_75t_SL \i44/i1  (.A(n33[2]),
    .Y(\i44/n1 ));
 AND3x4_ASAP7_75t_SL \i44/i10  (.A(\i44/n525 ),
    .B(\i44/n534 ),
    .C(\i44/n513 ),
    .Y(n32[1]));
 NAND2xp33_ASAP7_75t_SL \i44/i100  (.A(\i44/n326 ),
    .B(\i44/n431 ),
    .Y(\i44/n449 ));
 NOR5xp2_ASAP7_75t_SL \i44/i101  (.A(\i44/n373 ),
    .B(\i44/n550 ),
    .C(\i44/n356 ),
    .D(\i44/n300 ),
    .E(\i44/n248 ),
    .Y(\i44/n448 ));
 NAND5xp2_ASAP7_75t_SL \i44/i102  (.A(\i44/n311 ),
    .B(\i44/n388 ),
    .C(\i44/n239 ),
    .D(\i44/n354 ),
    .E(\i44/n296 ),
    .Y(\i44/n447 ));
 NAND3xp33_ASAP7_75t_L \i44/i103  (.A(\i44/n305 ),
    .B(\i44/n339 ),
    .C(\i44/n415 ),
    .Y(\i44/n446 ));
 NOR5xp2_ASAP7_75t_SL \i44/i104  (.A(\i44/n304 ),
    .B(\i44/n317 ),
    .C(\i44/n294 ),
    .D(\i44/n130 ),
    .E(\i44/n106 ),
    .Y(\i44/n445 ));
 NAND5xp2_ASAP7_75t_SL \i44/i105  (.A(\i44/n28 ),
    .B(\i44/n561 ),
    .C(\i44/n239 ),
    .D(\i44/n103 ),
    .E(\i44/n214 ),
    .Y(\i44/n444 ));
 NAND4xp25_ASAP7_75t_SL \i44/i106  (.A(\i44/n242 ),
    .B(\i44/n256 ),
    .C(\i44/n360 ),
    .D(\i44/n21 ),
    .Y(\i44/n443 ));
 NOR5xp2_ASAP7_75t_SL \i44/i107  (.A(\i44/n262 ),
    .B(\i44/n560 ),
    .C(\i44/n247 ),
    .D(\i44/n208 ),
    .E(\i44/n206 ),
    .Y(\i44/n442 ));
 NOR2xp33_ASAP7_75t_SL \i44/i108  (.A(\i44/n404 ),
    .B(\i44/n436 ),
    .Y(\i44/n441 ));
 NOR2xp33_ASAP7_75t_SL \i44/i109  (.A(\i44/n392 ),
    .B(\i44/n423 ),
    .Y(\i44/n440 ));
 NOR2x1p5_ASAP7_75t_SL \i44/i11  (.A(\i44/n535 ),
    .B(\i44/n526 ),
    .Y(n32[5]));
 NAND3x1_ASAP7_75t_SL \i44/i110  (.A(\i44/n260 ),
    .B(\i44/n422 ),
    .C(\i44/n388 ),
    .Y(\i44/n457 ));
 NAND3x1_ASAP7_75t_SL \i44/i111  (.A(\i44/n383 ),
    .B(\i44/n361 ),
    .C(\i44/n327 ),
    .Y(\i44/n456 ));
 AOI21xp5_ASAP7_75t_L \i44/i112  (.A1(\i44/n78 ),
    .A2(\i44/n265 ),
    .B(\i44/n184 ),
    .Y(\i44/n433 ));
 NAND2xp5_ASAP7_75t_SL \i44/i113  (.A(\i44/n359 ),
    .B(\i44/n391 ),
    .Y(\i44/n432 ));
 NOR2xp33_ASAP7_75t_SL \i44/i114  (.A(\i44/n390 ),
    .B(\i44/n29 ),
    .Y(\i44/n431 ));
 NOR2xp33_ASAP7_75t_SL \i44/i115  (.A(\i44/n367 ),
    .B(\i44/n378 ),
    .Y(\i44/n430 ));
 NOR2xp67_ASAP7_75t_SL \i44/i116  (.A(\i44/n193 ),
    .B(\i44/n375 ),
    .Y(\i44/n429 ));
 NOR2xp33_ASAP7_75t_SL \i44/i117  (.A(\i44/n573 ),
    .B(\i44/n373 ),
    .Y(\i44/n428 ));
 NOR4xp25_ASAP7_75t_SL \i44/i118  (.A(\i44/n342 ),
    .B(\i44/n568 ),
    .C(\i44/n573 ),
    .D(\i44/n572 ),
    .Y(\i44/n427 ));
 NAND2xp5_ASAP7_75t_SL \i44/i119  (.A(\i44/n290 ),
    .B(\i44/n351 ),
    .Y(\i44/n426 ));
 AND2x2_ASAP7_75t_SL \i44/i12  (.A(\i44/n536 ),
    .B(\i44/n519 ),
    .Y(n32[0]));
 NOR4xp25_ASAP7_75t_SL \i44/i120  (.A(\i44/n126 ),
    .B(\i44/n283 ),
    .C(\i44/n250 ),
    .D(\i44/n266 ),
    .Y(\i44/n425 ));
 NOR3xp33_ASAP7_75t_SL \i44/i121  (.A(\i44/n288 ),
    .B(\i44/n241 ),
    .C(\i44/n287 ),
    .Y(\i44/n424 ));
 NAND2xp33_ASAP7_75t_SL \i44/i122  (.A(\i44/n338 ),
    .B(\i44/n26 ),
    .Y(\i44/n423 ));
 NOR2x1p5_ASAP7_75t_SL \i44/i123  (.A(\i44/n312 ),
    .B(\i44/n337 ),
    .Y(\i44/n422 ));
 NAND2xp33_ASAP7_75t_SL \i44/i124  (.A(\i44/n389 ),
    .B(\i44/n371 ),
    .Y(\i44/n421 ));
 NAND3xp33_ASAP7_75t_SL \i44/i125  (.A(\i44/n27 ),
    .B(\i44/n240 ),
    .C(\i44/n272 ),
    .Y(\i44/n420 ));
 NOR3xp33_ASAP7_75t_SL \i44/i126  (.A(\i44/n243 ),
    .B(\i44/n257 ),
    .C(\i44/n222 ),
    .Y(\i44/n439 ));
 NAND2xp5_ASAP7_75t_SL \i44/i127  (.A(\i44/n15 ),
    .B(\i44/n242 ),
    .Y(\i44/n438 ));
 NOR2x1_ASAP7_75t_SL \i44/i128  (.A(\i44/n310 ),
    .B(\i44/n335 ),
    .Y(\i44/n437 ));
 NAND2xp5_ASAP7_75t_SL \i44/i129  (.A(\i44/n239 ),
    .B(\i44/n343 ),
    .Y(\i44/n436 ));
 NOR3xp33_ASAP7_75t_SL \i44/i13  (.A(\i44/n508 ),
    .B(\i44/n504 ),
    .C(\i44/n511 ),
    .Y(\i44/n536 ));
 NOR2x1_ASAP7_75t_SL \i44/i130  (.A(\i44/n313 ),
    .B(\i44/n376 ),
    .Y(\i44/n435 ));
 NOR3x1_ASAP7_75t_SL \i44/i131  (.A(\i44/n247 ),
    .B(\i44/n237 ),
    .C(\i44/n204 ),
    .Y(\i44/n434 ));
 INVx1_ASAP7_75t_SL \i44/i132  (.A(\i44/n417 ),
    .Y(\i44/n418 ));
 INVx1_ASAP7_75t_SL \i44/i133  (.A(\i44/n30 ),
    .Y(\i44/n416 ));
 NOR4xp25_ASAP7_75t_SL \i44/i134  (.A(\i44/n226 ),
    .B(\i44/n269 ),
    .C(\i44/n255 ),
    .D(\i44/n220 ),
    .Y(\i44/n415 ));
 AOI211xp5_ASAP7_75t_SL \i44/i135  (.A1(\i44/n77 ),
    .A2(\i44/n72 ),
    .B(\i44/n337 ),
    .C(\i44/n199 ),
    .Y(\i44/n414 ));
 AOI211xp5_ASAP7_75t_SL \i44/i136  (.A1(\i44/n133 ),
    .A2(\i44/n61 ),
    .B(\i44/n355 ),
    .C(\i44/n286 ),
    .Y(\i44/n413 ));
 NAND2xp33_ASAP7_75t_L \i44/i137  (.A(\i44/n328 ),
    .B(\i44/n353 ),
    .Y(\i44/n412 ));
 NAND5xp2_ASAP7_75t_SL \i44/i138  (.A(\i44/n267 ),
    .B(\i44/n281 ),
    .C(\i44/n292 ),
    .D(\i44/n201 ),
    .E(\i44/n127 ),
    .Y(\i44/n411 ));
 NOR4xp25_ASAP7_75t_SL \i44/i139  (.A(\i44/n363 ),
    .B(\i44/n165 ),
    .C(\i44/n167 ),
    .D(\i44/n189 ),
    .Y(\i44/n410 ));
 NOR2x2_ASAP7_75t_SL \i44/i14  (.A(\i44/n528 ),
    .B(\i44/n529 ),
    .Y(n32[2]));
 OAI221xp5_ASAP7_75t_SL \i44/i140  (.A1(\i44/n97 ),
    .A2(\i44/n131 ),
    .B1(\i44/n131 ),
    .B2(\i44/n18 ),
    .C(\i44/n338 ),
    .Y(\i44/n409 ));
 NOR2xp33_ASAP7_75t_SL \i44/i141  (.A(\i44/n318 ),
    .B(\i44/n322 ),
    .Y(\i44/n408 ));
 AOI211xp5_ASAP7_75t_SL \i44/i142  (.A1(\i44/n187 ),
    .A2(\i44/n79 ),
    .B(\i44/n302 ),
    .C(\i44/n210 ),
    .Y(\i44/n407 ));
 OA21x2_ASAP7_75t_SL \i44/i143  (.A1(\i44/n537 ),
    .A2(\i44/n78 ),
    .B(\i44/n561 ),
    .Y(\i44/n406 ));
 NOR4xp25_ASAP7_75t_SL \i44/i144  (.A(\i44/n295 ),
    .B(\i44/n198 ),
    .C(\i44/n232 ),
    .D(\i44/n204 ),
    .Y(\i44/n405 ));
 NAND5xp2_ASAP7_75t_SL \i44/i145  (.A(\i44/n166 ),
    .B(\i44/n113 ),
    .C(\i44/n178 ),
    .D(\i44/n169 ),
    .E(\i44/n105 ),
    .Y(\i44/n404 ));
 NOR3xp33_ASAP7_75t_SL \i44/i146  (.A(\i44/n336 ),
    .B(\i44/n200 ),
    .C(\i44/n102 ),
    .Y(\i44/n403 ));
 NAND2xp5_ASAP7_75t_SL \i44/i147  (.A(\i44/n316 ),
    .B(\i44/n28 ),
    .Y(\i44/n402 ));
 NAND5xp2_ASAP7_75t_SL \i44/i148  (.A(\i44/n238 ),
    .B(\i44/n120 ),
    .C(\i44/n230 ),
    .D(\i44/n219 ),
    .E(\i44/n218 ),
    .Y(\i44/n401 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i44/i149  (.A1(\i44/n82 ),
    .A2(\i44/n108 ),
    .B(\i44/n84 ),
    .C(\i44/n307 ),
    .Y(\i44/n400 ));
 NAND4xp75_ASAP7_75t_SL \i44/i15  (.A(\i44/n494 ),
    .B(\i44/n514 ),
    .C(\i44/n492 ),
    .D(\i44/n574 ),
    .Y(\i44/n535 ));
 NAND4xp25_ASAP7_75t_SL \i44/i150  (.A(\i44/n349 ),
    .B(\i44/n282 ),
    .C(\i44/n128 ),
    .D(\i44/n202 ),
    .Y(\i44/n399 ));
 NAND5xp2_ASAP7_75t_SL \i44/i151  (.A(\i44/n188 ),
    .B(\i44/n168 ),
    .C(\i44/n274 ),
    .D(\i44/n123 ),
    .E(\i44/n117 ),
    .Y(\i44/n398 ));
 NAND2xp5_ASAP7_75t_SL \i44/i152  (.A(\i44/n315 ),
    .B(\i44/n341 ),
    .Y(\i44/n397 ));
 NAND3xp33_ASAP7_75t_SL \i44/i153  (.A(\i44/n334 ),
    .B(\i44/n104 ),
    .C(\i44/n110 ),
    .Y(\i44/n396 ));
 NAND2xp5_ASAP7_75t_SL \i44/i154  (.A(\i44/n260 ),
    .B(\i44/n388 ),
    .Y(\i44/n395 ));
 NOR2xp33_ASAP7_75t_L \i44/i155  (.A(\i44/n365 ),
    .B(\i44/n378 ),
    .Y(\i44/n419 ));
 NAND2xp5_ASAP7_75t_SL \i44/i156  (.A(\i44/n261 ),
    .B(\i44/n389 ),
    .Y(\i44/n394 ));
 NOR2x1p5_ASAP7_75t_SL \i44/i157  (.A(\i44/n320 ),
    .B(\i44/n369 ),
    .Y(\i44/n417 ));
 NAND3x1_ASAP7_75t_SL \i44/i158  (.A(\i44/n299 ),
    .B(\i44/n159 ),
    .C(\i44/n172 ),
    .Y(\i44/n30 ));
 INVxp67_ASAP7_75t_SL \i44/i159  (.A(\i44/n392 ),
    .Y(\i44/n393 ));
 NOR3xp33_ASAP7_75t_SL \i44/i16  (.A(\i44/n512 ),
    .B(\i44/n477 ),
    .C(\i44/n522 ),
    .Y(\i44/n534 ));
 INVxp67_ASAP7_75t_SL \i44/i160  (.A(\i44/n8 ),
    .Y(\i44/n391 ));
 INVxp67_ASAP7_75t_SL \i44/i161  (.A(\i44/n386 ),
    .Y(\i44/n387 ));
 INVxp67_ASAP7_75t_SL \i44/i162  (.A(\i44/n384 ),
    .Y(\i44/n385 ));
 INVx2_ASAP7_75t_SL \i44/i163  (.A(\i44/n382 ),
    .Y(\i44/n383 ));
 INVxp67_ASAP7_75t_SL \i44/i164  (.A(\i44/n380 ),
    .Y(\i44/n381 ));
 INVxp67_ASAP7_75t_SL \i44/i165  (.A(\i44/n376 ),
    .Y(\i44/n377 ));
 INVxp67_ASAP7_75t_SL \i44/i166  (.A(\i44/n567 ),
    .Y(\i44/n374 ));
 INVx1_ASAP7_75t_SL \i44/i167  (.A(\i44/n371 ),
    .Y(\i44/n372 ));
 OAI31xp33_ASAP7_75t_SL \i44/i168  (.A1(\i44/n79 ),
    .A2(\i44/n3 ),
    .A3(\i44/n62 ),
    .B(\i44/n58 ),
    .Y(\i44/n370 ));
 NAND2x1_ASAP7_75t_SL \i44/i169  (.A(\i44/n254 ),
    .B(\i44/n252 ),
    .Y(\i44/n369 ));
 NAND4xp75_ASAP7_75t_SL \i44/i17  (.A(\i44/n493 ),
    .B(\i44/n524 ),
    .C(\i44/n498 ),
    .D(\i44/n488 ),
    .Y(\i44/n533 ));
 NOR2xp33_ASAP7_75t_SL \i44/i170  (.A(\i44/n293 ),
    .B(\i44/n288 ),
    .Y(\i44/n368 ));
 NAND2xp33_ASAP7_75t_SL \i44/i171  (.A(\i44/n240 ),
    .B(\i44/n239 ),
    .Y(\i44/n367 ));
 OAI21xp5_ASAP7_75t_SL \i44/i172  (.A1(\i44/n60 ),
    .A2(\i44/n156 ),
    .B(\i44/n216 ),
    .Y(\i44/n366 ));
 NAND2xp5_ASAP7_75t_SL \i44/i173  (.A(\i44/n203 ),
    .B(\i44/n240 ),
    .Y(\i44/n365 ));
 AOI211xp5_ASAP7_75t_SL \i44/i174  (.A1(\i44/n95 ),
    .A2(\i44/n35 ),
    .B(\i44/n135 ),
    .C(\i44/n141 ),
    .Y(\i44/n364 ));
 AOI31xp33_ASAP7_75t_SL \i44/i175  (.A1(\i44/n60 ),
    .A2(\i44/n19 ),
    .A3(\i44/n70 ),
    .B(\i44/n55 ),
    .Y(\i44/n363 ));
 NOR3xp33_ASAP7_75t_SL \i44/i176  (.A(\i44/n241 ),
    .B(\i44/n155 ),
    .C(\i44/n139 ),
    .Y(\i44/n362 ));
 NOR3xp33_ASAP7_75t_SL \i44/i177  (.A(\i44/n132 ),
    .B(\i44/n148 ),
    .C(\i44/n293 ),
    .Y(\i44/n361 ));
 OAI31xp33_ASAP7_75t_SL \i44/i178  (.A1(\i44/n56 ),
    .A2(\i44/n58 ),
    .A3(\i44/n75 ),
    .B(\i44/n95 ),
    .Y(\i44/n360 ));
 AOI221xp5_ASAP7_75t_SL \i44/i179  (.A1(\i44/n82 ),
    .A2(\i44/n98 ),
    .B1(\i44/n562 ),
    .B2(\i44/n71 ),
    .C(\i44/n221 ),
    .Y(\i44/n359 ));
 AND3x4_ASAP7_75t_SL \i44/i18  (.A(\i44/n515 ),
    .B(\i44/n530 ),
    .C(\i44/n520 ),
    .Y(n32[7]));
 OAI31xp33_ASAP7_75t_R \i44/i180  (.A1(\i44/n79 ),
    .A2(\i44/n80 ),
    .A3(\i44/n82 ),
    .B(\i44/n75 ),
    .Y(\i44/n358 ));
 AOI21xp5_ASAP7_75t_SL \i44/i181  (.A1(\i44/n184 ),
    .A2(\i44/n70 ),
    .B(\i44/n93 ),
    .Y(\i44/n392 ));
 AOI21xp5_ASAP7_75t_L \i44/i182  (.A1(\i44/n70 ),
    .A2(\i44/n194 ),
    .B(\i44/n92 ),
    .Y(\i44/n357 ));
 OAI221xp5_ASAP7_75t_SL \i44/i183  (.A1(\i44/n20 ),
    .A2(\i44/n97 ),
    .B1(\i44/n57 ),
    .B2(\i44/n63 ),
    .C(\i44/n249 ),
    .Y(\i44/n356 ));
 AOI21xp33_ASAP7_75t_SL \i44/i184  (.A1(\i44/n194 ),
    .A2(\i44/n539 ),
    .B(\i44/n81 ),
    .Y(\i44/n355 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i44/i185  (.A1(\i44/n90 ),
    .A2(\i44/n6 ),
    .B(\i44/n94 ),
    .C(\i44/n22 ),
    .Y(\i44/n354 ));
 NOR3xp33_ASAP7_75t_SL \i44/i186  (.A(\i44/n263 ),
    .B(\i44/n132 ),
    .C(\i44/n163 ),
    .Y(\i44/n353 ));
 NAND3xp33_ASAP7_75t_SL \i44/i187  (.A(\i44/n23 ),
    .B(\i44/n25 ),
    .C(\i44/n192 ),
    .Y(\i44/n352 ));
 AOI22xp5_ASAP7_75t_SL \i44/i188  (.A1(\i44/n66 ),
    .A2(\i44/n180 ),
    .B1(\i44/n71 ),
    .B2(\i44/n62 ),
    .Y(\i44/n351 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i44/i189  (.A1(\i44/n92 ),
    .A2(\i44/n538 ),
    .B(\i44/n74 ),
    .C(\i44/n136 ),
    .Y(\i44/n350 ));
 NAND4xp75_ASAP7_75t_SL \i44/i19  (.A(\i44/n497 ),
    .B(\i44/n578 ),
    .C(\i44/n506 ),
    .D(\i44/n523 ),
    .Y(\i44/n532 ));
 OAI21xp5_ASAP7_75t_SL \i44/i190  (.A1(\i44/n69 ),
    .A2(\i44/n549 ),
    .B(\i44/n79 ),
    .Y(\i44/n349 ));
 NAND4xp25_ASAP7_75t_SL \i44/i191  (.A(\i44/n207 ),
    .B(\i44/n202 ),
    .C(\i44/n170 ),
    .D(\i44/n173 ),
    .Y(\i44/n348 ));
 NAND2xp33_ASAP7_75t_SL \i44/i192  (.A(\i44/n276 ),
    .B(\i44/n162 ),
    .Y(\i44/n347 ));
 OAI211xp5_ASAP7_75t_SL \i44/i193  (.A1(\i44/n81 ),
    .A2(\i44/n73 ),
    .B(\i44/n175 ),
    .C(\i44/n179 ),
    .Y(\i44/n390 ));
 NOR2xp67_ASAP7_75t_SL \i44/i194  (.A(\i44/n559 ),
    .B(\i44/n294 ),
    .Y(\i44/n389 ));
 AOI21x1_ASAP7_75t_SL \i44/i195  (.A1(\i44/n62 ),
    .A2(\i44/n69 ),
    .B(\i44/n302 ),
    .Y(\i44/n388 ));
 NAND2xp5_ASAP7_75t_SL \i44/i196  (.A(\i44/n278 ),
    .B(\i44/n253 ),
    .Y(\i44/n29 ));
 NOR2xp33_ASAP7_75t_SL \i44/i197  (.A(\i44/n279 ),
    .B(\i44/n295 ),
    .Y(\i44/n386 ));
 OAI211xp5_ASAP7_75t_SL \i44/i198  (.A1(\i44/n70 ),
    .A2(\i44/n81 ),
    .B(\i44/n216 ),
    .C(\i44/n217 ),
    .Y(\i44/n384 ));
 OR2x2_ASAP7_75t_SL \i44/i199  (.A(\i44/n228 ),
    .B(\i44/n557 ),
    .Y(\i44/n382 ));
 INVx1_ASAP7_75t_SL \i44/i2  (.A(\i44/n468 ),
    .Y(\i44/n2 ));
 NAND2x1_ASAP7_75t_SL \i44/i20  (.A(\i44/n485 ),
    .B(\i44/n516 ),
    .Y(\i44/n531 ));
 AOI21xp5_ASAP7_75t_SL \i44/i200  (.A1(\i44/n80 ),
    .A2(\i44/n545 ),
    .B(\i44/n291 ),
    .Y(\i44/n380 ));
 OAI211xp5_ASAP7_75t_SL \i44/i201  (.A1(\i44/n97 ),
    .A2(\i44/n85 ),
    .B(\i44/n212 ),
    .C(\i44/n150 ),
    .Y(\i44/n379 ));
 NAND2xp5_ASAP7_75t_SL \i44/i202  (.A(\i44/n296 ),
    .B(\i44/n297 ),
    .Y(\i44/n378 ));
 NAND2xp5_ASAP7_75t_SL \i44/i203  (.A(\i44/n27 ),
    .B(\i44/n223 ),
    .Y(\i44/n376 ));
 NAND2xp5_ASAP7_75t_SL \i44/i204  (.A(\i44/n275 ),
    .B(\i44/n303 ),
    .Y(\i44/n375 ));
 NAND2xp5_ASAP7_75t_SL \i44/i205  (.A(\i44/n209 ),
    .B(\i44/n234 ),
    .Y(\i44/n373 ));
 NOR2x1_ASAP7_75t_SL \i44/i206  (.A(\i44/n277 ),
    .B(\i44/n248 ),
    .Y(\i44/n371 ));
 INVxp67_ASAP7_75t_SL \i44/i207  (.A(\i44/n342 ),
    .Y(\i44/n343 ));
 INVx1_ASAP7_75t_SL \i44/i208  (.A(\i44/n339 ),
    .Y(\i44/n340 ));
 INVx1_ASAP7_75t_SL \i44/i209  (.A(\i44/n334 ),
    .Y(\i44/n335 ));
 NOR2xp67_ASAP7_75t_SL \i44/i21  (.A(\i44/n517 ),
    .B(\i44/n478 ),
    .Y(\i44/n530 ));
 NAND4xp25_ASAP7_75t_SL \i44/i210  (.A(\i44/n129 ),
    .B(\i44/n151 ),
    .C(\i44/n136 ),
    .D(\i44/n134 ),
    .Y(\i44/n331 ));
 AOI31xp33_ASAP7_75t_SL \i44/i211  (.A1(\i44/n152 ),
    .A2(\i44/n78 ),
    .A3(\i44/n55 ),
    .B(\i44/n539 ),
    .Y(\i44/n330 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i44/i212  (.A1(\i44/n94 ),
    .A2(\i44/n59 ),
    .B(\i44/n75 ),
    .C(\i44/n157 ),
    .Y(\i44/n329 ));
 NOR4xp25_ASAP7_75t_SL \i44/i213  (.A(\i44/n126 ),
    .B(\i44/n142 ),
    .C(\i44/n215 ),
    .D(\i44/n101 ),
    .Y(\i44/n328 ));
 AOI211xp5_ASAP7_75t_SL \i44/i214  (.A1(\i44/n153 ),
    .A2(\i44/n546 ),
    .B(\i44/n200 ),
    .C(\i44/n111 ),
    .Y(\i44/n327 ));
 AOI21xp5_ASAP7_75t_SL \i44/i215  (.A1(\i44/n185 ),
    .A2(\i44/n94 ),
    .B(\i44/n268 ),
    .Y(\i44/n326 ));
 NOR2xp33_ASAP7_75t_L \i44/i216  (.A(\i44/n558 ),
    .B(\i44/n548 ),
    .Y(\i44/n325 ));
 OAI31xp33_ASAP7_75t_SL \i44/i217  (.A1(\i44/n66 ),
    .A2(\i44/n562 ),
    .A3(\i44/n95 ),
    .B(\i44/n545 ),
    .Y(\i44/n324 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i44/i218  (.A1(\i44/n81 ),
    .A2(\i44/n538 ),
    .B(\i44/n89 ),
    .C(\i44/n264 ),
    .Y(\i44/n323 ));
 OAI22xp5_ASAP7_75t_SL \i44/i219  (.A1(\i44/n85 ),
    .A2(\i44/n186 ),
    .B1(\i44/n73 ),
    .B2(\i44/n109 ),
    .Y(\i44/n322 ));
 NAND4xp75_ASAP7_75t_SL \i44/i22  (.A(\i44/n489 ),
    .B(\i44/n501 ),
    .C(\i44/n483 ),
    .D(\i44/n486 ),
    .Y(\i44/n529 ));
 NOR2xp33_ASAP7_75t_SL \i44/i220  (.A(\i44/n245 ),
    .B(\i44/n224 ),
    .Y(\i44/n321 ));
 OAI222xp33_ASAP7_75t_SL \i44/i221  (.A1(\i44/n92 ),
    .A2(\i44/n539 ),
    .B1(\i44/n538 ),
    .B2(\i44/n19 ),
    .C1(\i44/n78 ),
    .C2(\i44/n73 ),
    .Y(\i44/n320 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i44/i222  (.A1(\i44/n66 ),
    .A2(\i44/n64 ),
    .B(\i44/n6 ),
    .C(\i44/n196 ),
    .Y(\i44/n319 ));
 NAND2xp33_ASAP7_75t_L \i44/i223  (.A(\i44/n125 ),
    .B(\i44/n235 ),
    .Y(\i44/n318 ));
 NAND2xp33_ASAP7_75t_SL \i44/i224  (.A(\i44/n285 ),
    .B(\i44/n149 ),
    .Y(\i44/n317 ));
 AOI22xp33_ASAP7_75t_SL \i44/i225  (.A1(\i44/n80 ),
    .A2(\i44/n122 ),
    .B1(\i44/n546 ),
    .B2(\i44/n82 ),
    .Y(\i44/n316 ));
 OAI21xp33_ASAP7_75t_SL \i44/i226  (.A1(\i44/n133 ),
    .A2(\i44/n80 ),
    .B(\i44/n546 ),
    .Y(\i44/n315 ));
 OA21x2_ASAP7_75t_SL \i44/i227  (.A1(\i44/n539 ),
    .A2(\i44/n156 ),
    .B(\i44/n144 ),
    .Y(\i44/n314 ));
 NAND2xp5_ASAP7_75t_SL \i44/i228  (.A(\i44/n229 ),
    .B(\i44/n301 ),
    .Y(\i44/n313 ));
 NAND4xp25_ASAP7_75t_SL \i44/i229  (.A(\i44/n146 ),
    .B(\i44/n174 ),
    .C(\i44/n119 ),
    .D(\i44/n116 ),
    .Y(\i44/n312 ));
 OR3x1_ASAP7_75t_SL \i44/i23  (.A(\i44/n509 ),
    .B(\i44/n507 ),
    .C(\i44/n490 ),
    .Y(\i44/n528 ));
 AOI221xp5_ASAP7_75t_SL \i44/i230  (.A1(\i44/n71 ),
    .A2(\i44/n54 ),
    .B1(\i44/n59 ),
    .B2(\i44/n72 ),
    .C(\i44/n556 ),
    .Y(\i44/n311 ));
 OAI221xp5_ASAP7_75t_SL \i44/i231  (.A1(\i44/n96 ),
    .A2(\i44/n89 ),
    .B1(\i44/n76 ),
    .B2(\i44/n18 ),
    .C(\i44/n124 ),
    .Y(\i44/n346 ));
 OAI222xp33_ASAP7_75t_SL \i44/i232  (.A1(\i44/n9 ),
    .A2(\i44/n60 ),
    .B1(\i44/n63 ),
    .B2(\i44/n73 ),
    .C1(\i44/n76 ),
    .C2(\i44/n83 ),
    .Y(\i44/n310 ));
 OAI221xp5_ASAP7_75t_SL \i44/i233  (.A1(\i44/n92 ),
    .A2(\i44/n83 ),
    .B1(\i44/n76 ),
    .B2(\i44/n74 ),
    .C(\i44/n246 ),
    .Y(\i44/n309 ));
 AND3x1_ASAP7_75t_SL \i44/i234  (.A(\i44/n143 ),
    .B(\i44/n151 ),
    .C(\i44/n270 ),
    .Y(\i44/n308 ));
 AOI22xp5_ASAP7_75t_SL \i44/i235  (.A1(\i44/n91 ),
    .A2(\i44/n182 ),
    .B1(\i44/n69 ),
    .B2(\i44/n94 ),
    .Y(\i44/n345 ));
 NAND2xp33_ASAP7_75t_SL \i44/i236  (.A(\i44/n231 ),
    .B(\i44/n271 ),
    .Y(\i44/n307 ));
 OAI221xp5_ASAP7_75t_SL \i44/i237  (.A1(\i44/n92 ),
    .A2(\i44/n87 ),
    .B1(\i44/n20 ),
    .B2(\i44/n19 ),
    .C(\i44/n284 ),
    .Y(\i44/n306 ));
 OAI222xp33_ASAP7_75t_SL \i44/i238  (.A1(\i44/n85 ),
    .A2(\i44/n87 ),
    .B1(\i44/n96 ),
    .B2(\i44/n83 ),
    .C1(\i44/n20 ),
    .C2(\i44/n70 ),
    .Y(\i44/n344 ));
 NAND3x1_ASAP7_75t_SL \i44/i239  (.A(\i44/n236 ),
    .B(\i44/n177 ),
    .C(\i44/n171 ),
    .Y(\i44/n342 ));
 OR3x1_ASAP7_75t_SL \i44/i24  (.A(\i44/n510 ),
    .B(\i44/n476 ),
    .C(\i44/n450 ),
    .Y(\i44/n527 ));
 AOI22x1_ASAP7_75t_SL \i44/i240  (.A1(\i44/n176 ),
    .A2(\i44/n95 ),
    .B1(\i44/n562 ),
    .B2(\i44/n75 ),
    .Y(\i44/n15 ));
 AOI22xp5_ASAP7_75t_SL \i44/i241  (.A1(\i44/n98 ),
    .A2(\i44/n114 ),
    .B1(\i44/n56 ),
    .B2(\i44/n79 ),
    .Y(\i44/n341 ));
 AOI221x1_ASAP7_75t_SL \i44/i242  (.A1(\i44/n95 ),
    .A2(\i44/n75 ),
    .B1(\i44/n82 ),
    .B2(\i44/n84 ),
    .C(\i44/n273 ),
    .Y(\i44/n339 ));
 AOI211x1_ASAP7_75t_SL \i44/i243  (.A1(\i44/n115 ),
    .A2(\i44/n565 ),
    .B(\i44/n213 ),
    .C(\i44/n215 ),
    .Y(\i44/n338 ));
 AO21x2_ASAP7_75t_SL \i44/i244  (.A1(\i44/n546 ),
    .A2(\i44/n3 ),
    .B(\i44/n571 ),
    .Y(\i44/n337 ));
 OAI21xp5_ASAP7_75t_SL \i44/i245  (.A1(\i44/n55 ),
    .A2(\i44/n89 ),
    .B(\i44/n280 ),
    .Y(\i44/n336 ));
 NOR2x1_ASAP7_75t_SL \i44/i246  (.A(\i44/n145 ),
    .B(\i44/n227 ),
    .Y(\i44/n334 ));
 OAI211xp5_ASAP7_75t_SL \i44/i247  (.A1(\i44/n74 ),
    .A2(\i44/n118 ),
    .B(\i44/n128 ),
    .C(\i44/n158 ),
    .Y(\i44/n333 ));
 NOR2xp33_ASAP7_75t_SL \i44/i248  (.A(\i44/n157 ),
    .B(\i44/n233 ),
    .Y(\i44/n28 ));
 NOR2xp33_ASAP7_75t_SL \i44/i249  (.A(\i44/n160 ),
    .B(\i44/n298 ),
    .Y(\i44/n305 ));
 NAND3xp33_ASAP7_75t_SL \i44/i25  (.A(\i44/n521 ),
    .B(\i44/n506 ),
    .C(\i44/n489 ),
    .Y(\i44/n526 ));
 AOI222xp33_ASAP7_75t_SL \i44/i250  (.A1(\i44/n82 ),
    .A2(\i44/n71 ),
    .B1(\i44/n6 ),
    .B2(\i44/n54 ),
    .C1(\i44/n79 ),
    .C2(\i44/n69 ),
    .Y(\i44/n332 ));
 INVx1_ASAP7_75t_SL \i44/i251  (.A(\i44/n303 ),
    .Y(\i44/n304 ));
 INVx1_ASAP7_75t_SL \i44/i252  (.A(\i44/n300 ),
    .Y(\i44/n301 ));
 INVx1_ASAP7_75t_SL \i44/i253  (.A(\i44/n298 ),
    .Y(\i44/n299 ));
 INVxp67_ASAP7_75t_SL \i44/i254  (.A(\i44/n291 ),
    .Y(\i44/n292 ));
 INVx1_ASAP7_75t_SL \i44/i255  (.A(\i44/n548 ),
    .Y(\i44/n289 ));
 OAI21xp33_ASAP7_75t_SL \i44/i256  (.A1(\i44/n551 ),
    .A2(\i44/n68 ),
    .B(\i44/n205 ),
    .Y(\i44/n287 ));
 NAND2xp5_ASAP7_75t_SL \i44/i257  (.A(\i44/n107 ),
    .B(\i44/n150 ),
    .Y(\i44/n286 ));
 OAI21xp5_ASAP7_75t_SL \i44/i258  (.A1(\i44/n562 ),
    .A2(\i44/n62 ),
    .B(\i44/n90 ),
    .Y(\i44/n285 ));
 NOR2xp33_ASAP7_75t_SL \i44/i259  (.A(\i44/n161 ),
    .B(\i44/n199 ),
    .Y(\i44/n284 ));
 NOR2x1_ASAP7_75t_SL \i44/i26  (.A(\i44/n432 ),
    .B(\i44/n507 ),
    .Y(\i44/n524 ));
 NAND2xp33_ASAP7_75t_L \i44/i260  (.A(\i44/n195 ),
    .B(\i44/n112 ),
    .Y(\i44/n283 ));
 OAI21xp5_ASAP7_75t_SL \i44/i261  (.A1(\i44/n77 ),
    .A2(\i44/n64 ),
    .B(\i44/n58 ),
    .Y(\i44/n282 ));
 NOR2xp33_ASAP7_75t_SL \i44/i262  (.A(\i44/n22 ),
    .B(\i44/n137 ),
    .Y(\i44/n281 ));
 OAI21xp5_ASAP7_75t_SL \i44/i263  (.A1(\i44/n80 ),
    .A2(\i44/n88 ),
    .B(\i44/n71 ),
    .Y(\i44/n280 ));
 OAI21xp5_ASAP7_75t_SL \i44/i264  (.A1(\i44/n537 ),
    .A2(\i44/n93 ),
    .B(\i44/n197 ),
    .Y(\i44/n279 ));
 AOI22xp5_ASAP7_75t_SL \i44/i265  (.A1(\i44/n90 ),
    .A2(\i44/n64 ),
    .B1(\i44/n84 ),
    .B2(\i44/n79 ),
    .Y(\i44/n278 ));
 OAI21xp5_ASAP7_75t_SL \i44/i266  (.A1(\i44/n19 ),
    .A2(\i44/n76 ),
    .B(\i44/n154 ),
    .Y(\i44/n277 ));
 OAI21xp33_ASAP7_75t_SL \i44/i267  (.A1(\i44/n80 ),
    .A2(\i44/n62 ),
    .B(\i44/n72 ),
    .Y(\i44/n276 ));
 AOI22xp33_ASAP7_75t_SL \i44/i268  (.A1(\i44/n54 ),
    .A2(\i44/n98 ),
    .B1(\i44/n56 ),
    .B2(\i44/n80 ),
    .Y(\i44/n275 ));
 OAI21xp5_ASAP7_75t_SL \i44/i269  (.A1(\i44/n84 ),
    .A2(\i44/n98 ),
    .B(\i44/n91 ),
    .Y(\i44/n274 ));
 NOR2x1_ASAP7_75t_SL \i44/i27  (.A(\i44/n491 ),
    .B(\i44/n487 ),
    .Y(\i44/n523 ));
 OA21x2_ASAP7_75t_SL \i44/i270  (.A1(\i44/n6 ),
    .A2(\i44/n98 ),
    .B(\i44/n94 ),
    .Y(\i44/n273 ));
 AOI22xp33_ASAP7_75t_SL \i44/i271  (.A1(\i44/n98 ),
    .A2(\i44/n562 ),
    .B1(\i44/n565 ),
    .B2(\i44/n3 ),
    .Y(\i44/n272 ));
 OAI21xp5_ASAP7_75t_SL \i44/i272  (.A1(\i44/n72 ),
    .A2(\i44/n56 ),
    .B(\i44/n91 ),
    .Y(\i44/n271 ));
 OAI21xp5_ASAP7_75t_SL \i44/i273  (.A1(\i44/n80 ),
    .A2(\i44/n77 ),
    .B(\i44/n98 ),
    .Y(\i44/n270 ));
 AOI21xp33_ASAP7_75t_SL \i44/i274  (.A1(\i44/n70 ),
    .A2(\i44/n89 ),
    .B(\i44/n55 ),
    .Y(\i44/n269 ));
 OAI21xp5_ASAP7_75t_SL \i44/i275  (.A1(\i44/n537 ),
    .A2(\i44/n76 ),
    .B(\i44/n26 ),
    .Y(\i44/n268 ));
 AOI22xp5_ASAP7_75t_SL \i44/i276  (.A1(\i44/n69 ),
    .A2(\i44/n66 ),
    .B1(\i44/n84 ),
    .B2(\i44/n64 ),
    .Y(\i44/n267 ));
 AOI21xp33_ASAP7_75t_SL \i44/i277  (.A1(\i44/n81 ),
    .A2(\i44/n55 ),
    .B(\i44/n74 ),
    .Y(\i44/n266 ));
 OAI21xp33_ASAP7_75t_SL \i44/i278  (.A1(\i44/n94 ),
    .A2(\i44/n80 ),
    .B(\i44/n58 ),
    .Y(\i44/n265 ));
 OAI21xp5_ASAP7_75t_SL \i44/i279  (.A1(\i44/n77 ),
    .A2(\i44/n66 ),
    .B(\i44/n84 ),
    .Y(\i44/n264 ));
 NAND3xp33_ASAP7_75t_SL \i44/i28  (.A(\i44/n471 ),
    .B(\i44/n582 ),
    .C(\i44/n469 ),
    .Y(\i44/n522 ));
 NAND2xp5_ASAP7_75t_SL \i44/i280  (.A(\i44/n91 ),
    .B(\i44/n185 ),
    .Y(\i44/n27 ));
 AOI22xp5_ASAP7_75t_SL \i44/i281  (.A1(\i44/n100 ),
    .A2(\i44/n86 ),
    .B1(\i44/n84 ),
    .B2(\i44/n3 ),
    .Y(\i44/n303 ));
 NAND2xp5_ASAP7_75t_L \i44/i282  (.A(\i44/n216 ),
    .B(\i44/n217 ),
    .Y(\i44/n263 ));
 OAI22xp5_ASAP7_75t_SL \i44/i283  (.A1(\i44/n68 ),
    .A2(\i44/n92 ),
    .B1(\i44/n99 ),
    .B2(\i44/n17 ),
    .Y(\i44/n302 ));
 OAI22xp5_ASAP7_75t_L \i44/i284  (.A1(\i44/n99 ),
    .A2(\i44/n76 ),
    .B1(\i44/n20 ),
    .B2(\i44/n73 ),
    .Y(\i44/n300 ));
 OAI22xp5_ASAP7_75t_SL \i44/i285  (.A1(\i44/n97 ),
    .A2(\i44/n63 ),
    .B1(\i44/n537 ),
    .B2(\i44/n85 ),
    .Y(\i44/n298 ));
 AOI22xp5_ASAP7_75t_SL \i44/i286  (.A1(\i44/n565 ),
    .A2(\i44/n95 ),
    .B1(\i44/n6 ),
    .B2(\i44/n88 ),
    .Y(\i44/n297 ));
 AOI22xp5_ASAP7_75t_R \i44/i287  (.A1(\i44/n565 ),
    .A2(\i44/n66 ),
    .B1(\i44/n100 ),
    .B2(\i44/n64 ),
    .Y(\i44/n296 ));
 OAI22xp5_ASAP7_75t_SL \i44/i288  (.A1(\i44/n74 ),
    .A2(\i44/n85 ),
    .B1(\i44/n76 ),
    .B2(\i44/n57 ),
    .Y(\i44/n295 ));
 OAI22xp5_ASAP7_75t_SL \i44/i289  (.A1(\i44/n99 ),
    .A2(\i44/n96 ),
    .B1(\i44/n539 ),
    .B2(\i44/n9 ),
    .Y(\i44/n294 ));
 NOR2x1_ASAP7_75t_SL \i44/i29  (.A(\i44/n496 ),
    .B(\i44/n459 ),
    .Y(\i44/n521 ));
 NAND2xp5_ASAP7_75t_L \i44/i290  (.A(\i44/n21 ),
    .B(\i44/n181 ),
    .Y(\i44/n293 ));
 OAI22xp5_ASAP7_75t_SL \i44/i291  (.A1(\i44/n537 ),
    .A2(\i44/n96 ),
    .B1(\i44/n73 ),
    .B2(\i44/n93 ),
    .Y(\i44/n291 ));
 OAI21xp5_ASAP7_75t_SL \i44/i292  (.A1(\i44/n80 ),
    .A2(\i44/n59 ),
    .B(\i44/n90 ),
    .Y(\i44/n290 ));
 NAND2xp33_ASAP7_75t_L \i44/i293  (.A(\i44/n128 ),
    .B(\i44/n158 ),
    .Y(\i44/n262 ));
 OAI21xp5_ASAP7_75t_SL \i44/i294  (.A1(\i44/n74 ),
    .A2(\i44/n63 ),
    .B(\i44/n127 ),
    .Y(\i44/n288 ));
 INVxp67_ASAP7_75t_SL \i44/i295  (.A(\i44/n258 ),
    .Y(\i44/n259 ));
 INVxp67_ASAP7_75t_SL \i44/i296  (.A(\i44/n256 ),
    .Y(\i44/n257 ));
 INVx1_ASAP7_75t_SL \i44/i297  (.A(\i44/n254 ),
    .Y(\i44/n255 ));
 INVx1_ASAP7_75t_SL \i44/i298  (.A(\i44/n251 ),
    .Y(\i44/n252 ));
 INVxp67_ASAP7_75t_SL \i44/i299  (.A(\i44/n249 ),
    .Y(\i44/n250 ));
 INVx2_ASAP7_75t_SL \i44/i3  (.A(\i44/n9 ),
    .Y(\i44/n3 ));
 NOR5xp2_ASAP7_75t_SL \i44/i30  (.A(\i44/n461 ),
    .B(\i44/n411 ),
    .C(\i44/n452 ),
    .D(\i44/n375 ),
    .E(\i44/n379 ),
    .Y(\i44/n520 ));
 INVxp67_ASAP7_75t_SL \i44/i300  (.A(\i44/n245 ),
    .Y(\i44/n246 ));
 INVxp67_ASAP7_75t_SL \i44/i301  (.A(\i44/n243 ),
    .Y(\i44/n244 ));
 OAI21xp5_ASAP7_75t_SL \i44/i302  (.A1(\i44/n64 ),
    .A2(\i44/n86 ),
    .B(\i44/n84 ),
    .Y(\i44/n238 ));
 OAI21xp5_ASAP7_75t_SL \i44/i303  (.A1(\i44/n18 ),
    .A2(\i44/n9 ),
    .B(\i44/n140 ),
    .Y(\i44/n237 ));
 OAI21xp5_ASAP7_75t_SL \i44/i304  (.A1(\i44/n65 ),
    .A2(\i44/n75 ),
    .B(\i44/n77 ),
    .Y(\i44/n236 ));
 OAI21xp33_ASAP7_75t_SL \i44/i305  (.A1(\i44/n562 ),
    .A2(\i44/n59 ),
    .B(\i44/n65 ),
    .Y(\i44/n235 ));
 AOI22xp5_ASAP7_75t_SL \i44/i306  (.A1(\i44/n546 ),
    .A2(\i44/n66 ),
    .B1(\i44/n58 ),
    .B2(\i44/n3 ),
    .Y(\i44/n234 ));
 OAI22xp5_ASAP7_75t_SL \i44/i307  (.A1(\i44/n96 ),
    .A2(\i44/n60 ),
    .B1(\i44/n57 ),
    .B2(\i44/n17 ),
    .Y(\i44/n233 ));
 AOI21xp33_ASAP7_75t_SL \i44/i308  (.A1(\i44/n76 ),
    .A2(\i44/n85 ),
    .B(\i44/n87 ),
    .Y(\i44/n232 ));
 OAI21xp5_ASAP7_75t_SL \i44/i309  (.A1(\i44/n54 ),
    .A2(\i44/n59 ),
    .B(\i44/n58 ),
    .Y(\i44/n231 ));
 NOR3xp33_ASAP7_75t_SL \i44/i31  (.A(\i44/n457 ),
    .B(\i44/n473 ),
    .C(\i44/n505 ),
    .Y(\i44/n519 ));
 OAI21xp5_ASAP7_75t_SL \i44/i310  (.A1(\i44/n546 ),
    .A2(\i44/n65 ),
    .B(\i44/n562 ),
    .Y(\i44/n230 ));
 AOI22xp33_ASAP7_75t_SL \i44/i311  (.A1(\i44/n565 ),
    .A2(\i44/n80 ),
    .B1(\i44/n6 ),
    .B2(\i44/n562 ),
    .Y(\i44/n229 ));
 OAI22xp33_ASAP7_75t_SL \i44/i312  (.A1(\i44/n68 ),
    .A2(\i44/n55 ),
    .B1(\i44/n92 ),
    .B2(\i44/n70 ),
    .Y(\i44/n228 ));
 AOI22xp5_ASAP7_75t_SL \i44/i313  (.A1(\i44/n100 ),
    .A2(\i44/n91 ),
    .B1(\i44/n90 ),
    .B2(\i44/n62 ),
    .Y(\i44/n261 ));
 OAI22xp33_ASAP7_75t_SL \i44/i314  (.A1(\i44/n20 ),
    .A2(\i44/n68 ),
    .B1(\i44/n85 ),
    .B2(\i44/n89 ),
    .Y(\i44/n227 ));
 OAI22xp5_ASAP7_75t_SL \i44/i315  (.A1(\i44/n97 ),
    .A2(\i44/n9 ),
    .B1(\i44/n18 ),
    .B2(\i44/n92 ),
    .Y(\i44/n226 ));
 OAI22xp5_ASAP7_75t_SL \i44/i316  (.A1(\i44/n70 ),
    .A2(\i44/n9 ),
    .B1(\i44/n89 ),
    .B2(\i44/n81 ),
    .Y(\i44/n225 ));
 AOI22xp5_ASAP7_75t_SL \i44/i317  (.A1(\i44/n54 ),
    .A2(\i44/n56 ),
    .B1(\i44/n100 ),
    .B2(\i44/n80 ),
    .Y(\i44/n260 ));
 OAI22xp33_ASAP7_75t_SL \i44/i318  (.A1(\i44/n538 ),
    .A2(\i44/n68 ),
    .B1(\i44/n17 ),
    .B2(\i44/n60 ),
    .Y(\i44/n224 ));
 AOI22xp5_ASAP7_75t_SL \i44/i319  (.A1(\i44/n71 ),
    .A2(\i44/n86 ),
    .B1(\i44/n56 ),
    .B2(\i44/n88 ),
    .Y(\i44/n223 ));
 NOR2x1_ASAP7_75t_SL \i44/i32  (.A(\i44/n502 ),
    .B(\i44/n462 ),
    .Y(\i44/n518 ));
 OAI22xp5_ASAP7_75t_SL \i44/i320  (.A1(\i44/n68 ),
    .A2(\i44/n96 ),
    .B1(\i44/n73 ),
    .B2(\i44/n17 ),
    .Y(\i44/n222 ));
 OAI21xp5_ASAP7_75t_SL \i44/i321  (.A1(\i44/n539 ),
    .A2(\i44/n63 ),
    .B(\i44/n138 ),
    .Y(\i44/n258 ));
 AOI22xp5_ASAP7_75t_SL \i44/i322  (.A1(\i44/n54 ),
    .A2(\i44/n72 ),
    .B1(\i44/n56 ),
    .B2(\i44/n62 ),
    .Y(\i44/n256 ));
 AOI22xp5_ASAP7_75t_SL \i44/i323  (.A1(\i44/n58 ),
    .A2(\i44/n59 ),
    .B1(\i44/n66 ),
    .B2(\i44/n71 ),
    .Y(\i44/n254 ));
 AOI22xp5_ASAP7_75t_SL \i44/i324  (.A1(\i44/n94 ),
    .A2(\i44/n100 ),
    .B1(\i44/n546 ),
    .B2(\i44/n79 ),
    .Y(\i44/n253 ));
 OAI22xp5_ASAP7_75t_SL \i44/i325  (.A1(\i44/n55 ),
    .A2(\i44/n18 ),
    .B1(\i44/n68 ),
    .B2(\i44/n78 ),
    .Y(\i44/n221 ));
 NAND2xp33_ASAP7_75t_SL \i44/i326  (.A(\i44/n218 ),
    .B(\i44/n219 ),
    .Y(\i44/n220 ));
 OAI22x1_ASAP7_75t_SL \i44/i327  (.A1(\i44/n19 ),
    .A2(\i44/n96 ),
    .B1(\i44/n57 ),
    .B2(\i44/n551 ),
    .Y(\i44/n251 ));
 AOI22xp5_ASAP7_75t_SL \i44/i328  (.A1(\i44/n58 ),
    .A2(\i44/n66 ),
    .B1(\i44/n56 ),
    .B2(\i44/n94 ),
    .Y(\i44/n249 ));
 AO22x2_ASAP7_75t_SL \i44/i329  (.A1(\i44/n98 ),
    .A2(\i44/n95 ),
    .B1(\i44/n61 ),
    .B2(\i44/n88 ),
    .Y(\i44/n248 ));
 NAND2xp5_ASAP7_75t_SL \i44/i33  (.A(\i44/n460 ),
    .B(\i44/n479 ),
    .Y(\i44/n517 ));
 OAI21xp5_ASAP7_75t_SL \i44/i330  (.A1(\i44/n83 ),
    .A2(\i44/n538 ),
    .B(\i44/n121 ),
    .Y(\i44/n247 ));
 OAI22xp5_ASAP7_75t_L \i44/i331  (.A1(\i44/n87 ),
    .A2(\i44/n55 ),
    .B1(\i44/n85 ),
    .B2(\i44/n539 ),
    .Y(\i44/n245 ));
 OAI22xp5_ASAP7_75t_SL \i44/i332  (.A1(\i44/n70 ),
    .A2(\i44/n538 ),
    .B1(\i44/n73 ),
    .B2(\i44/n85 ),
    .Y(\i44/n243 ));
 AOI22xp5_ASAP7_75t_SL \i44/i333  (.A1(\i44/n54 ),
    .A2(\i44/n58 ),
    .B1(\i44/n75 ),
    .B2(\i44/n88 ),
    .Y(\i44/n242 ));
 OAI22xp5_ASAP7_75t_SL \i44/i334  (.A1(\i44/n60 ),
    .A2(\i44/n67 ),
    .B1(\i44/n73 ),
    .B2(\i44/n551 ),
    .Y(\i44/n241 ));
 AOI22xp5_ASAP7_75t_SL \i44/i335  (.A1(\i44/n65 ),
    .A2(\i44/n88 ),
    .B1(\i44/n56 ),
    .B2(\i44/n66 ),
    .Y(\i44/n240 ));
 AOI22xp5_ASAP7_75t_SL \i44/i336  (.A1(\i44/n100 ),
    .A2(\i44/n59 ),
    .B1(\i44/n545 ),
    .B2(\i44/n79 ),
    .Y(\i44/n239 ));
 INVxp67_ASAP7_75t_SL \i44/i337  (.A(\i44/n213 ),
    .Y(\i44/n214 ));
 INVx1_ASAP7_75t_SL \i44/i338  (.A(\i44/n211 ),
    .Y(\i44/n212 ));
 INVxp67_ASAP7_75t_SL \i44/i339  (.A(\i44/n209 ),
    .Y(\i44/n210 ));
 NOR3x1_ASAP7_75t_SL \i44/i34  (.A(\i44/n30 ),
    .B(\i44/n475 ),
    .C(\i44/n402 ),
    .Y(\i44/n525 ));
 INVxp67_ASAP7_75t_SL \i44/i340  (.A(\i44/n207 ),
    .Y(\i44/n208 ));
 INVxp67_ASAP7_75t_SL \i44/i341  (.A(\i44/n205 ),
    .Y(\i44/n206 ));
 INVxp67_ASAP7_75t_SL \i44/i342  (.A(\i44/n568 ),
    .Y(\i44/n203 ));
 INVxp67_ASAP7_75t_SL \i44/i343  (.A(\i44/n197 ),
    .Y(\i44/n198 ));
 INVxp67_ASAP7_75t_SL \i44/i344  (.A(\i44/n195 ),
    .Y(\i44/n196 ));
 INVxp67_ASAP7_75t_SL \i44/i345  (.A(\i44/n192 ),
    .Y(\i44/n193 ));
 INVxp67_ASAP7_75t_SL \i44/i346  (.A(\i44/n190 ),
    .Y(\i44/n191 ));
 INVxp67_ASAP7_75t_SL \i44/i347  (.A(\i44/n188 ),
    .Y(\i44/n189 ));
 INVxp67_ASAP7_75t_SL \i44/i348  (.A(\i44/n186 ),
    .Y(\i44/n187 ));
 INVx1_ASAP7_75t_SL \i44/i349  (.A(\i44/n185 ),
    .Y(\i44/n184 ));
 NOR3xp33_ASAP7_75t_SL \i44/i35  (.A(\i44/n421 ),
    .B(\i44/n30 ),
    .C(\i44/n499 ),
    .Y(\i44/n515 ));
 NAND2xp5_ASAP7_75t_SL \i44/i350  (.A(\i44/n72 ),
    .B(\i44/n91 ),
    .Y(\i44/n219 ));
 NAND2xp5_ASAP7_75t_SL \i44/i351  (.A(\i44/n90 ),
    .B(\i44/n88 ),
    .Y(\i44/n183 ));
 NAND2xp5_ASAP7_75t_SL \i44/i352  (.A(\i44/n89 ),
    .B(\i44/n87 ),
    .Y(\i44/n182 ));
 NAND2xp5_ASAP7_75t_SL \i44/i353  (.A(\i44/n56 ),
    .B(\i44/n95 ),
    .Y(\i44/n181 ));
 NAND2xp33_ASAP7_75t_SL \i44/i354  (.A(\i44/n70 ),
    .B(\i44/n537 ),
    .Y(\i44/n180 ));
 NAND2xp5_ASAP7_75t_SL \i44/i355  (.A(\i44/n64 ),
    .B(\i44/n69 ),
    .Y(\i44/n179 ));
 NAND2xp5_ASAP7_75t_SL \i44/i356  (.A(\i44/n64 ),
    .B(\i44/n71 ),
    .Y(\i44/n218 ));
 NAND2xp5_ASAP7_75t_SL \i44/i357  (.A(\i44/n69 ),
    .B(\i44/n77 ),
    .Y(\i44/n217 ));
 NAND2xp5_ASAP7_75t_SL \i44/i358  (.A(\i44/n71 ),
    .B(\i44/n91 ),
    .Y(\i44/n178 ));
 NAND2xp5_ASAP7_75t_SL \i44/i359  (.A(\i44/n3 ),
    .B(\i44/n69 ),
    .Y(\i44/n177 ));
 NOR2xp67_ASAP7_75t_SL \i44/i36  (.A(\i44/n480 ),
    .B(\i44/n30 ),
    .Y(\i44/n514 ));
 NAND2xp5_ASAP7_75t_SL \i44/i360  (.A(\i44/n73 ),
    .B(\i44/n18 ),
    .Y(\i44/n176 ));
 NAND2xp5_ASAP7_75t_SL \i44/i361  (.A(\i44/n90 ),
    .B(\i44/n94 ),
    .Y(\i44/n175 ));
 NAND2xp5_ASAP7_75t_SL \i44/i362  (.A(\i44/n72 ),
    .B(\i44/n3 ),
    .Y(\i44/n174 ));
 NAND2xp5_ASAP7_75t_SL \i44/i363  (.A(\i44/n79 ),
    .B(\i44/n75 ),
    .Y(\i44/n173 ));
 NAND2xp5_ASAP7_75t_SL \i44/i364  (.A(\i44/n71 ),
    .B(\i44/n79 ),
    .Y(\i44/n172 ));
 NAND2xp5_ASAP7_75t_SL \i44/i365  (.A(\i44/n54 ),
    .B(\i44/n61 ),
    .Y(\i44/n171 ));
 NAND2xp5_ASAP7_75t_SL \i44/i366  (.A(\i44/n61 ),
    .B(\i44/n77 ),
    .Y(\i44/n170 ));
 NAND2xp5_ASAP7_75t_SL \i44/i367  (.A(\i44/n72 ),
    .B(\i44/n94 ),
    .Y(\i44/n169 ));
 NAND2xp5_ASAP7_75t_SL \i44/i368  (.A(\i44/n54 ),
    .B(\i44/n84 ),
    .Y(\i44/n216 ));
 AND2x2_ASAP7_75t_SL \i44/i369  (.A(\i44/n61 ),
    .B(\i44/n80 ),
    .Y(\i44/n215 ));
 NOR3xp33_ASAP7_75t_SL \i44/i37  (.A(\i44/n458 ),
    .B(\i44/n453 ),
    .C(\i44/n2 ),
    .Y(\i44/n513 ));
 AND2x2_ASAP7_75t_SL \i44/i370  (.A(\i44/n90 ),
    .B(\i44/n77 ),
    .Y(\i44/n213 ));
 AND2x2_ASAP7_75t_SL \i44/i371  (.A(\i44/n100 ),
    .B(\i44/n79 ),
    .Y(\i44/n211 ));
 NAND2xp5_ASAP7_75t_SL \i44/i372  (.A(\i44/n79 ),
    .B(\i44/n6 ),
    .Y(\i44/n26 ));
 NAND2xp5_ASAP7_75t_SL \i44/i373  (.A(\i44/n84 ),
    .B(\i44/n94 ),
    .Y(\i44/n209 ));
 NAND2xp5_ASAP7_75t_SL \i44/i374  (.A(\i44/n98 ),
    .B(\i44/n59 ),
    .Y(\i44/n207 ));
 NAND2xp5_ASAP7_75t_SL \i44/i375  (.A(\i44/n545 ),
    .B(\i44/n77 ),
    .Y(\i44/n205 ));
 AND2x2_ASAP7_75t_SL \i44/i376  (.A(\i44/n72 ),
    .B(\i44/n66 ),
    .Y(\i44/n204 ));
 NAND2xp5_ASAP7_75t_SL \i44/i377  (.A(\i44/n565 ),
    .B(\i44/n3 ),
    .Y(\i44/n168 ));
 NAND2xp5_ASAP7_75t_SL \i44/i378  (.A(\i44/n82 ),
    .B(\i44/n565 ),
    .Y(\i44/n202 ));
 NOR2xp33_ASAP7_75t_SL \i44/i379  (.A(\i44/n74 ),
    .B(\i44/n85 ),
    .Y(\i44/n167 ));
 NAND4xp25_ASAP7_75t_SL \i44/i38  (.A(\i44/n440 ),
    .B(\i44/n541 ),
    .C(\i44/n434 ),
    .D(\i44/n467 ),
    .Y(\i44/n512 ));
 NAND2xp5_ASAP7_75t_SL \i44/i380  (.A(\i44/n545 ),
    .B(\i44/n64 ),
    .Y(\i44/n201 ));
 NAND2xp5_ASAP7_75t_SL \i44/i381  (.A(\i44/n66 ),
    .B(\i44/n69 ),
    .Y(\i44/n166 ));
 NOR2xp33_ASAP7_75t_SL \i44/i382  (.A(\i44/n68 ),
    .B(\i44/n85 ),
    .Y(\i44/n200 ));
 AND2x2_ASAP7_75t_SL \i44/i383  (.A(\i44/n71 ),
    .B(\i44/n3 ),
    .Y(\i44/n199 ));
 NOR2xp33_ASAP7_75t_SL \i44/i384  (.A(\i44/n19 ),
    .B(\i44/n17 ),
    .Y(\i44/n165 ));
 NAND2xp5_ASAP7_75t_SL \i44/i385  (.A(\i44/n565 ),
    .B(\i44/n59 ),
    .Y(\i44/n197 ));
 NOR2xp33_ASAP7_75t_SL \i44/i386  (.A(\i44/n545 ),
    .B(\i44/n90 ),
    .Y(\i44/n164 ));
 NOR2xp33_ASAP7_75t_SL \i44/i387  (.A(\i44/n68 ),
    .B(\i44/n93 ),
    .Y(\i44/n163 ));
 NAND2xp5_ASAP7_75t_SL \i44/i388  (.A(\i44/n90 ),
    .B(\i44/n3 ),
    .Y(\i44/n195 ));
 NOR2xp33_ASAP7_75t_L \i44/i389  (.A(\i44/n98 ),
    .B(\i44/n58 ),
    .Y(\i44/n194 ));
 NAND3xp33_ASAP7_75t_L \i44/i39  (.A(\i44/n419 ),
    .B(\i44/n541 ),
    .C(\i44/n484 ),
    .Y(\i44/n511 ));
 NAND2xp5_ASAP7_75t_SL \i44/i390  (.A(\i44/n545 ),
    .B(\i44/n86 ),
    .Y(\i44/n25 ));
 NAND2xp5_ASAP7_75t_SL \i44/i391  (.A(\i44/n98 ),
    .B(\i44/n62 ),
    .Y(\i44/n192 ));
 NAND2xp5_ASAP7_75t_SL \i44/i392  (.A(\i44/n94 ),
    .B(\i44/n71 ),
    .Y(\i44/n190 ));
 NAND2xp5_ASAP7_75t_SL \i44/i393  (.A(\i44/n98 ),
    .B(\i44/n79 ),
    .Y(\i44/n188 ));
 NAND2xp5_ASAP7_75t_SL \i44/i394  (.A(\i44/n72 ),
    .B(\i44/n82 ),
    .Y(\i44/n162 ));
 NOR2xp33_ASAP7_75t_SL \i44/i395  (.A(\i44/n90 ),
    .B(\i44/n72 ),
    .Y(\i44/n186 ));
 NOR2x1_ASAP7_75t_SL \i44/i396  (.A(\i44/n89 ),
    .B(\i44/n63 ),
    .Y(\i44/n161 ));
 OR2x2_ASAP7_75t_SL \i44/i397  (.A(\i44/n58 ),
    .B(\i44/n565 ),
    .Y(\i44/n185 ));
 INVxp67_ASAP7_75t_SL \i44/i398  (.A(\i44/n159 ),
    .Y(\i44/n160 ));
 INVxp67_ASAP7_75t_SL \i44/i399  (.A(\i44/n154 ),
    .Y(\i44/n155 ));
 INVx2_ASAP7_75t_SL \i44/i4  (.A(\i44/n552 ),
    .Y(\i44/n4 ));
 NAND3xp33_ASAP7_75t_SL \i44/i40  (.A(\i44/n543 ),
    .B(\i44/n468 ),
    .C(\i44/n454 ),
    .Y(\i44/n510 ));
 INVx1_ASAP7_75t_SL \i44/i400  (.A(\i44/n152 ),
    .Y(\i44/n153 ));
 INVxp67_ASAP7_75t_SL \i44/i401  (.A(\i44/n146 ),
    .Y(\i44/n147 ));
 INVxp67_ASAP7_75t_SL \i44/i402  (.A(\i44/n144 ),
    .Y(\i44/n145 ));
 INVxp67_ASAP7_75t_SL \i44/i403  (.A(\i44/n142 ),
    .Y(\i44/n143 ));
 INVxp67_ASAP7_75t_SL \i44/i404  (.A(\i44/n140 ),
    .Y(\i44/n141 ));
 INVxp67_ASAP7_75t_SL \i44/i405  (.A(\i44/n540 ),
    .Y(\i44/n139 ));
 INVxp67_ASAP7_75t_SL \i44/i406  (.A(\i44/n137 ),
    .Y(\i44/n138 ));
 INVxp67_ASAP7_75t_SL \i44/i407  (.A(\i44/n129 ),
    .Y(\i44/n130 ));
 INVx1_ASAP7_75t_SL \i44/i408  (.A(\i44/n125 ),
    .Y(\i44/n126 ));
 INVx2_ASAP7_75t_SL \i44/i409  (.A(\i44/n21 ),
    .Y(\i44/n22 ));
 NAND2xp5_ASAP7_75t_L \i44/i41  (.A(\i44/n575 ),
    .B(\i44/n500 ),
    .Y(\i44/n509 ));
 NAND2xp5_ASAP7_75t_SL \i44/i410  (.A(\i44/n546 ),
    .B(\i44/n80 ),
    .Y(\i44/n124 ));
 NAND2xp5_ASAP7_75t_SL \i44/i411  (.A(\i44/n58 ),
    .B(\i44/n82 ),
    .Y(\i44/n123 ));
 NAND2xp5_ASAP7_75t_SL \i44/i412  (.A(\i44/n65 ),
    .B(\i44/n80 ),
    .Y(\i44/n24 ));
 NAND2xp5_ASAP7_75t_SL \i44/i413  (.A(\i44/n83 ),
    .B(\i44/n74 ),
    .Y(\i44/n122 ));
 NAND2xp5_ASAP7_75t_SL \i44/i414  (.A(\i44/n65 ),
    .B(\i44/n82 ),
    .Y(\i44/n121 ));
 NAND2xp5_ASAP7_75t_SL \i44/i415  (.A(\i44/n82 ),
    .B(\i44/n56 ),
    .Y(\i44/n120 ));
 NAND2xp5_ASAP7_75t_SL \i44/i416  (.A(\i44/n84 ),
    .B(\i44/n66 ),
    .Y(\i44/n119 ));
 NOR2xp33_ASAP7_75t_SL \i44/i417  (.A(\i44/n94 ),
    .B(\i44/n3 ),
    .Y(\i44/n118 ));
 NAND2xp5_ASAP7_75t_R \i44/i418  (.A(\i44/n75 ),
    .B(\i44/n62 ),
    .Y(\i44/n117 ));
 NAND2xp5_ASAP7_75t_SL \i44/i419  (.A(\i44/n56 ),
    .B(\i44/n77 ),
    .Y(\i44/n116 ));
 NAND2xp33_ASAP7_75t_SL \i44/i42  (.A(\i44/n465 ),
    .B(\i44/n482 ),
    .Y(\i44/n508 ));
 NAND2xp5_ASAP7_75t_L \i44/i420  (.A(\i44/n20 ),
    .B(\i44/n55 ),
    .Y(\i44/n115 ));
 NAND2xp33_ASAP7_75t_SL \i44/i421  (.A(\i44/n67 ),
    .B(\i44/n9 ),
    .Y(\i44/n114 ));
 NAND2xp5_ASAP7_75t_SL \i44/i422  (.A(\i44/n6 ),
    .B(\i44/n64 ),
    .Y(\i44/n113 ));
 NAND2xp5_ASAP7_75t_SL \i44/i423  (.A(\i44/n100 ),
    .B(\i44/n562 ),
    .Y(\i44/n159 ));
 NAND2xp5_ASAP7_75t_SL \i44/i424  (.A(\i44/n546 ),
    .B(\i44/n64 ),
    .Y(\i44/n112 ));
 NOR2xp33_ASAP7_75t_SL \i44/i425  (.A(\i44/n63 ),
    .B(\i44/n537 ),
    .Y(\i44/n111 ));
 NAND2xp5_ASAP7_75t_SL \i44/i426  (.A(\i44/n100 ),
    .B(\i44/n3 ),
    .Y(\i44/n158 ));
 AND2x2_ASAP7_75t_SL \i44/i427  (.A(\i44/n6 ),
    .B(\i44/n82 ),
    .Y(\i44/n157 ));
 NOR2xp33_ASAP7_75t_SL \i44/i428  (.A(\i44/n94 ),
    .B(\i44/n86 ),
    .Y(\i44/n156 ));
 NAND2xp5_ASAP7_75t_SL \i44/i429  (.A(\i44/n90 ),
    .B(\i44/n66 ),
    .Y(\i44/n154 ));
 NOR2x1_ASAP7_75t_SL \i44/i43  (.A(\i44/n490 ),
    .B(\i44/n481 ),
    .Y(\i44/n516 ));
 NOR2x1_ASAP7_75t_SL \i44/i430  (.A(\i44/n77 ),
    .B(\i44/n88 ),
    .Y(\i44/n152 ));
 NAND2xp5_ASAP7_75t_SL \i44/i431  (.A(\i44/n6 ),
    .B(\i44/n86 ),
    .Y(\i44/n151 ));
 NAND2xp5_ASAP7_75t_SL \i44/i432  (.A(\i44/n84 ),
    .B(\i44/n62 ),
    .Y(\i44/n150 ));
 NAND2xp5_ASAP7_75t_SL \i44/i433  (.A(\i44/n56 ),
    .B(\i44/n80 ),
    .Y(\i44/n110 ));
 NAND2xp5_ASAP7_75t_SL \i44/i434  (.A(\i44/n61 ),
    .B(\i44/n64 ),
    .Y(\i44/n149 ));
 AND2x2_ASAP7_75t_SL \i44/i435  (.A(\i44/n6 ),
    .B(\i44/n59 ),
    .Y(\i44/n148 ));
 NOR2xp33_ASAP7_75t_SL \i44/i436  (.A(\i44/n77 ),
    .B(\i44/n64 ),
    .Y(\i44/n109 ));
 NAND2xp5_ASAP7_75t_SL \i44/i437  (.A(\i44/n546 ),
    .B(\i44/n94 ),
    .Y(\i44/n146 ));
 NAND2xp5_ASAP7_75t_SL \i44/i438  (.A(\i44/n546 ),
    .B(\i44/n59 ),
    .Y(\i44/n144 ));
 NOR2xp67_ASAP7_75t_SL \i44/i439  (.A(\i44/n60 ),
    .B(\i44/n92 ),
    .Y(\i44/n142 ));
 NAND2xp33_ASAP7_75t_L \i44/i44  (.A(\i44/n470 ),
    .B(\i44/n442 ),
    .Y(\i44/n505 ));
 NAND2xp5_ASAP7_75t_SL \i44/i440  (.A(\i44/n56 ),
    .B(\i44/n59 ),
    .Y(\i44/n140 ));
 NAND2xp33_ASAP7_75t_L \i44/i441  (.A(\i44/n538 ),
    .B(\i44/n551 ),
    .Y(\i44/n108 ));
 NOR2xp67_ASAP7_75t_L \i44/i442  (.A(\i44/n55 ),
    .B(\i44/n537 ),
    .Y(\i44/n137 ));
 NAND2xp5_ASAP7_75t_SL \i44/i443  (.A(\i44/n58 ),
    .B(\i44/n86 ),
    .Y(\i44/n23 ));
 NAND2xp5_ASAP7_75t_SL \i44/i444  (.A(\i44/n58 ),
    .B(\i44/n88 ),
    .Y(\i44/n136 ));
 AND2x2_ASAP7_75t_SL \i44/i445  (.A(\i44/n100 ),
    .B(\i44/n88 ),
    .Y(\i44/n135 ));
 NAND2xp5_ASAP7_75t_SL \i44/i446  (.A(\i44/n3 ),
    .B(\i44/n65 ),
    .Y(\i44/n134 ));
 NAND2xp5_ASAP7_75t_SL \i44/i447  (.A(\i44/n17 ),
    .B(\i44/n20 ),
    .Y(\i44/n133 ));
 NAND2xp33_ASAP7_75t_L \i44/i448  (.A(\i44/n3 ),
    .B(\i44/n84 ),
    .Y(\i44/n107 ));
 AND2x2_ASAP7_75t_SL \i44/i449  (.A(\i44/n100 ),
    .B(\i44/n66 ),
    .Y(\i44/n132 ));
 NAND2xp33_ASAP7_75t_L \i44/i45  (.A(\i44/n575 ),
    .B(\i44/n448 ),
    .Y(\i44/n504 ));
 NOR2xp33_ASAP7_75t_SL \i44/i450  (.A(\i44/n67 ),
    .B(\i44/n539 ),
    .Y(\i44/n106 ));
 NOR2xp67_ASAP7_75t_SL \i44/i451  (.A(\i44/n562 ),
    .B(\i44/n80 ),
    .Y(\i44/n131 ));
 NAND2xp5_ASAP7_75t_SL \i44/i452  (.A(\i44/n6 ),
    .B(\i44/n88 ),
    .Y(\i44/n105 ));
 NAND2xp5_ASAP7_75t_SL \i44/i453  (.A(\i44/n65 ),
    .B(\i44/n62 ),
    .Y(\i44/n129 ));
 NAND2xp5_ASAP7_75t_SL \i44/i454  (.A(\i44/n56 ),
    .B(\i44/n3 ),
    .Y(\i44/n104 ));
 NAND2xp5_ASAP7_75t_SL \i44/i455  (.A(\i44/n84 ),
    .B(\i44/n88 ),
    .Y(\i44/n128 ));
 NAND2xp5_ASAP7_75t_SL \i44/i456  (.A(\i44/n65 ),
    .B(\i44/n86 ),
    .Y(\i44/n103 ));
 NAND2xp5_ASAP7_75t_SL \i44/i457  (.A(\i44/n100 ),
    .B(\i44/n82 ),
    .Y(\i44/n127 ));
 NOR2xp33_ASAP7_75t_SL \i44/i458  (.A(\i44/n99 ),
    .B(\i44/n17 ),
    .Y(\i44/n102 ));
 NOR2xp33_ASAP7_75t_SL \i44/i459  (.A(\i44/n99 ),
    .B(\i44/n63 ),
    .Y(\i44/n101 ));
 NOR2xp33_ASAP7_75t_SL \i44/i46  (.A(\i44/n447 ),
    .B(\i44/n472 ),
    .Y(\i44/n503 ));
 NAND2xp5_ASAP7_75t_SL \i44/i460  (.A(\i44/n65 ),
    .B(\i44/n91 ),
    .Y(\i44/n125 ));
 NAND2x1_ASAP7_75t_SL \i44/i461  (.A(\i44/n6 ),
    .B(\i44/n62 ),
    .Y(\i44/n21 ));
 INVx2_ASAP7_75t_SL \i44/i462  (.A(\i44/n100 ),
    .Y(\i44/n99 ));
 INVx1_ASAP7_75t_SL \i44/i463  (.A(\i44/n98 ),
    .Y(\i44/n97 ));
 INVx3_ASAP7_75t_SL \i44/i464  (.A(\i44/n96 ),
    .Y(\i44/n95 ));
 INVx2_ASAP7_75t_SL \i44/i465  (.A(\i44/n94 ),
    .Y(\i44/n93 ));
 INVx4_ASAP7_75t_SL \i44/i466  (.A(\i44/n92 ),
    .Y(\i44/n91 ));
 INVx3_ASAP7_75t_SL \i44/i467  (.A(\i44/n90 ),
    .Y(\i44/n89 ));
 INVx2_ASAP7_75t_SL \i44/i468  (.A(\i44/n546 ),
    .Y(\i44/n87 ));
 INVx4_ASAP7_75t_SL \i44/i469  (.A(\i44/n86 ),
    .Y(\i44/n85 ));
 NAND3xp33_ASAP7_75t_SL \i44/i47  (.A(\i44/n437 ),
    .B(\i44/n445 ),
    .C(\i44/n414 ),
    .Y(\i44/n502 ));
 INVx2_ASAP7_75t_SL \i44/i470  (.A(\i44/n84 ),
    .Y(\i44/n83 ));
 INVx3_ASAP7_75t_SL \i44/i471  (.A(\i44/n82 ),
    .Y(\i44/n81 ));
 INVx2_ASAP7_75t_SL \i44/i472  (.A(\i44/n79 ),
    .Y(\i44/n78 ));
 INVx4_ASAP7_75t_SL \i44/i473  (.A(\i44/n77 ),
    .Y(\i44/n76 ));
 INVx2_ASAP7_75t_SL \i44/i474  (.A(\i44/n75 ),
    .Y(\i44/n74 ));
 INVx3_ASAP7_75t_SL \i44/i475  (.A(\i44/n73 ),
    .Y(\i44/n72 ));
 AND2x4_ASAP7_75t_SL \i44/i476  (.A(\i44/n44 ),
    .B(\i44/n49 ),
    .Y(\i44/n100 ));
 AND2x4_ASAP7_75t_SL \i44/i477  (.A(\i44/n47 ),
    .B(\i44/n44 ),
    .Y(\i44/n98 ));
 OR2x4_ASAP7_75t_SL \i44/i478  (.A(\i44/n36 ),
    .B(\i44/n7 ),
    .Y(\i44/n96 ));
 AND2x4_ASAP7_75t_SL \i44/i479  (.A(\i44/n41 ),
    .B(\i44/n4 ),
    .Y(\i44/n94 ));
 NOR2x1_ASAP7_75t_SL \i44/i48  (.A(\i44/n395 ),
    .B(\i44/n456 ),
    .Y(\i44/n501 ));
 OR2x6_ASAP7_75t_SL \i44/i480  (.A(\i44/n39 ),
    .B(\i44/n53 ),
    .Y(\i44/n92 ));
 AND2x4_ASAP7_75t_SL \i44/i481  (.A(\i44/n35 ),
    .B(\i44/n51 ),
    .Y(\i44/n90 ));
 AND2x4_ASAP7_75t_SL \i44/i482  (.A(\i44/n38 ),
    .B(\i44/n42 ),
    .Y(\i44/n88 ));
 NAND2x1p5_ASAP7_75t_SL \i44/i483  (.A(\i44/n38 ),
    .B(\i44/n42 ),
    .Y(\i44/n20 ));
 AND2x4_ASAP7_75t_SL \i44/i484  (.A(\i44/n52 ),
    .B(\i44/n37 ),
    .Y(\i44/n86 ));
 AND2x4_ASAP7_75t_SL \i44/i485  (.A(\i44/n35 ),
    .B(\i44/n46 ),
    .Y(\i44/n84 ));
 AND2x4_ASAP7_75t_SL \i44/i486  (.A(\i44/n38 ),
    .B(\i44/n40 ),
    .Y(\i44/n82 ));
 AND2x4_ASAP7_75t_SL \i44/i487  (.A(\i44/n41 ),
    .B(\i44/n5 ),
    .Y(\i44/n80 ));
 AND2x4_ASAP7_75t_SL \i44/i488  (.A(\i44/n41 ),
    .B(\i44/n38 ),
    .Y(\i44/n79 ));
 AND2x4_ASAP7_75t_SL \i44/i489  (.A(\i44/n38 ),
    .B(\i44/n37 ),
    .Y(\i44/n77 ));
 NOR2xp33_ASAP7_75t_SL \i44/i49  (.A(\i44/n463 ),
    .B(\i44/n375 ),
    .Y(\i44/n500 ));
 AND2x4_ASAP7_75t_SL \i44/i490  (.A(\i44/n47 ),
    .B(\i44/n45 ),
    .Y(\i44/n75 ));
 OR2x6_ASAP7_75t_SL \i44/i491  (.A(\i44/n48 ),
    .B(\i44/n34 ),
    .Y(\i44/n73 ));
 INVx2_ASAP7_75t_SL \i44/i492  (.A(\i44/n71 ),
    .Y(\i44/n19 ));
 INVx3_ASAP7_75t_SL \i44/i493  (.A(\i44/n545 ),
    .Y(\i44/n70 ));
 INVx3_ASAP7_75t_SL \i44/i494  (.A(\i44/n69 ),
    .Y(\i44/n68 ));
 INVx4_ASAP7_75t_SL \i44/i495  (.A(\i44/n67 ),
    .Y(\i44/n66 ));
 INVx4_ASAP7_75t_SL \i44/i496  (.A(\i44/n64 ),
    .Y(\i44/n63 ));
 INVx3_ASAP7_75t_SL \i44/i497  (.A(\i44/n62 ),
    .Y(\i44/n17 ));
 INVx4_ASAP7_75t_SL \i44/i498  (.A(\i44/n61 ),
    .Y(\i44/n60 ));
 INVx3_ASAP7_75t_SL \i44/i499  (.A(\i44/n58 ),
    .Y(\i44/n57 ));
 INVx1_ASAP7_75t_SL \i44/i5  (.A(\i44/n36 ),
    .Y(\i44/n5 ));
 NAND2xp5_ASAP7_75t_SL \i44/i50  (.A(\i44/n470 ),
    .B(\i44/n466 ),
    .Y(\i44/n499 ));
 INVx13_ASAP7_75t_SL \i44/i500  (.A(\i44/n55 ),
    .Y(\i44/n54 ));
 AND2x4_ASAP7_75t_SL \i44/i501  (.A(\i44/n44 ),
    .B(\i44/n51 ),
    .Y(\i44/n71 ));
 OR2x2_ASAP7_75t_SL \i44/i502  (.A(\i44/n10 ),
    .B(\i44/n50 ),
    .Y(\i44/n18 ));
 AND2x4_ASAP7_75t_SL \i44/i503  (.A(\i44/n46 ),
    .B(\i44/n44 ),
    .Y(\i44/n69 ));
 NAND2x1p5_ASAP7_75t_SL \i44/i504  (.A(\i44/n41 ),
    .B(\i44/n52 ),
    .Y(\i44/n67 ));
 NAND2x1p5_ASAP7_75t_SL \i44/i505  (.A(\i44/n4 ),
    .B(\i44/n40 ),
    .Y(\i44/n9 ));
 AND2x4_ASAP7_75t_SL \i44/i506  (.A(\i44/n46 ),
    .B(\i44/n11 ),
    .Y(\i44/n65 ));
 AND2x4_ASAP7_75t_SL \i44/i507  (.A(\i44/n40 ),
    .B(\i44/n5 ),
    .Y(\i44/n64 ));
 AND2x4_ASAP7_75t_SL \i44/i508  (.A(\i44/n37 ),
    .B(\i44/n5 ),
    .Y(\i44/n62 ));
 AND2x4_ASAP7_75t_SL \i44/i509  (.A(\i44/n49 ),
    .B(\i44/n11 ),
    .Y(\i44/n61 ));
 NOR2x1_ASAP7_75t_SL \i44/i51  (.A(\i44/n379 ),
    .B(\i44/n472 ),
    .Y(\i44/n498 ));
 AND2x4_ASAP7_75t_SL \i44/i510  (.A(\i44/n4 ),
    .B(\i44/n42 ),
    .Y(\i44/n59 ));
 AND2x4_ASAP7_75t_SL \i44/i511  (.A(\i44/n46 ),
    .B(\i44/n45 ),
    .Y(\i44/n58 ));
 AND2x4_ASAP7_75t_SL \i44/i512  (.A(\i44/n51 ),
    .B(\i44/n45 ),
    .Y(\i44/n56 ));
 OR2x6_ASAP7_75t_SL \i44/i513  (.A(\i44/n33 ),
    .B(\i44/n43 ),
    .Y(\i44/n55 ));
 INVx2_ASAP7_75t_SL \i44/i514  (.A(\i44/n52 ),
    .Y(\i44/n53 ));
 INVx2_ASAP7_75t_SL \i44/i515  (.A(\i44/n50 ),
    .Y(\i44/n51 ));
 INVx3_ASAP7_75t_SL \i44/i516  (.A(\i44/n48 ),
    .Y(\i44/n49 ));
 NAND2xp5_ASAP7_75t_SL \i44/i517  (.A(\i44/n12 ),
    .B(\i44/n1 ),
    .Y(\i44/n43 ));
 AND2x2_ASAP7_75t_SL \i44/i518  (.A(\i44/n12 ),
    .B(\i44/n1 ),
    .Y(\i44/n52 ));
 NAND2xp5_ASAP7_75t_SL \i44/i519  (.A(\i44/n0 ),
    .B(n33[5]),
    .Y(\i44/n50 ));
 NOR2x1_ASAP7_75t_SL \i44/i52  (.A(\i44/n446 ),
    .B(\i44/n457 ),
    .Y(\i44/n497 ));
 NAND2x1p5_ASAP7_75t_SL \i44/i520  (.A(n33[4]),
    .B(n33[5]),
    .Y(\i44/n48 ));
 AND2x4_ASAP7_75t_SL \i44/i521  (.A(\i44/n31 ),
    .B(\i44/n0 ),
    .Y(\i44/n47 ));
 AND2x2_ASAP7_75t_SL \i44/i522  (.A(n33[4]),
    .B(\i44/n31 ),
    .Y(\i44/n46 ));
 AND2x2_ASAP7_75t_SL \i44/i523  (.A(n33[7]),
    .B(\i44/n16 ),
    .Y(\i44/n45 ));
 AND2x2_ASAP7_75t_SL \i44/i524  (.A(\i44/n14 ),
    .B(\i44/n16 ),
    .Y(\i44/n44 ));
 INVx2_ASAP7_75t_SL \i44/i525  (.A(\i44/n7 ),
    .Y(\i44/n42 ));
 INVx1_ASAP7_75t_SL \i44/i526  (.A(\i44/n40 ),
    .Y(\i44/n39 ));
 INVx2_ASAP7_75t_SL \i44/i527  (.A(\i44/n553 ),
    .Y(\i44/n37 ));
 INVx2_ASAP7_75t_SL \i44/i528  (.A(\i44/n35 ),
    .Y(\i44/n34 ));
 NAND2xp5_ASAP7_75t_SL \i44/i529  (.A(\i44/n32 ),
    .B(\i44/n13 ),
    .Y(\i44/n33 ));
 NAND2xp5_ASAP7_75t_SL \i44/i53  (.A(\i44/n413 ),
    .B(\i44/n451 ),
    .Y(\i44/n496 ));
 AND2x2_ASAP7_75t_SL \i44/i530  (.A(n33[0]),
    .B(n33[1]),
    .Y(\i44/n41 ));
 AND2x4_ASAP7_75t_SL \i44/i531  (.A(n33[0]),
    .B(\i44/n32 ),
    .Y(\i44/n40 ));
 AND2x4_ASAP7_75t_SL \i44/i532  (.A(n33[2]),
    .B(n33[3]),
    .Y(\i44/n38 ));
 NAND2x1_ASAP7_75t_SL \i44/i533  (.A(n33[3]),
    .B(\i44/n1 ),
    .Y(\i44/n36 ));
 AND2x2_ASAP7_75t_SL \i44/i534  (.A(n33[7]),
    .B(n33[6]),
    .Y(\i44/n35 ));
 INVx1_ASAP7_75t_SL \i44/i535  (.A(n33[1]),
    .Y(\i44/n32 ));
 INVx3_ASAP7_75t_SL \i44/i536  (.A(n33[5]),
    .Y(\i44/n31 ));
 INVx2_ASAP7_75t_SL \i44/i537  (.A(n33[6]),
    .Y(\i44/n16 ));
 INVx2_ASAP7_75t_SL \i44/i538  (.A(n33[7]),
    .Y(\i44/n14 ));
 INVx2_ASAP7_75t_SL \i44/i539  (.A(n33[0]),
    .Y(\i44/n13 ));
 NOR5xp2_ASAP7_75t_SL \i44/i54  (.A(\i44/n333 ),
    .B(\i44/n567 ),
    .C(\i44/n346 ),
    .D(\i44/n29 ),
    .E(\i44/n309 ),
    .Y(\i44/n495 ));
 INVx2_ASAP7_75t_SL \i44/i540  (.A(n33[3]),
    .Y(\i44/n12 ));
 AND2x2_ASAP7_75t_L \i44/i541  (.A(\i44/n14 ),
    .B(n33[6]),
    .Y(\i44/n11 ));
 NAND2xp5_ASAP7_75t_SL \i44/i542  (.A(\i44/n14 ),
    .B(n33[6]),
    .Y(\i44/n10 ));
 OR2x2_ASAP7_75t_SL \i44/i543  (.A(\i44/n148 ),
    .B(\i44/n557 ),
    .Y(\i44/n8 ));
 OR2x2_ASAP7_75t_SL \i44/i544  (.A(n33[0]),
    .B(n33[1]),
    .Y(\i44/n7 ));
 INVx4_ASAP7_75t_SL \i44/i545  (.A(\i44/n65 ),
    .Y(\i44/n537 ));
 NAND2x1p5_ASAP7_75t_L \i44/i546  (.A(\i44/n4 ),
    .B(\i44/n42 ),
    .Y(\i44/n538 ));
 INVx3_ASAP7_75t_SL \i44/i547  (.A(\i44/n56 ),
    .Y(\i44/n539 ));
 NAND2xp5_ASAP7_75t_SL \i44/i548  (.A(\i44/n54 ),
    .B(\i44/n100 ),
    .Y(\i44/n540 ));
 NOR2x1_ASAP7_75t_SL \i44/i549  (.A(\i44/n572 ),
    .B(\i44/n563 ),
    .Y(\i44/n541 ));
 NOR2x1_ASAP7_75t_SL \i44/i55  (.A(\i44/n2 ),
    .B(\i44/n458 ),
    .Y(\i44/n494 ));
 NOR2xp33_ASAP7_75t_SL \i44/i550  (.A(\i44/n563 ),
    .B(\i44/n373 ),
    .Y(\i44/n542 ));
 NOR2xp33_ASAP7_75t_SL \i44/i551  (.A(\i44/n564 ),
    .B(\i44/n333 ),
    .Y(\i44/n543 ));
 OA21x2_ASAP7_75t_SL \i44/i552  (.A1(\i44/n60 ),
    .A2(\i44/n554 ),
    .B(\i44/n24 ),
    .Y(\i44/n544 ));
 AND2x4_ASAP7_75t_SL \i44/i553  (.A(\i44/n49 ),
    .B(\i44/n45 ),
    .Y(\i44/n545 ));
 AND2x4_ASAP7_75t_SL \i44/i554  (.A(\i44/n35 ),
    .B(\i44/n47 ),
    .Y(\i44/n546 ));
 NOR2x1_ASAP7_75t_SL \i44/i555  (.A(\i44/n17 ),
    .B(\i44/n547 ),
    .Y(\i44/n548 ));
 NOR2x1_ASAP7_75t_SL \i44/i556  (.A(\i44/n545 ),
    .B(\i44/n546 ),
    .Y(\i44/n547 ));
 INVxp67_ASAP7_75t_SL \i44/i557  (.A(\i44/n547 ),
    .Y(\i44/n549 ));
 OAI221xp5_ASAP7_75t_SL \i44/i558  (.A1(\i44/n547 ),
    .A2(\i44/n96 ),
    .B1(\i44/n67 ),
    .B2(\i44/n74 ),
    .C(\i44/n190 ),
    .Y(\i44/n550 ));
 INVx2_ASAP7_75t_SL \i44/i559  (.A(\i44/n80 ),
    .Y(\i44/n551 ));
 NAND2x1_ASAP7_75t_SL \i44/i56  (.A(\i44/n455 ),
    .B(\i44/n435 ),
    .Y(\i44/n507 ));
 OR2x2_ASAP7_75t_SL \i44/i560  (.A(\i44/n1 ),
    .B(n33[3]),
    .Y(\i44/n552 ));
 NAND2xp5_ASAP7_75t_SL \i44/i561  (.A(\i44/n13 ),
    .B(n33[1]),
    .Y(\i44/n553 ));
 NOR2xp33_ASAP7_75t_SL \i44/i562  (.A(\i44/n554 ),
    .B(\i44/n57 ),
    .Y(\i44/n555 ));
 OR2x2_ASAP7_75t_SL \i44/i563  (.A(\i44/n552 ),
    .B(\i44/n553 ),
    .Y(\i44/n554 ));
 OAI22xp5_ASAP7_75t_SL \i44/i564  (.A1(\i44/n60 ),
    .A2(\i44/n538 ),
    .B1(\i44/n554 ),
    .B2(\i44/n57 ),
    .Y(\i44/n556 ));
 OAI22xp5_ASAP7_75t_SL \i44/i565  (.A1(\i44/n60 ),
    .A2(\i44/n85 ),
    .B1(\i44/n73 ),
    .B2(\i44/n554 ),
    .Y(\i44/n557 ));
 OAI21xp5_ASAP7_75t_SL \i44/i566  (.A1(\i44/n83 ),
    .A2(\i44/n554 ),
    .B(\i44/n149 ),
    .Y(\i44/n558 ));
 OAI22xp33_ASAP7_75t_SL \i44/i567  (.A1(\i44/n57 ),
    .A2(\i44/n96 ),
    .B1(\i44/n554 ),
    .B2(\i44/n68 ),
    .Y(\i44/n559 ));
 AOI31xp33_ASAP7_75t_SL \i44/i568  (.A1(\i44/n60 ),
    .A2(\i44/n87 ),
    .A3(\i44/n74 ),
    .B(\i44/n554 ),
    .Y(\i44/n560 ));
 AO21x1_ASAP7_75t_SL \i44/i569  (.A1(\i44/n554 ),
    .A2(\i44/n183 ),
    .B(\i44/n164 ),
    .Y(\i44/n561 ));
 NOR2x1_ASAP7_75t_SL \i44/i57  (.A(\i44/n473 ),
    .B(\i44/n457 ),
    .Y(\i44/n493 ));
 INVx4_ASAP7_75t_SL \i44/i570  (.A(\i44/n554 ),
    .Y(\i44/n562 ));
 OAI221xp5_ASAP7_75t_SL \i44/i571  (.A1(\i44/n537 ),
    .A2(\i44/n538 ),
    .B1(\i44/n554 ),
    .B2(\i44/n539 ),
    .C(\i44/n540 ),
    .Y(\i44/n563 ));
 OAI221xp5_ASAP7_75t_L \i44/i572  (.A1(\i44/n537 ),
    .A2(\i44/n538 ),
    .B1(\i44/n554 ),
    .B2(\i44/n539 ),
    .C(\i44/n540 ),
    .Y(\i44/n564 ));
 AND2x4_ASAP7_75t_SL \i44/i573  (.A(\i44/n47 ),
    .B(\i44/n11 ),
    .Y(\i44/n565 ));
 OAI221xp5_ASAP7_75t_SL \i44/i574  (.A1(\i44/n63 ),
    .A2(\i44/n566 ),
    .B1(\i44/n60 ),
    .B2(\i44/n554 ),
    .C(\i44/n24 ),
    .Y(\i44/n567 ));
 INVx4_ASAP7_75t_SL \i44/i575  (.A(\i44/n565 ),
    .Y(\i44/n566 ));
 NOR2xp67_ASAP7_75t_R \i44/i576  (.A(\i44/n554 ),
    .B(\i44/n566 ),
    .Y(\i44/n568 ));
 OA21x2_ASAP7_75t_SL \i44/i577  (.A1(\i44/n566 ),
    .A2(\i44/n17 ),
    .B(\i44/n201 ),
    .Y(\i44/n569 ));
 AOI21xp33_ASAP7_75t_SL \i44/i578  (.A1(\i44/n73 ),
    .A2(\i44/n566 ),
    .B(\i44/n55 ),
    .Y(\i44/n570 ));
 OAI22x1_ASAP7_75t_SL \i44/i579  (.A1(\i44/n81 ),
    .A2(\i44/n68 ),
    .B1(\i44/n78 ),
    .B2(\i44/n566 ),
    .Y(\i44/n571 ));
 NOR2x1_ASAP7_75t_SL \i44/i58  (.A(\i44/n394 ),
    .B(\i44/n456 ),
    .Y(\i44/n506 ));
 OAI22x1_ASAP7_75t_SL \i44/i580  (.A1(\i44/n566 ),
    .A2(\i44/n85 ),
    .B1(\i44/n74 ),
    .B2(\i44/n92 ),
    .Y(\i44/n572 ));
 NOR2xp67_ASAP7_75t_SL \i44/i581  (.A(\i44/n566 ),
    .B(\i44/n76 ),
    .Y(\i44/n573 ));
 AND4x1_ASAP7_75t_SL \i44/i582  (.A(\i44/n332 ),
    .B(\i44/n377 ),
    .C(\i44/n576 ),
    .D(\i44/n569 ),
    .Y(\i44/n574 ));
 AND4x1_ASAP7_75t_SL \i44/i583  (.A(\i44/n321 ),
    .B(\i44/n380 ),
    .C(\i44/n345 ),
    .D(\i44/n332 ),
    .Y(\i44/n575 ));
 AOI21xp5_ASAP7_75t_SL \i44/i584  (.A1(\i44/n61 ),
    .A2(\i44/n79 ),
    .B(\i44/n556 ),
    .Y(\i44/n576 ));
 AND2x2_ASAP7_75t_SL \i44/i585  (.A(\i44/n577 ),
    .B(\i44/n469 ),
    .Y(\i44/n578 ));
 AOI21xp33_ASAP7_75t_SL \i44/i586  (.A1(\i44/n54 ),
    .A2(\i44/n75 ),
    .B(\i44/n135 ),
    .Y(\i44/n577 ));
 NAND3xp33_ASAP7_75t_SL \i44/i587  (.A(\i44/n579 ),
    .B(\i44/n297 ),
    .C(\i44/n368 ),
    .Y(\i44/n580 ));
 AO21x1_ASAP7_75t_SL \i44/i588  (.A1(\i44/n566 ),
    .A2(\i44/n60 ),
    .B(\i44/n93 ),
    .Y(\i44/n579 ));
 NOR3xp33_ASAP7_75t_SL \i44/i589  (.A(\i44/n581 ),
    .B(\i44/n366 ),
    .C(\i44/n571 ),
    .Y(\i44/n582 ));
 INVxp67_ASAP7_75t_SL \i44/i59  (.A(\i44/n491 ),
    .Y(\i44/n492 ));
 OAI21xp5_ASAP7_75t_SL \i44/i590  (.A1(\i44/n73 ),
    .A2(\i44/n20 ),
    .B(\i44/n134 ),
    .Y(\i44/n581 ));
 INVx2_ASAP7_75t_SL \i44/i6  (.A(\i44/n18 ),
    .Y(\i44/n6 ));
 INVxp67_ASAP7_75t_SL \i44/i60  (.A(\i44/n487 ),
    .Y(\i44/n488 ));
 AND5x1_ASAP7_75t_SL \i44/i61  (.A(\i44/n408 ),
    .B(\i44/n576 ),
    .C(\i44/n400 ),
    .D(\i44/n319 ),
    .E(\i44/n290 ),
    .Y(\i44/n486 ));
 NOR3xp33_ASAP7_75t_SL \i44/i62  (.A(\i44/n420 ),
    .B(\i44/n399 ),
    .C(\i44/n381 ),
    .Y(\i44/n485 ));
 NOR3xp33_ASAP7_75t_SL \i44/i63  (.A(\i44/n443 ),
    .B(\i44/n382 ),
    .C(\i44/n331 ),
    .Y(\i44/n484 ));
 AND5x1_ASAP7_75t_SL \i44/i64  (.A(\i44/n371 ),
    .B(\i44/n385 ),
    .C(\i44/n364 ),
    .D(\i44/n374 ),
    .E(\i44/n299 ),
    .Y(\i44/n483 ));
 NOR2xp33_ASAP7_75t_SL \i44/i65  (.A(\i44/n444 ),
    .B(\i44/n449 ),
    .Y(\i44/n482 ));
 NAND4xp25_ASAP7_75t_SL \i44/i66  (.A(\i44/n428 ),
    .B(\i44/n541 ),
    .C(\i44/n439 ),
    .D(\i44/n424 ),
    .Y(\i44/n481 ));
 NAND5xp2_ASAP7_75t_SL \i44/i67  (.A(\i44/n407 ),
    .B(\i44/n362 ),
    .C(\i44/n259 ),
    .D(\i44/n244 ),
    .E(\i44/n15 ),
    .Y(\i44/n480 ));
 NOR4xp25_ASAP7_75t_SL \i44/i68  (.A(\i44/n397 ),
    .B(\i44/n567 ),
    .C(\i44/n347 ),
    .D(\i44/n323 ),
    .Y(\i44/n479 ));
 NAND4xp25_ASAP7_75t_SL \i44/i69  (.A(\i44/n417 ),
    .B(\i44/n430 ),
    .C(\i44/n542 ),
    .D(\i44/n434 ),
    .Y(\i44/n478 ));
 NOR2x2_ASAP7_75t_SL \i44/i7  (.A(\i44/n532 ),
    .B(\i44/n531 ),
    .Y(n32[4]));
 NAND4xp25_ASAP7_75t_SL \i44/i70  (.A(\i44/n441 ),
    .B(\i44/n439 ),
    .C(\i44/n544 ),
    .D(\i44/n289 ),
    .Y(\i44/n477 ));
 NAND3xp33_ASAP7_75t_SL \i44/i71  (.A(\i44/n434 ),
    .B(\i44/n406 ),
    .C(\i44/n23 ),
    .Y(\i44/n491 ));
 NAND4xp75_ASAP7_75t_SL \i44/i72  (.A(\i44/n338 ),
    .B(\i44/n308 ),
    .C(\i44/n393 ),
    .D(\i44/n26 ),
    .Y(\i44/n490 ));
 NAND2xp33_ASAP7_75t_L \i44/i73  (.A(\i44/n416 ),
    .B(\i44/n474 ),
    .Y(\i44/n476 ));
 AND2x2_ASAP7_75t_SL \i44/i74  (.A(\i44/n419 ),
    .B(\i44/n464 ),
    .Y(\i44/n489 ));
 NAND2x1p5_ASAP7_75t_SL \i44/i75  (.A(\i44/n471 ),
    .B(\i44/n429 ),
    .Y(\i44/n487 ));
 INVxp67_ASAP7_75t_SL \i44/i76  (.A(\i44/n474 ),
    .Y(\i44/n475 ));
 NOR5xp2_ASAP7_75t_SL \i44/i77  (.A(\i44/n357 ),
    .B(\i44/n330 ),
    .C(\i44/n251 ),
    .D(\i44/n211 ),
    .E(\i44/n555 ),
    .Y(\i44/n467 ));
 NOR3xp33_ASAP7_75t_SL \i44/i78  (.A(\i44/n438 ),
    .B(\i44/n352 ),
    .C(\i44/n344 ),
    .Y(\i44/n466 ));
 NOR2xp33_ASAP7_75t_SL \i44/i79  (.A(\i44/n396 ),
    .B(\i44/n418 ),
    .Y(\i44/n465 ));
 NOR2x2_ASAP7_75t_SL \i44/i8  (.A(\i44/n527 ),
    .B(\i44/n533 ),
    .Y(n32[3]));
 NOR2xp33_ASAP7_75t_SL \i44/i80  (.A(\i44/n436 ),
    .B(\i44/n387 ),
    .Y(\i44/n464 ));
 NOR2x1_ASAP7_75t_SL \i44/i81  (.A(\i44/n401 ),
    .B(\i44/n372 ),
    .Y(\i44/n474 ));
 NAND3xp33_ASAP7_75t_SL \i44/i82  (.A(\i44/n341 ),
    .B(\i44/n370 ),
    .C(\i44/n253 ),
    .Y(\i44/n463 ));
 NAND2xp5_ASAP7_75t_L \i44/i83  (.A(\i44/n435 ),
    .B(\i44/n405 ),
    .Y(\i44/n462 ));
 NAND2xp5_ASAP7_75t_SL \i44/i84  (.A(\i44/n386 ),
    .B(\i44/n427 ),
    .Y(\i44/n461 ));
 NAND3xp33_ASAP7_75t_SL \i44/i85  (.A(\i44/n576 ),
    .B(\i44/n325 ),
    .C(\i44/n569 ),
    .Y(\i44/n473 ));
 NOR3xp33_ASAP7_75t_SL \i44/i86  (.A(\i44/n409 ),
    .B(\i44/n8 ),
    .C(\i44/n306 ),
    .Y(\i44/n460 ));
 NAND2xp5_ASAP7_75t_SL \i44/i87  (.A(\i44/n25 ),
    .B(\i44/n417 ),
    .Y(\i44/n472 ));
 OR3x1_ASAP7_75t_SL \i44/i88  (.A(\i44/n333 ),
    .B(\i44/n346 ),
    .C(\i44/n29 ),
    .Y(\i44/n459 ));
 NOR2x1_ASAP7_75t_SL \i44/i89  (.A(\i44/n344 ),
    .B(\i44/n438 ),
    .Y(\i44/n471 ));
 AND5x2_ASAP7_75t_SL \i44/i9  (.A(\i44/n525 ),
    .B(\i44/n516 ),
    .C(\i44/n518 ),
    .D(\i44/n503 ),
    .E(\i44/n495 ),
    .Y(n32[6]));
 NOR2xp33_ASAP7_75t_L \i44/i90  (.A(\i44/n398 ),
    .B(\i44/n384 ),
    .Y(\i44/n470 ));
 NOR2xp33_ASAP7_75t_L \i44/i91  (.A(\i44/n550 ),
    .B(\i44/n426 ),
    .Y(\i44/n469 ));
 NOR3x1_ASAP7_75t_SL \i44/i92  (.A(\i44/n340 ),
    .B(\i44/n225 ),
    .C(\i44/n390 ),
    .Y(\i44/n468 ));
 NOR3xp33_ASAP7_75t_SL \i44/i93  (.A(\i44/n348 ),
    .B(\i44/n258 ),
    .C(\i44/n336 ),
    .Y(\i44/n455 ));
 NOR2xp33_ASAP7_75t_SL \i44/i94  (.A(\i44/n580 ),
    .B(\i44/n412 ),
    .Y(\i44/n454 ));
 NAND3xp33_ASAP7_75t_SL \i44/i95  (.A(\i44/n332 ),
    .B(\i44/n403 ),
    .C(\i44/n345 ),
    .Y(\i44/n453 ));
 NAND4xp25_ASAP7_75t_SL \i44/i96  (.A(\i44/n314 ),
    .B(\i44/n329 ),
    .C(\i44/n358 ),
    .D(\i44/n324 ),
    .Y(\i44/n452 ));
 NAND2x1_ASAP7_75t_SL \i44/i97  (.A(\i44/n425 ),
    .B(\i44/n437 ),
    .Y(\i44/n458 ));
 NOR5xp2_ASAP7_75t_SL \i44/i98  (.A(\i44/n433 ),
    .B(\i44/n350 ),
    .C(\i44/n147 ),
    .D(\i44/n570 ),
    .E(\i44/n191 ),
    .Y(\i44/n451 ));
 NAND3xp33_ASAP7_75t_SL \i44/i99  (.A(\i44/n389 ),
    .B(\i44/n410 ),
    .C(\i44/n261 ),
    .Y(\i44/n450 ));
 XOR2xp5_ASAP7_75t_SL i440 (.A(n1163),
    .B(n969),
    .Y(n1032));
 XNOR2xp5_ASAP7_75t_SL i441 (.A(n811),
    .B(n1192),
    .Y(n1031));
 AOI31xp33_ASAP7_75t_SL i442 (.A1(n819),
    .A2(n878),
    .A3(n1[3]),
    .B(n294),
    .Y(n1030));
 A2O1A1O1Ixp25_ASAP7_75t_SL i443 (.A1(n1[0]),
    .A2(n1[1]),
    .B(n292),
    .C(n819),
    .D(n294),
    .Y(n1029));
 A2O1A1Ixp33_ASAP7_75t_SL i444 (.A1(n1[2]),
    .A2(n293),
    .B(n877),
    .C(n819),
    .Y(n1028));
 AOI21xp5_ASAP7_75t_SL i445 (.A1(n819),
    .A2(n172),
    .B(n294),
    .Y(n1027));
 OAI22xp5_ASAP7_75t_SL i446 (.A1(n874),
    .A2(n125),
    .B1(n475),
    .B2(n221),
    .Y(n1026));
 OAI22xp5_ASAP7_75t_SL i447 (.A1(n873),
    .A2(n509),
    .B1(n872),
    .B2(n508),
    .Y(n1025));
 OAI22xp5_ASAP7_75t_SL i448 (.A1(n867),
    .A2(n788),
    .B1(n866),
    .B2(n787),
    .Y(n1024));
 OAI22xp5_ASAP7_75t_L i449 (.A1(n865),
    .A2(n800),
    .B1(n801),
    .B2(n864),
    .Y(n1023));
 INVx1_ASAP7_75t_SL \i45/i0  (.A(n31[7]),
    .Y(\i45/n0 ));
 INVx2_ASAP7_75t_SL \i45/i1  (.A(n31[5]),
    .Y(\i45/n1 ));
 NOR2x2_ASAP7_75t_SL \i45/i10  (.A(\i45/n556 ),
    .B(\i45/n562 ),
    .Y(n30[3]));
 NAND3xp33_ASAP7_75t_SL \i45/i100  (.A(\i45/n415 ),
    .B(\i45/n437 ),
    .C(\i45/n279 ),
    .Y(\i45/n480 ));
 NAND2xp33_ASAP7_75t_SL \i45/i101  (.A(\i45/n348 ),
    .B(\i45/n459 ),
    .Y(\i45/n479 ));
 NOR5xp2_ASAP7_75t_SL \i45/i102  (.A(\i45/n398 ),
    .B(\i45/n357 ),
    .C(\i45/n381 ),
    .D(\i45/n320 ),
    .E(\i45/n266 ),
    .Y(\i45/n478 ));
 NAND5xp2_ASAP7_75t_SL \i45/i103  (.A(\i45/n333 ),
    .B(\i45/n413 ),
    .C(\i45/n255 ),
    .D(\i45/n379 ),
    .E(\i45/n316 ),
    .Y(\i45/n477 ));
 NAND3xp33_ASAP7_75t_L \i45/i104  (.A(\i45/n326 ),
    .B(\i45/n363 ),
    .C(\i45/n442 ),
    .Y(\i45/n476 ));
 NOR5xp2_ASAP7_75t_SL \i45/i105  (.A(\i45/n324 ),
    .B(\i45/n339 ),
    .C(\i45/n314 ),
    .D(\i45/n139 ),
    .E(\i45/n115 ),
    .Y(\i45/n475 ));
 NAND5xp2_ASAP7_75t_SL \i45/i106  (.A(\i45/n32 ),
    .B(\i45/n414 ),
    .C(\i45/n255 ),
    .D(\i45/n111 ),
    .E(\i45/n227 ),
    .Y(\i45/n474 ));
 NAND4xp25_ASAP7_75t_SL \i45/i107  (.A(\i45/n260 ),
    .B(\i45/n274 ),
    .C(\i45/n385 ),
    .D(\i45/n22 ),
    .Y(\i45/n473 ));
 NOR5xp2_ASAP7_75t_SL \i45/i108  (.A(\i45/n280 ),
    .B(\i45/n329 ),
    .C(\i45/n265 ),
    .D(\i45/n221 ),
    .E(\i45/n219 ),
    .Y(\i45/n472 ));
 NOR2xp33_ASAP7_75t_SL \i45/i109  (.A(\i45/n431 ),
    .B(\i45/n466 ),
    .Y(\i45/n471 ));
 AND5x2_ASAP7_75t_SL \i45/i11  (.A(\i45/n554 ),
    .B(\i45/n545 ),
    .C(\i45/n547 ),
    .D(\i45/n532 ),
    .E(\i45/n524 ),
    .Y(n30[6]));
 NOR2xp33_ASAP7_75t_SL \i45/i110  (.A(\i45/n419 ),
    .B(\i45/n451 ),
    .Y(\i45/n470 ));
 NAND3x1_ASAP7_75t_SL \i45/i111  (.A(\i45/n278 ),
    .B(\i45/n449 ),
    .C(\i45/n413 ),
    .Y(\i45/n487 ));
 NAND3x1_ASAP7_75t_SL \i45/i112  (.A(\i45/n408 ),
    .B(\i45/n386 ),
    .C(\i45/n349 ),
    .Y(\i45/n486 ));
 AOI21xp5_ASAP7_75t_L \i45/i113  (.A1(\i45/n90 ),
    .A2(\i45/n283 ),
    .B(\i45/n195 ),
    .Y(\i45/n462 ));
 NOR2xp33_ASAP7_75t_SL \i45/i114  (.A(\i45/n398 ),
    .B(\i45/n354 ),
    .Y(\i45/n461 ));
 NAND2xp5_ASAP7_75t_SL \i45/i115  (.A(\i45/n384 ),
    .B(\i45/n418 ),
    .Y(\i45/n460 ));
 NOR2xp33_ASAP7_75t_SL \i45/i116  (.A(\i45/n417 ),
    .B(\i45/n573 ),
    .Y(\i45/n459 ));
 NOR2xp33_ASAP7_75t_SL \i45/i117  (.A(\i45/n392 ),
    .B(\i45/n403 ),
    .Y(\i45/n458 ));
 NOR2xp67_ASAP7_75t_SL \i45/i118  (.A(\i45/n205 ),
    .B(\i45/n400 ),
    .Y(\i45/n457 ));
 NOR2xp33_ASAP7_75t_L \i45/i119  (.A(\i45/n28 ),
    .B(\i45/n398 ),
    .Y(\i45/n456 ));
 AND3x4_ASAP7_75t_SL \i45/i12  (.A(\i45/n554 ),
    .B(\i45/n563 ),
    .C(\i45/n542 ),
    .Y(n30[1]));
 NOR4xp25_ASAP7_75t_SL \i45/i120  (.A(\i45/n30 ),
    .B(\i45/n367 ),
    .C(\i45/n28 ),
    .D(\i45/n215 ),
    .Y(\i45/n455 ));
 NAND2xp5_ASAP7_75t_SL \i45/i121  (.A(\i45/n310 ),
    .B(\i45/n376 ),
    .Y(\i45/n454 ));
 NOR4xp25_ASAP7_75t_SL \i45/i122  (.A(\i45/n135 ),
    .B(\i45/n302 ),
    .C(\i45/n268 ),
    .D(\i45/n284 ),
    .Y(\i45/n453 ));
 NOR3xp33_ASAP7_75t_SL \i45/i123  (.A(\i45/n307 ),
    .B(\i45/n258 ),
    .C(\i45/n306 ),
    .Y(\i45/n452 ));
 NAND2xp33_ASAP7_75t_SL \i45/i124  (.A(\i45/n362 ),
    .B(\i45/n29 ),
    .Y(\i45/n451 ));
 NOR2xp33_ASAP7_75t_SL \i45/i125  (.A(\i45/n354 ),
    .B(\i45/n356 ),
    .Y(\i45/n450 ));
 NOR2x1p5_ASAP7_75t_SL \i45/i126  (.A(\i45/n334 ),
    .B(\i45/n361 ),
    .Y(\i45/n449 ));
 NAND2xp33_ASAP7_75t_SL \i45/i127  (.A(\i45/n415 ),
    .B(\i45/n396 ),
    .Y(\i45/n448 ));
 NAND3xp33_ASAP7_75t_SL \i45/i128  (.A(\i45/n31 ),
    .B(\i45/n256 ),
    .C(\i45/n290 ),
    .Y(\i45/n447 ));
 NOR3xp33_ASAP7_75t_SL \i45/i129  (.A(\i45/n261 ),
    .B(\i45/n275 ),
    .C(\i45/n237 ),
    .Y(\i45/n469 ));
 NOR2x1p5_ASAP7_75t_SL \i45/i13  (.A(\i45/n564 ),
    .B(\i45/n555 ),
    .Y(n30[5]));
 NAND2xp5_ASAP7_75t_SL \i45/i130  (.A(\i45/n366 ),
    .B(\i45/n260 ),
    .Y(\i45/n468 ));
 NOR2x1_ASAP7_75t_SL \i45/i131  (.A(\i45/n332 ),
    .B(\i45/n359 ),
    .Y(\i45/n467 ));
 NAND2xp5_ASAP7_75t_SL \i45/i132  (.A(\i45/n255 ),
    .B(\i45/n368 ),
    .Y(\i45/n466 ));
 NOR2x1_ASAP7_75t_SL \i45/i133  (.A(\i45/n335 ),
    .B(\i45/n401 ),
    .Y(\i45/n465 ));
 NOR2x1_ASAP7_75t_SL \i45/i134  (.A(\i45/n30 ),
    .B(\i45/n354 ),
    .Y(\i45/n464 ));
 NOR3x1_ASAP7_75t_SL \i45/i135  (.A(\i45/n265 ),
    .B(\i45/n252 ),
    .C(\i45/n217 ),
    .Y(\i45/n463 ));
 INVx1_ASAP7_75t_SL \i45/i136  (.A(\i45/n444 ),
    .Y(\i45/n445 ));
 INVx1_ASAP7_75t_SL \i45/i137  (.A(\i45/n34 ),
    .Y(\i45/n443 ));
 NOR4xp25_ASAP7_75t_SL \i45/i138  (.A(\i45/n241 ),
    .B(\i45/n287 ),
    .C(\i45/n273 ),
    .D(\i45/n233 ),
    .Y(\i45/n442 ));
 AOI211xp5_ASAP7_75t_SL \i45/i139  (.A1(\i45/n89 ),
    .A2(\i45/n84 ),
    .B(\i45/n361 ),
    .C(\i45/n211 ),
    .Y(\i45/n441 ));
 AND2x2_ASAP7_75t_SL \i45/i14  (.A(\i45/n565 ),
    .B(\i45/n548 ),
    .Y(n30[0]));
 AOI211xp5_ASAP7_75t_SL \i45/i140  (.A1(\i45/n142 ),
    .A2(\i45/n67 ),
    .B(\i45/n380 ),
    .C(\i45/n305 ),
    .Y(\i45/n440 ));
 NAND2xp33_ASAP7_75t_SL \i45/i141  (.A(\i45/n350 ),
    .B(\i45/n378 ),
    .Y(\i45/n439 ));
 NAND5xp2_ASAP7_75t_SL \i45/i142  (.A(\i45/n285 ),
    .B(\i45/n300 ),
    .C(\i45/n312 ),
    .D(\i45/n213 ),
    .E(\i45/n136 ),
    .Y(\i45/n438 ));
 NOR4xp25_ASAP7_75t_SL \i45/i143  (.A(\i45/n388 ),
    .B(\i45/n175 ),
    .C(\i45/n177 ),
    .D(\i45/n201 ),
    .Y(\i45/n437 ));
 OAI221xp5_ASAP7_75t_SL \i45/i144  (.A1(\i45/n140 ),
    .A2(\i45/n106 ),
    .B1(\i45/n140 ),
    .B2(\i45/n19 ),
    .C(\i45/n362 ),
    .Y(\i45/n436 ));
 NOR2xp33_ASAP7_75t_SL \i45/i145  (.A(\i45/n340 ),
    .B(\i45/n344 ),
    .Y(\i45/n435 ));
 AOI211xp5_ASAP7_75t_SL \i45/i146  (.A1(\i45/n199 ),
    .A2(\i45/n571 ),
    .B(\i45/n322 ),
    .C(\i45/n223 ),
    .Y(\i45/n434 ));
 OA21x2_ASAP7_75t_SL \i45/i147  (.A1(\i45/n73 ),
    .A2(\i45/n90 ),
    .B(\i45/n414 ),
    .Y(\i45/n433 ));
 NOR4xp25_ASAP7_75t_SL \i45/i148  (.A(\i45/n315 ),
    .B(\i45/n210 ),
    .C(\i45/n247 ),
    .D(\i45/n217 ),
    .Y(\i45/n432 ));
 NAND5xp2_ASAP7_75t_SL \i45/i149  (.A(\i45/n176 ),
    .B(\i45/n122 ),
    .C(\i45/n188 ),
    .D(\i45/n179 ),
    .E(\i45/n113 ),
    .Y(\i45/n431 ));
 NOR3xp33_ASAP7_75t_SL \i45/i15  (.A(\i45/n537 ),
    .B(\i45/n533 ),
    .C(\i45/n540 ),
    .Y(\i45/n565 ));
 NOR3xp33_ASAP7_75t_SL \i45/i150  (.A(\i45/n360 ),
    .B(\i45/n212 ),
    .C(\i45/n110 ),
    .Y(\i45/n430 ));
 NAND2xp5_ASAP7_75t_SL \i45/i151  (.A(\i45/n338 ),
    .B(\i45/n32 ),
    .Y(\i45/n429 ));
 NAND5xp2_ASAP7_75t_SL \i45/i152  (.A(\i45/n253 ),
    .B(\i45/n129 ),
    .C(\i45/n245 ),
    .D(\i45/n232 ),
    .E(\i45/n231 ),
    .Y(\i45/n428 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i45/i153  (.A1(\i45/n93 ),
    .A2(\i45/n117 ),
    .B(\i45/n95 ),
    .C(\i45/n328 ),
    .Y(\i45/n427 ));
 NAND4xp25_ASAP7_75t_SL \i45/i154  (.A(\i45/n374 ),
    .B(\i45/n301 ),
    .C(\i45/n137 ),
    .D(\i45/n214 ),
    .Y(\i45/n426 ));
 NAND5xp2_ASAP7_75t_SL \i45/i155  (.A(\i45/n200 ),
    .B(\i45/n178 ),
    .C(\i45/n292 ),
    .D(\i45/n132 ),
    .E(\i45/n126 ),
    .Y(\i45/n425 ));
 NAND2xp5_ASAP7_75t_SL \i45/i156  (.A(\i45/n337 ),
    .B(\i45/n365 ),
    .Y(\i45/n424 ));
 NAND3xp33_ASAP7_75t_SL \i45/i157  (.A(\i45/n358 ),
    .B(\i45/n112 ),
    .C(\i45/n119 ),
    .Y(\i45/n423 ));
 NAND2xp5_ASAP7_75t_SL \i45/i158  (.A(\i45/n413 ),
    .B(\i45/n278 ),
    .Y(\i45/n422 ));
 NOR2xp33_ASAP7_75t_L \i45/i159  (.A(\i45/n390 ),
    .B(\i45/n403 ),
    .Y(\i45/n446 ));
 NOR2x2_ASAP7_75t_SL \i45/i16  (.A(\i45/n557 ),
    .B(\i45/n558 ),
    .Y(n30[2]));
 NAND2xp5_ASAP7_75t_SL \i45/i160  (.A(\i45/n279 ),
    .B(\i45/n415 ),
    .Y(\i45/n421 ));
 NOR2x1p5_ASAP7_75t_SL \i45/i161  (.A(\i45/n342 ),
    .B(\i45/n394 ),
    .Y(\i45/n444 ));
 NAND3x1_ASAP7_75t_SL \i45/i162  (.A(\i45/n319 ),
    .B(\i45/n169 ),
    .C(\i45/n182 ),
    .Y(\i45/n34 ));
 INVxp67_ASAP7_75t_SL \i45/i163  (.A(\i45/n419 ),
    .Y(\i45/n420 ));
 INVxp67_ASAP7_75t_SL \i45/i164  (.A(\i45/n10 ),
    .Y(\i45/n418 ));
 INVxp67_ASAP7_75t_SL \i45/i165  (.A(\i45/n411 ),
    .Y(\i45/n412 ));
 INVxp67_ASAP7_75t_SL \i45/i166  (.A(\i45/n409 ),
    .Y(\i45/n410 ));
 INVx2_ASAP7_75t_SL \i45/i167  (.A(\i45/n407 ),
    .Y(\i45/n408 ));
 INVxp67_ASAP7_75t_SL \i45/i168  (.A(\i45/n405 ),
    .Y(\i45/n406 ));
 INVxp67_ASAP7_75t_SL \i45/i169  (.A(\i45/n401 ),
    .Y(\i45/n402 ));
 NAND4xp75_ASAP7_75t_SL \i45/i17  (.A(\i45/n523 ),
    .B(\i45/n543 ),
    .C(\i45/n521 ),
    .D(\i45/n575 ),
    .Y(\i45/n564 ));
 INVxp67_ASAP7_75t_SL \i45/i170  (.A(\i45/n33 ),
    .Y(\i45/n399 ));
 INVx1_ASAP7_75t_SL \i45/i171  (.A(\i45/n396 ),
    .Y(\i45/n397 ));
 OAI31xp33_ASAP7_75t_SL \i45/i172  (.A1(\i45/n571 ),
    .A2(\i45/n4 ),
    .A3(\i45/n68 ),
    .B(\i45/n63 ),
    .Y(\i45/n395 ));
 NAND2x1_ASAP7_75t_SL \i45/i173  (.A(\i45/n272 ),
    .B(\i45/n270 ),
    .Y(\i45/n394 ));
 NOR2xp33_ASAP7_75t_SL \i45/i174  (.A(\i45/n313 ),
    .B(\i45/n307 ),
    .Y(\i45/n393 ));
 NAND2xp33_ASAP7_75t_SL \i45/i175  (.A(\i45/n256 ),
    .B(\i45/n255 ),
    .Y(\i45/n392 ));
 OAI21xp5_ASAP7_75t_SL \i45/i176  (.A1(\i45/n66 ),
    .A2(\i45/n166 ),
    .B(\i45/n229 ),
    .Y(\i45/n391 ));
 NAND2xp5_ASAP7_75t_SL \i45/i177  (.A(\i45/n216 ),
    .B(\i45/n256 ),
    .Y(\i45/n390 ));
 AOI211xp5_ASAP7_75t_SL \i45/i178  (.A1(\i45/n104 ),
    .A2(\i45/n38 ),
    .B(\i45/n144 ),
    .C(\i45/n151 ),
    .Y(\i45/n389 ));
 AOI31xp33_ASAP7_75t_SL \i45/i179  (.A1(\i45/n66 ),
    .A2(\i45/n20 ),
    .A3(\i45/n79 ),
    .B(\i45/n59 ),
    .Y(\i45/n388 ));
 NOR3xp33_ASAP7_75t_SL \i45/i18  (.A(\i45/n541 ),
    .B(\i45/n506 ),
    .C(\i45/n551 ),
    .Y(\i45/n563 ));
 NOR3xp33_ASAP7_75t_SL \i45/i180  (.A(\i45/n258 ),
    .B(\i45/n165 ),
    .C(\i45/n149 ),
    .Y(\i45/n387 ));
 NOR3xp33_ASAP7_75t_SL \i45/i181  (.A(\i45/n141 ),
    .B(\i45/n158 ),
    .C(\i45/n313 ),
    .Y(\i45/n386 ));
 OAI31xp33_ASAP7_75t_R \i45/i182  (.A1(\i45/n61 ),
    .A2(\i45/n63 ),
    .A3(\i45/n87 ),
    .B(\i45/n104 ),
    .Y(\i45/n385 ));
 AOI221xp5_ASAP7_75t_SL \i45/i183  (.A1(\i45/n93 ),
    .A2(\i45/n107 ),
    .B1(\i45/n69 ),
    .B2(\i45/n81 ),
    .C(\i45/n234 ),
    .Y(\i45/n384 ));
 OAI31xp33_ASAP7_75t_R \i45/i184  (.A1(\i45/n571 ),
    .A2(\i45/n91 ),
    .A3(\i45/n93 ),
    .B(\i45/n87 ),
    .Y(\i45/n383 ));
 AOI21xp5_ASAP7_75t_R \i45/i185  (.A1(\i45/n195 ),
    .A2(\i45/n79 ),
    .B(\i45/n566 ),
    .Y(\i45/n419 ));
 AOI21xp5_ASAP7_75t_L \i45/i186  (.A1(\i45/n79 ),
    .A2(\i45/n206 ),
    .B(\i45/n103 ),
    .Y(\i45/n382 ));
 OAI221xp5_ASAP7_75t_SL \i45/i187  (.A1(\i45/n21 ),
    .A2(\i45/n106 ),
    .B1(\i45/n62 ),
    .B2(\i45/n71 ),
    .C(\i45/n267 ),
    .Y(\i45/n381 ));
 AOI21xp33_ASAP7_75t_SL \i45/i188  (.A1(\i45/n206 ),
    .A2(\i45/n60 ),
    .B(\i45/n92 ),
    .Y(\i45/n380 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i45/i189  (.A1(\i45/n101 ),
    .A2(\i45/n7 ),
    .B(\i45/n569 ),
    .C(\i45/n23 ),
    .Y(\i45/n379 ));
 NAND4xp75_ASAP7_75t_SL \i45/i19  (.A(\i45/n522 ),
    .B(\i45/n553 ),
    .C(\i45/n527 ),
    .D(\i45/n517 ),
    .Y(\i45/n562 ));
 NOR3xp33_ASAP7_75t_SL \i45/i190  (.A(\i45/n281 ),
    .B(\i45/n141 ),
    .C(\i45/n173 ),
    .Y(\i45/n378 ));
 NAND3xp33_ASAP7_75t_SL \i45/i191  (.A(\i45/n24 ),
    .B(\i45/n27 ),
    .C(\i45/n204 ),
    .Y(\i45/n377 ));
 AOI22xp33_ASAP7_75t_SL \i45/i192  (.A1(\i45/n190 ),
    .A2(\i45/n75 ),
    .B1(\i45/n81 ),
    .B2(\i45/n68 ),
    .Y(\i45/n376 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i45/i193  (.A1(\i45/n103 ),
    .A2(\i45/n64 ),
    .B(\i45/n86 ),
    .C(\i45/n145 ),
    .Y(\i45/n375 ));
 OAI21xp5_ASAP7_75t_SL \i45/i194  (.A1(\i45/n78 ),
    .A2(\i45/n197 ),
    .B(\i45/n571 ),
    .Y(\i45/n374 ));
 NAND4xp25_ASAP7_75t_SL \i45/i195  (.A(\i45/n220 ),
    .B(\i45/n214 ),
    .C(\i45/n180 ),
    .D(\i45/n183 ),
    .Y(\i45/n373 ));
 NAND2xp33_ASAP7_75t_SL \i45/i196  (.A(\i45/n295 ),
    .B(\i45/n172 ),
    .Y(\i45/n372 ));
 OAI211xp5_ASAP7_75t_SL \i45/i197  (.A1(\i45/n92 ),
    .A2(\i45/n85 ),
    .B(\i45/n185 ),
    .C(\i45/n189 ),
    .Y(\i45/n417 ));
 NOR2x1_ASAP7_75t_SL \i45/i198  (.A(\i45/n194 ),
    .B(\i45/n257 ),
    .Y(\i45/n416 ));
 NOR2xp33_ASAP7_75t_SL \i45/i199  (.A(\i45/n254 ),
    .B(\i45/n314 ),
    .Y(\i45/n415 ));
 INVx2_ASAP7_75t_SL \i45/i2  (.A(n31[2]),
    .Y(\i45/n2 ));
 AND3x4_ASAP7_75t_SL \i45/i20  (.A(\i45/n544 ),
    .B(\i45/n559 ),
    .C(\i45/n549 ),
    .Y(n30[7]));
 AO21x1_ASAP7_75t_SL \i45/i200  (.A1(\i45/n70 ),
    .A2(\i45/n193 ),
    .B(\i45/n174 ),
    .Y(\i45/n414 ));
 AOI21xp5_ASAP7_75t_SL \i45/i201  (.A1(\i45/n68 ),
    .A2(\i45/n78 ),
    .B(\i45/n322 ),
    .Y(\i45/n413 ));
 NOR2xp33_ASAP7_75t_SL \i45/i202  (.A(\i45/n298 ),
    .B(\i45/n315 ),
    .Y(\i45/n411 ));
 OAI211xp5_ASAP7_75t_SL \i45/i203  (.A1(\i45/n79 ),
    .A2(\i45/n92 ),
    .B(\i45/n229 ),
    .C(\i45/n230 ),
    .Y(\i45/n409 ));
 OR2x2_ASAP7_75t_SL \i45/i204  (.A(\i45/n243 ),
    .B(\i45/n271 ),
    .Y(\i45/n407 ));
 AOI21xp5_ASAP7_75t_SL \i45/i205  (.A1(\i45/n91 ),
    .A2(\i45/n80 ),
    .B(\i45/n311 ),
    .Y(\i45/n405 ));
 OAI211xp5_ASAP7_75t_SL \i45/i206  (.A1(\i45/n106 ),
    .A2(\i45/n96 ),
    .B(\i45/n225 ),
    .C(\i45/n160 ),
    .Y(\i45/n404 ));
 NAND2xp5_ASAP7_75t_SL \i45/i207  (.A(\i45/n316 ),
    .B(\i45/n317 ),
    .Y(\i45/n403 ));
 NAND2xp5_ASAP7_75t_SL \i45/i208  (.A(\i45/n31 ),
    .B(\i45/n238 ),
    .Y(\i45/n401 ));
 NAND2xp5_ASAP7_75t_SL \i45/i209  (.A(\i45/n294 ),
    .B(\i45/n323 ),
    .Y(\i45/n400 ));
 NAND4xp75_ASAP7_75t_SL \i45/i21  (.A(\i45/n526 ),
    .B(\i45/n578 ),
    .C(\i45/n535 ),
    .D(\i45/n552 ),
    .Y(\i45/n561 ));
 OAI221xp5_ASAP7_75t_SL \i45/i210  (.A1(\i45/n71 ),
    .A2(\i45/n82 ),
    .B1(\i45/n66 ),
    .B2(\i45/n70 ),
    .C(\i45/n25 ),
    .Y(\i45/n33 ));
 NAND2xp5_ASAP7_75t_SL \i45/i211  (.A(\i45/n222 ),
    .B(\i45/n249 ),
    .Y(\i45/n398 ));
 NOR2x1_ASAP7_75t_SL \i45/i212  (.A(\i45/n296 ),
    .B(\i45/n266 ),
    .Y(\i45/n396 ));
 INVxp67_ASAP7_75t_SL \i45/i213  (.A(\i45/n367 ),
    .Y(\i45/n368 ));
 INVx1_ASAP7_75t_SL \i45/i214  (.A(\i45/n363 ),
    .Y(\i45/n364 ));
 INVx1_ASAP7_75t_SL \i45/i215  (.A(\i45/n358 ),
    .Y(\i45/n359 ));
 NAND4xp25_ASAP7_75t_SL \i45/i216  (.A(\i45/n138 ),
    .B(\i45/n161 ),
    .C(\i45/n145 ),
    .D(\i45/n143 ),
    .Y(\i45/n353 ));
 AOI31xp33_ASAP7_75t_SL \i45/i217  (.A1(\i45/n162 ),
    .A2(\i45/n90 ),
    .A3(\i45/n59 ),
    .B(\i45/n60 ),
    .Y(\i45/n352 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i45/i218  (.A1(\i45/n569 ),
    .A2(\i45/n65 ),
    .B(\i45/n87 ),
    .C(\i45/n167 ),
    .Y(\i45/n351 ));
 NOR4xp25_ASAP7_75t_SL \i45/i219  (.A(\i45/n135 ),
    .B(\i45/n152 ),
    .C(\i45/n228 ),
    .D(\i45/n109 ),
    .Y(\i45/n350 ));
 NAND2x1_ASAP7_75t_SL \i45/i22  (.A(\i45/n514 ),
    .B(\i45/n545 ),
    .Y(\i45/n560 ));
 AOI211xp5_ASAP7_75t_SL \i45/i220  (.A1(\i45/n163 ),
    .A2(\i45/n570 ),
    .B(\i45/n212 ),
    .C(\i45/n120 ),
    .Y(\i45/n349 ));
 AOI21xp5_ASAP7_75t_SL \i45/i221  (.A1(\i45/n196 ),
    .A2(\i45/n569 ),
    .B(\i45/n286 ),
    .Y(\i45/n348 ));
 NOR2xp33_ASAP7_75t_L \i45/i222  (.A(\i45/n236 ),
    .B(\i45/n308 ),
    .Y(\i45/n347 ));
 OAI31xp33_ASAP7_75t_SL \i45/i223  (.A1(\i45/n75 ),
    .A2(\i45/n69 ),
    .A3(\i45/n104 ),
    .B(\i45/n80 ),
    .Y(\i45/n346 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i45/i224  (.A1(\i45/n92 ),
    .A2(\i45/n64 ),
    .B(\i45/n100 ),
    .C(\i45/n282 ),
    .Y(\i45/n345 ));
 OAI22xp5_ASAP7_75t_SL \i45/i225  (.A1(\i45/n96 ),
    .A2(\i45/n198 ),
    .B1(\i45/n85 ),
    .B2(\i45/n118 ),
    .Y(\i45/n344 ));
 NOR2xp33_ASAP7_75t_SL \i45/i226  (.A(\i45/n263 ),
    .B(\i45/n239 ),
    .Y(\i45/n343 ));
 OAI222xp33_ASAP7_75t_SL \i45/i227  (.A1(\i45/n103 ),
    .A2(\i45/n60 ),
    .B1(\i45/n64 ),
    .B2(\i45/n20 ),
    .C1(\i45/n90 ),
    .C2(\i45/n85 ),
    .Y(\i45/n342 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i45/i228  (.A1(\i45/n75 ),
    .A2(\i45/n72 ),
    .B(\i45/n7 ),
    .C(\i45/n208 ),
    .Y(\i45/n341 ));
 NAND2xp33_ASAP7_75t_L \i45/i229  (.A(\i45/n134 ),
    .B(\i45/n250 ),
    .Y(\i45/n340 ));
 NOR2xp67_ASAP7_75t_SL \i45/i23  (.A(\i45/n507 ),
    .B(\i45/n546 ),
    .Y(\i45/n559 ));
 NAND2xp33_ASAP7_75t_SL \i45/i230  (.A(\i45/n304 ),
    .B(\i45/n159 ),
    .Y(\i45/n339 ));
 AOI22xp5_ASAP7_75t_SL \i45/i231  (.A1(\i45/n91 ),
    .A2(\i45/n131 ),
    .B1(\i45/n570 ),
    .B2(\i45/n93 ),
    .Y(\i45/n338 ));
 OAI21xp33_ASAP7_75t_SL \i45/i232  (.A1(\i45/n142 ),
    .A2(\i45/n91 ),
    .B(\i45/n570 ),
    .Y(\i45/n337 ));
 OA21x2_ASAP7_75t_SL \i45/i233  (.A1(\i45/n60 ),
    .A2(\i45/n166 ),
    .B(\i45/n154 ),
    .Y(\i45/n336 ));
 NAND2xp5_ASAP7_75t_SL \i45/i234  (.A(\i45/n244 ),
    .B(\i45/n321 ),
    .Y(\i45/n335 ));
 NAND4xp25_ASAP7_75t_SL \i45/i235  (.A(\i45/n156 ),
    .B(\i45/n184 ),
    .C(\i45/n128 ),
    .D(\i45/n125 ),
    .Y(\i45/n334 ));
 AOI221xp5_ASAP7_75t_SL \i45/i236  (.A1(\i45/n81 ),
    .A2(\i45/n58 ),
    .B1(\i45/n65 ),
    .B2(\i45/n84 ),
    .C(\i45/n257 ),
    .Y(\i45/n333 ));
 OAI221xp5_ASAP7_75t_SL \i45/i237  (.A1(\i45/n105 ),
    .A2(\i45/n100 ),
    .B1(\i45/n88 ),
    .B2(\i45/n19 ),
    .C(\i45/n133 ),
    .Y(\i45/n371 ));
 OAI222xp33_ASAP7_75t_SL \i45/i238  (.A1(\i45/n12 ),
    .A2(\i45/n66 ),
    .B1(\i45/n71 ),
    .B2(\i45/n85 ),
    .C1(\i45/n88 ),
    .C2(\i45/n94 ),
    .Y(\i45/n332 ));
 OAI221xp5_ASAP7_75t_SL \i45/i239  (.A1(\i45/n103 ),
    .A2(\i45/n94 ),
    .B1(\i45/n88 ),
    .B2(\i45/n86 ),
    .C(\i45/n264 ),
    .Y(\i45/n331 ));
 NAND4xp75_ASAP7_75t_SL \i45/i24  (.A(\i45/n518 ),
    .B(\i45/n530 ),
    .C(\i45/n512 ),
    .D(\i45/n515 ),
    .Y(\i45/n558 ));
 AND3x1_ASAP7_75t_SL \i45/i240  (.A(\i45/n153 ),
    .B(\i45/n161 ),
    .C(\i45/n288 ),
    .Y(\i45/n330 ));
 AOI22xp5_ASAP7_75t_SL \i45/i241  (.A1(\i45/n102 ),
    .A2(\i45/n192 ),
    .B1(\i45/n78 ),
    .B2(\i45/n569 ),
    .Y(\i45/n370 ));
 AOI31xp33_ASAP7_75t_SL \i45/i242  (.A1(\i45/n66 ),
    .A2(\i45/n98 ),
    .A3(\i45/n86 ),
    .B(\i45/n70 ),
    .Y(\i45/n329 ));
 NAND2xp33_ASAP7_75t_SL \i45/i243  (.A(\i45/n246 ),
    .B(\i45/n289 ),
    .Y(\i45/n328 ));
 OAI221xp5_ASAP7_75t_SL \i45/i244  (.A1(\i45/n103 ),
    .A2(\i45/n98 ),
    .B1(\i45/n21 ),
    .B2(\i45/n20 ),
    .C(\i45/n303 ),
    .Y(\i45/n327 ));
 OAI222xp33_ASAP7_75t_SL \i45/i245  (.A1(\i45/n96 ),
    .A2(\i45/n98 ),
    .B1(\i45/n105 ),
    .B2(\i45/n94 ),
    .C1(\i45/n21 ),
    .C2(\i45/n79 ),
    .Y(\i45/n369 ));
 NAND3x1_ASAP7_75t_SL \i45/i246  (.A(\i45/n251 ),
    .B(\i45/n187 ),
    .C(\i45/n181 ),
    .Y(\i45/n367 ));
 AOI22xp5_ASAP7_75t_SL \i45/i247  (.A1(\i45/n186 ),
    .A2(\i45/n104 ),
    .B1(\i45/n69 ),
    .B2(\i45/n87 ),
    .Y(\i45/n366 ));
 AOI22xp5_ASAP7_75t_SL \i45/i248  (.A1(\i45/n107 ),
    .A2(\i45/n123 ),
    .B1(\i45/n61 ),
    .B2(\i45/n571 ),
    .Y(\i45/n365 ));
 AOI221x1_ASAP7_75t_SL \i45/i249  (.A1(\i45/n104 ),
    .A2(\i45/n87 ),
    .B1(\i45/n93 ),
    .B2(\i45/n95 ),
    .C(\i45/n291 ),
    .Y(\i45/n363 ));
 OR3x1_ASAP7_75t_SL \i45/i25  (.A(\i45/n538 ),
    .B(\i45/n536 ),
    .C(\i45/n519 ),
    .Y(\i45/n557 ));
 AOI211x1_ASAP7_75t_SL \i45/i250  (.A1(\i45/n124 ),
    .A2(\i45/n83 ),
    .B(\i45/n226 ),
    .C(\i45/n228 ),
    .Y(\i45/n362 ));
 AO21x2_ASAP7_75t_SL \i45/i251  (.A1(\i45/n570 ),
    .A2(\i45/n4 ),
    .B(\i45/n259 ),
    .Y(\i45/n361 ));
 OAI21xp5_ASAP7_75t_SL \i45/i252  (.A1(\i45/n59 ),
    .A2(\i45/n100 ),
    .B(\i45/n299 ),
    .Y(\i45/n360 ));
 NOR2x1_ASAP7_75t_SL \i45/i253  (.A(\i45/n155 ),
    .B(\i45/n242 ),
    .Y(\i45/n358 ));
 OAI221xp5_ASAP7_75t_SL \i45/i254  (.A1(\i45/n26 ),
    .A2(\i45/n105 ),
    .B1(\i45/n76 ),
    .B2(\i45/n86 ),
    .C(\i45/n202 ),
    .Y(\i45/n357 ));
 OAI211xp5_ASAP7_75t_SL \i45/i255  (.A1(\i45/n86 ),
    .A2(\i45/n127 ),
    .B(\i45/n137 ),
    .C(\i45/n168 ),
    .Y(\i45/n356 ));
 NOR2x1_ASAP7_75t_SL \i45/i256  (.A(\i45/n167 ),
    .B(\i45/n248 ),
    .Y(\i45/n32 ));
 NOR2xp33_ASAP7_75t_SL \i45/i257  (.A(\i45/n170 ),
    .B(\i45/n318 ),
    .Y(\i45/n326 ));
 AOI222xp33_ASAP7_75t_SL \i45/i258  (.A1(\i45/n93 ),
    .A2(\i45/n81 ),
    .B1(\i45/n7 ),
    .B2(\i45/n58 ),
    .C1(\i45/n571 ),
    .C2(\i45/n78 ),
    .Y(\i45/n355 ));
 OAI221xp5_ASAP7_75t_SL \i45/i259  (.A1(\i45/n73 ),
    .A2(\i45/n64 ),
    .B1(\i45/n70 ),
    .B2(\i45/n60 ),
    .C(\i45/n148 ),
    .Y(\i45/n354 ));
 OR3x1_ASAP7_75t_SL \i45/i26  (.A(\i45/n539 ),
    .B(\i45/n505 ),
    .C(\i45/n480 ),
    .Y(\i45/n556 ));
 INVx1_ASAP7_75t_SL \i45/i260  (.A(\i45/n323 ),
    .Y(\i45/n324 ));
 INVx1_ASAP7_75t_SL \i45/i261  (.A(\i45/n320 ),
    .Y(\i45/n321 ));
 INVx1_ASAP7_75t_SL \i45/i262  (.A(\i45/n318 ),
    .Y(\i45/n319 ));
 INVxp67_ASAP7_75t_SL \i45/i263  (.A(\i45/n311 ),
    .Y(\i45/n312 ));
 INVx1_ASAP7_75t_SL \i45/i264  (.A(\i45/n308 ),
    .Y(\i45/n309 ));
 OAI21xp33_ASAP7_75t_SL \i45/i265  (.A1(\i45/n567 ),
    .A2(\i45/n77 ),
    .B(\i45/n218 ),
    .Y(\i45/n306 ));
 NAND2xp5_ASAP7_75t_SL \i45/i266  (.A(\i45/n116 ),
    .B(\i45/n160 ),
    .Y(\i45/n305 ));
 OAI21xp5_ASAP7_75t_SL \i45/i267  (.A1(\i45/n69 ),
    .A2(\i45/n68 ),
    .B(\i45/n101 ),
    .Y(\i45/n304 ));
 NOR2xp33_ASAP7_75t_SL \i45/i268  (.A(\i45/n171 ),
    .B(\i45/n211 ),
    .Y(\i45/n303 ));
 NAND2xp33_ASAP7_75t_L \i45/i269  (.A(\i45/n207 ),
    .B(\i45/n121 ),
    .Y(\i45/n302 ));
 NAND3xp33_ASAP7_75t_SL \i45/i27  (.A(\i45/n550 ),
    .B(\i45/n535 ),
    .C(\i45/n518 ),
    .Y(\i45/n555 ));
 OAI21xp33_ASAP7_75t_SL \i45/i270  (.A1(\i45/n89 ),
    .A2(\i45/n72 ),
    .B(\i45/n63 ),
    .Y(\i45/n301 ));
 NOR2xp33_ASAP7_75t_SL \i45/i271  (.A(\i45/n23 ),
    .B(\i45/n146 ),
    .Y(\i45/n300 ));
 OAI21xp5_ASAP7_75t_SL \i45/i272  (.A1(\i45/n91 ),
    .A2(\i45/n99 ),
    .B(\i45/n81 ),
    .Y(\i45/n299 ));
 OAI21xp5_ASAP7_75t_SL \i45/i273  (.A1(\i45/n73 ),
    .A2(\i45/n566 ),
    .B(\i45/n209 ),
    .Y(\i45/n298 ));
 AOI22xp5_ASAP7_75t_SL \i45/i274  (.A1(\i45/n101 ),
    .A2(\i45/n72 ),
    .B1(\i45/n95 ),
    .B2(\i45/n571 ),
    .Y(\i45/n297 ));
 OAI21xp5_ASAP7_75t_SL \i45/i275  (.A1(\i45/n20 ),
    .A2(\i45/n88 ),
    .B(\i45/n164 ),
    .Y(\i45/n296 ));
 OAI21xp5_ASAP7_75t_SL \i45/i276  (.A1(\i45/n91 ),
    .A2(\i45/n68 ),
    .B(\i45/n84 ),
    .Y(\i45/n295 ));
 AOI22xp5_ASAP7_75t_R \i45/i277  (.A1(\i45/n58 ),
    .A2(\i45/n107 ),
    .B1(\i45/n61 ),
    .B2(\i45/n91 ),
    .Y(\i45/n294 ));
 OA21x2_ASAP7_75t_SL \i45/i278  (.A1(\i45/n82 ),
    .A2(\i45/n18 ),
    .B(\i45/n213 ),
    .Y(\i45/n325 ));
 AOI21xp33_ASAP7_75t_SL \i45/i279  (.A1(\i45/n85 ),
    .A2(\i45/n82 ),
    .B(\i45/n59 ),
    .Y(\i45/n293 ));
 NOR2x1_ASAP7_75t_SL \i45/i28  (.A(\i45/n460 ),
    .B(\i45/n536 ),
    .Y(\i45/n553 ));
 OAI21xp5_ASAP7_75t_SL \i45/i280  (.A1(\i45/n95 ),
    .A2(\i45/n107 ),
    .B(\i45/n102 ),
    .Y(\i45/n292 ));
 OA21x2_ASAP7_75t_SL \i45/i281  (.A1(\i45/n7 ),
    .A2(\i45/n107 ),
    .B(\i45/n569 ),
    .Y(\i45/n291 ));
 AOI22xp33_ASAP7_75t_SL \i45/i282  (.A1(\i45/n107 ),
    .A2(\i45/n69 ),
    .B1(\i45/n83 ),
    .B2(\i45/n4 ),
    .Y(\i45/n290 ));
 OAI21xp5_ASAP7_75t_SL \i45/i283  (.A1(\i45/n84 ),
    .A2(\i45/n61 ),
    .B(\i45/n102 ),
    .Y(\i45/n289 ));
 OAI21xp5_ASAP7_75t_SL \i45/i284  (.A1(\i45/n91 ),
    .A2(\i45/n89 ),
    .B(\i45/n107 ),
    .Y(\i45/n288 ));
 AOI21xp33_ASAP7_75t_SL \i45/i285  (.A1(\i45/n79 ),
    .A2(\i45/n100 ),
    .B(\i45/n59 ),
    .Y(\i45/n287 ));
 OAI21xp5_ASAP7_75t_SL \i45/i286  (.A1(\i45/n73 ),
    .A2(\i45/n88 ),
    .B(\i45/n29 ),
    .Y(\i45/n286 ));
 AOI22xp5_ASAP7_75t_SL \i45/i287  (.A1(\i45/n78 ),
    .A2(\i45/n75 ),
    .B1(\i45/n95 ),
    .B2(\i45/n72 ),
    .Y(\i45/n285 ));
 AOI21xp33_ASAP7_75t_SL \i45/i288  (.A1(\i45/n92 ),
    .A2(\i45/n59 ),
    .B(\i45/n86 ),
    .Y(\i45/n284 ));
 OAI21xp5_ASAP7_75t_SL \i45/i289  (.A1(\i45/n569 ),
    .A2(\i45/n91 ),
    .B(\i45/n63 ),
    .Y(\i45/n283 ));
 NOR2x1_ASAP7_75t_SL \i45/i29  (.A(\i45/n520 ),
    .B(\i45/n516 ),
    .Y(\i45/n552 ));
 OAI21xp5_ASAP7_75t_SL \i45/i290  (.A1(\i45/n89 ),
    .A2(\i45/n75 ),
    .B(\i45/n95 ),
    .Y(\i45/n282 ));
 NAND2xp5_ASAP7_75t_SL \i45/i291  (.A(\i45/n102 ),
    .B(\i45/n196 ),
    .Y(\i45/n31 ));
 AOI22xp5_ASAP7_75t_SL \i45/i292  (.A1(\i45/n568 ),
    .A2(\i45/n97 ),
    .B1(\i45/n95 ),
    .B2(\i45/n4 ),
    .Y(\i45/n323 ));
 NAND2xp5_ASAP7_75t_L \i45/i293  (.A(\i45/n229 ),
    .B(\i45/n230 ),
    .Y(\i45/n281 ));
 OAI22xp5_ASAP7_75t_SL \i45/i294  (.A1(\i45/n77 ),
    .A2(\i45/n103 ),
    .B1(\i45/n108 ),
    .B2(\i45/n18 ),
    .Y(\i45/n322 ));
 OAI22xp5_ASAP7_75t_SL \i45/i295  (.A1(\i45/n108 ),
    .A2(\i45/n88 ),
    .B1(\i45/n21 ),
    .B2(\i45/n85 ),
    .Y(\i45/n320 ));
 OAI22xp5_ASAP7_75t_SL \i45/i296  (.A1(\i45/n106 ),
    .A2(\i45/n71 ),
    .B1(\i45/n73 ),
    .B2(\i45/n96 ),
    .Y(\i45/n318 ));
 AOI22xp5_ASAP7_75t_SL \i45/i297  (.A1(\i45/n83 ),
    .A2(\i45/n104 ),
    .B1(\i45/n7 ),
    .B2(\i45/n99 ),
    .Y(\i45/n317 ));
 AOI22xp5_ASAP7_75t_SL \i45/i298  (.A1(\i45/n83 ),
    .A2(\i45/n75 ),
    .B1(\i45/n568 ),
    .B2(\i45/n72 ),
    .Y(\i45/n316 ));
 OAI22xp5_ASAP7_75t_SL \i45/i299  (.A1(\i45/n86 ),
    .A2(\i45/n96 ),
    .B1(\i45/n88 ),
    .B2(\i45/n62 ),
    .Y(\i45/n315 ));
 INVx2_ASAP7_75t_SL \i45/i3  (.A(n31[0]),
    .Y(\i45/n3 ));
 NAND3xp33_ASAP7_75t_SL \i45/i30  (.A(\i45/n500 ),
    .B(\i45/n582 ),
    .C(\i45/n498 ),
    .Y(\i45/n551 ));
 OAI22xp5_ASAP7_75t_SL \i45/i300  (.A1(\i45/n108 ),
    .A2(\i45/n105 ),
    .B1(\i45/n60 ),
    .B2(\i45/n12 ),
    .Y(\i45/n314 ));
 NAND2xp5_ASAP7_75t_L \i45/i301  (.A(\i45/n22 ),
    .B(\i45/n191 ),
    .Y(\i45/n313 ));
 OAI22xp5_ASAP7_75t_SL \i45/i302  (.A1(\i45/n73 ),
    .A2(\i45/n105 ),
    .B1(\i45/n85 ),
    .B2(\i45/n566 ),
    .Y(\i45/n311 ));
 OAI21xp5_ASAP7_75t_SL \i45/i303  (.A1(\i45/n91 ),
    .A2(\i45/n65 ),
    .B(\i45/n101 ),
    .Y(\i45/n310 ));
 NOR2x1_ASAP7_75t_SL \i45/i304  (.A(\i45/n18 ),
    .B(\i45/n26 ),
    .Y(\i45/n308 ));
 NAND2xp33_ASAP7_75t_L \i45/i305  (.A(\i45/n137 ),
    .B(\i45/n168 ),
    .Y(\i45/n280 ));
 OAI21xp5_ASAP7_75t_SL \i45/i306  (.A1(\i45/n86 ),
    .A2(\i45/n71 ),
    .B(\i45/n136 ),
    .Y(\i45/n307 ));
 INVxp67_ASAP7_75t_SL \i45/i307  (.A(\i45/n276 ),
    .Y(\i45/n277 ));
 INVxp67_ASAP7_75t_SL \i45/i308  (.A(\i45/n274 ),
    .Y(\i45/n275 ));
 INVx1_ASAP7_75t_SL \i45/i309  (.A(\i45/n272 ),
    .Y(\i45/n273 ));
 NOR2xp33_ASAP7_75t_SL \i45/i31  (.A(\i45/n525 ),
    .B(\i45/n489 ),
    .Y(\i45/n550 ));
 INVx1_ASAP7_75t_SL \i45/i310  (.A(\i45/n269 ),
    .Y(\i45/n270 ));
 INVxp67_ASAP7_75t_SL \i45/i311  (.A(\i45/n267 ),
    .Y(\i45/n268 ));
 INVxp67_ASAP7_75t_R \i45/i312  (.A(\i45/n263 ),
    .Y(\i45/n264 ));
 INVxp67_ASAP7_75t_SL \i45/i313  (.A(\i45/n261 ),
    .Y(\i45/n262 ));
 OAI22xp33_ASAP7_75t_SL \i45/i314  (.A1(\i45/n62 ),
    .A2(\i45/n105 ),
    .B1(\i45/n70 ),
    .B2(\i45/n77 ),
    .Y(\i45/n254 ));
 OAI21xp5_ASAP7_75t_SL \i45/i315  (.A1(\i45/n72 ),
    .A2(\i45/n97 ),
    .B(\i45/n95 ),
    .Y(\i45/n253 ));
 OAI21xp33_ASAP7_75t_SL \i45/i316  (.A1(\i45/n19 ),
    .A2(\i45/n12 ),
    .B(\i45/n150 ),
    .Y(\i45/n252 ));
 OAI21xp5_ASAP7_75t_SL \i45/i317  (.A1(\i45/n74 ),
    .A2(\i45/n87 ),
    .B(\i45/n89 ),
    .Y(\i45/n251 ));
 OAI21xp5_ASAP7_75t_SL \i45/i318  (.A1(\i45/n69 ),
    .A2(\i45/n65 ),
    .B(\i45/n74 ),
    .Y(\i45/n250 ));
 AOI22xp5_ASAP7_75t_SL \i45/i319  (.A1(\i45/n570 ),
    .A2(\i45/n75 ),
    .B1(\i45/n63 ),
    .B2(\i45/n4 ),
    .Y(\i45/n249 ));
 NOR5xp2_ASAP7_75t_SL \i45/i32  (.A(\i45/n491 ),
    .B(\i45/n438 ),
    .C(\i45/n482 ),
    .D(\i45/n400 ),
    .E(\i45/n404 ),
    .Y(\i45/n549 ));
 OAI22xp5_ASAP7_75t_SL \i45/i320  (.A1(\i45/n105 ),
    .A2(\i45/n66 ),
    .B1(\i45/n62 ),
    .B2(\i45/n18 ),
    .Y(\i45/n248 ));
 AOI21xp33_ASAP7_75t_SL \i45/i321  (.A1(\i45/n88 ),
    .A2(\i45/n96 ),
    .B(\i45/n98 ),
    .Y(\i45/n247 ));
 OAI21xp5_ASAP7_75t_SL \i45/i322  (.A1(\i45/n58 ),
    .A2(\i45/n65 ),
    .B(\i45/n63 ),
    .Y(\i45/n246 ));
 OAI21xp5_ASAP7_75t_SL \i45/i323  (.A1(\i45/n570 ),
    .A2(\i45/n74 ),
    .B(\i45/n69 ),
    .Y(\i45/n245 ));
 AOI22xp33_ASAP7_75t_SL \i45/i324  (.A1(\i45/n83 ),
    .A2(\i45/n91 ),
    .B1(\i45/n7 ),
    .B2(\i45/n69 ),
    .Y(\i45/n244 ));
 OAI22xp33_ASAP7_75t_SL \i45/i325  (.A1(\i45/n77 ),
    .A2(\i45/n59 ),
    .B1(\i45/n103 ),
    .B2(\i45/n79 ),
    .Y(\i45/n243 ));
 AOI22xp5_ASAP7_75t_SL \i45/i326  (.A1(\i45/n568 ),
    .A2(\i45/n102 ),
    .B1(\i45/n101 ),
    .B2(\i45/n68 ),
    .Y(\i45/n279 ));
 OAI22xp33_ASAP7_75t_SL \i45/i327  (.A1(\i45/n21 ),
    .A2(\i45/n77 ),
    .B1(\i45/n96 ),
    .B2(\i45/n100 ),
    .Y(\i45/n242 ));
 OAI22xp5_ASAP7_75t_SL \i45/i328  (.A1(\i45/n106 ),
    .A2(\i45/n12 ),
    .B1(\i45/n19 ),
    .B2(\i45/n103 ),
    .Y(\i45/n241 ));
 OAI22xp5_ASAP7_75t_SL \i45/i329  (.A1(\i45/n79 ),
    .A2(\i45/n12 ),
    .B1(\i45/n100 ),
    .B2(\i45/n92 ),
    .Y(\i45/n240 ));
 NOR3xp33_ASAP7_75t_SL \i45/i33  (.A(\i45/n487 ),
    .B(\i45/n502 ),
    .C(\i45/n534 ),
    .Y(\i45/n548 ));
 AOI22xp5_ASAP7_75t_SL \i45/i330  (.A1(\i45/n58 ),
    .A2(\i45/n61 ),
    .B1(\i45/n568 ),
    .B2(\i45/n91 ),
    .Y(\i45/n278 ));
 OAI22xp33_ASAP7_75t_SL \i45/i331  (.A1(\i45/n64 ),
    .A2(\i45/n77 ),
    .B1(\i45/n18 ),
    .B2(\i45/n66 ),
    .Y(\i45/n239 ));
 AOI22xp5_ASAP7_75t_SL \i45/i332  (.A1(\i45/n81 ),
    .A2(\i45/n97 ),
    .B1(\i45/n61 ),
    .B2(\i45/n99 ),
    .Y(\i45/n238 ));
 OAI22xp5_ASAP7_75t_SL \i45/i333  (.A1(\i45/n77 ),
    .A2(\i45/n105 ),
    .B1(\i45/n85 ),
    .B2(\i45/n18 ),
    .Y(\i45/n237 ));
 OAI21xp5_ASAP7_75t_SL \i45/i334  (.A1(\i45/n94 ),
    .A2(\i45/n70 ),
    .B(\i45/n159 ),
    .Y(\i45/n236 ));
 OAI21xp5_ASAP7_75t_SL \i45/i335  (.A1(\i45/n60 ),
    .A2(\i45/n71 ),
    .B(\i45/n147 ),
    .Y(\i45/n276 ));
 AOI22xp5_ASAP7_75t_SL \i45/i336  (.A1(\i45/n58 ),
    .A2(\i45/n84 ),
    .B1(\i45/n61 ),
    .B2(\i45/n68 ),
    .Y(\i45/n274 ));
 AOI22xp5_ASAP7_75t_SL \i45/i337  (.A1(\i45/n63 ),
    .A2(\i45/n65 ),
    .B1(\i45/n75 ),
    .B2(\i45/n81 ),
    .Y(\i45/n272 ));
 OA21x2_ASAP7_75t_SL \i45/i338  (.A1(\i45/n66 ),
    .A2(\i45/n70 ),
    .B(\i45/n25 ),
    .Y(\i45/n235 ));
 OAI22xp5_ASAP7_75t_SL \i45/i339  (.A1(\i45/n66 ),
    .A2(\i45/n96 ),
    .B1(\i45/n85 ),
    .B2(\i45/n70 ),
    .Y(\i45/n271 ));
 NOR2x1_ASAP7_75t_SL \i45/i34  (.A(\i45/n531 ),
    .B(\i45/n492 ),
    .Y(\i45/n547 ));
 OAI22xp5_ASAP7_75t_SL \i45/i340  (.A1(\i45/n59 ),
    .A2(\i45/n19 ),
    .B1(\i45/n77 ),
    .B2(\i45/n90 ),
    .Y(\i45/n234 ));
 NAND2xp33_ASAP7_75t_SL \i45/i341  (.A(\i45/n231 ),
    .B(\i45/n232 ),
    .Y(\i45/n233 ));
 OAI22x1_ASAP7_75t_SL \i45/i342  (.A1(\i45/n20 ),
    .A2(\i45/n105 ),
    .B1(\i45/n62 ),
    .B2(\i45/n567 ),
    .Y(\i45/n269 ));
 AOI22xp5_ASAP7_75t_SL \i45/i343  (.A1(\i45/n63 ),
    .A2(\i45/n75 ),
    .B1(\i45/n61 ),
    .B2(\i45/n569 ),
    .Y(\i45/n267 ));
 AO22x2_ASAP7_75t_SL \i45/i344  (.A1(\i45/n107 ),
    .A2(\i45/n104 ),
    .B1(\i45/n67 ),
    .B2(\i45/n99 ),
    .Y(\i45/n266 ));
 OAI21xp5_ASAP7_75t_SL \i45/i345  (.A1(\i45/n94 ),
    .A2(\i45/n64 ),
    .B(\i45/n130 ),
    .Y(\i45/n265 ));
 OAI22xp33_ASAP7_75t_SL \i45/i346  (.A1(\i45/n98 ),
    .A2(\i45/n59 ),
    .B1(\i45/n96 ),
    .B2(\i45/n60 ),
    .Y(\i45/n263 ));
 OAI22xp5_ASAP7_75t_SL \i45/i347  (.A1(\i45/n79 ),
    .A2(\i45/n64 ),
    .B1(\i45/n85 ),
    .B2(\i45/n96 ),
    .Y(\i45/n261 ));
 AOI22xp5_ASAP7_75t_SL \i45/i348  (.A1(\i45/n58 ),
    .A2(\i45/n63 ),
    .B1(\i45/n87 ),
    .B2(\i45/n99 ),
    .Y(\i45/n260 ));
 OAI22xp5_ASAP7_75t_SL \i45/i349  (.A1(\i45/n92 ),
    .A2(\i45/n77 ),
    .B1(\i45/n90 ),
    .B2(\i45/n82 ),
    .Y(\i45/n259 ));
 NAND2xp5_ASAP7_75t_SL \i45/i35  (.A(\i45/n490 ),
    .B(\i45/n508 ),
    .Y(\i45/n546 ));
 OAI22xp5_ASAP7_75t_SL \i45/i350  (.A1(\i45/n66 ),
    .A2(\i45/n76 ),
    .B1(\i45/n85 ),
    .B2(\i45/n567 ),
    .Y(\i45/n258 ));
 OAI22xp5_ASAP7_75t_SL \i45/i351  (.A1(\i45/n82 ),
    .A2(\i45/n96 ),
    .B1(\i45/n86 ),
    .B2(\i45/n103 ),
    .Y(\i45/n30 ));
 OAI22xp5_ASAP7_75t_SL \i45/i352  (.A1(\i45/n66 ),
    .A2(\i45/n64 ),
    .B1(\i45/n70 ),
    .B2(\i45/n62 ),
    .Y(\i45/n257 ));
 AOI22xp5_ASAP7_75t_SL \i45/i353  (.A1(\i45/n74 ),
    .A2(\i45/n99 ),
    .B1(\i45/n61 ),
    .B2(\i45/n75 ),
    .Y(\i45/n256 ));
 AOI22xp5_ASAP7_75t_SL \i45/i354  (.A1(\i45/n568 ),
    .A2(\i45/n65 ),
    .B1(\i45/n80 ),
    .B2(\i45/n571 ),
    .Y(\i45/n255 ));
 INVxp67_ASAP7_75t_SL \i45/i355  (.A(\i45/n226 ),
    .Y(\i45/n227 ));
 INVx1_ASAP7_75t_SL \i45/i356  (.A(\i45/n224 ),
    .Y(\i45/n225 ));
 INVxp67_ASAP7_75t_SL \i45/i357  (.A(\i45/n222 ),
    .Y(\i45/n223 ));
 INVxp67_ASAP7_75t_SL \i45/i358  (.A(\i45/n220 ),
    .Y(\i45/n221 ));
 INVxp67_ASAP7_75t_SL \i45/i359  (.A(\i45/n218 ),
    .Y(\i45/n219 ));
 NOR3x1_ASAP7_75t_SL \i45/i36  (.A(\i45/n34 ),
    .B(\i45/n504 ),
    .C(\i45/n429 ),
    .Y(\i45/n554 ));
 INVxp67_ASAP7_75t_SL \i45/i360  (.A(\i45/n215 ),
    .Y(\i45/n216 ));
 INVxp67_ASAP7_75t_SL \i45/i361  (.A(\i45/n209 ),
    .Y(\i45/n210 ));
 INVxp67_ASAP7_75t_SL \i45/i362  (.A(\i45/n207 ),
    .Y(\i45/n208 ));
 INVxp67_ASAP7_75t_SL \i45/i363  (.A(\i45/n204 ),
    .Y(\i45/n205 ));
 INVxp67_ASAP7_75t_SL \i45/i364  (.A(\i45/n202 ),
    .Y(\i45/n203 ));
 INVxp67_ASAP7_75t_SL \i45/i365  (.A(\i45/n200 ),
    .Y(\i45/n201 ));
 INVxp67_ASAP7_75t_SL \i45/i366  (.A(\i45/n198 ),
    .Y(\i45/n199 ));
 INVxp67_ASAP7_75t_SL \i45/i367  (.A(\i45/n26 ),
    .Y(\i45/n197 ));
 INVx1_ASAP7_75t_SL \i45/i368  (.A(\i45/n196 ),
    .Y(\i45/n195 ));
 NAND2xp5_ASAP7_75t_SL \i45/i369  (.A(\i45/n84 ),
    .B(\i45/n102 ),
    .Y(\i45/n232 ));
 NOR3xp33_ASAP7_75t_SL \i45/i37  (.A(\i45/n448 ),
    .B(\i45/n34 ),
    .C(\i45/n528 ),
    .Y(\i45/n544 ));
 AND2x2_ASAP7_75t_SL \i45/i370  (.A(\i45/n67 ),
    .B(\i45/n571 ),
    .Y(\i45/n194 ));
 NAND2xp5_ASAP7_75t_SL \i45/i371  (.A(\i45/n101 ),
    .B(\i45/n99 ),
    .Y(\i45/n193 ));
 NAND2xp5_ASAP7_75t_SL \i45/i372  (.A(\i45/n100 ),
    .B(\i45/n98 ),
    .Y(\i45/n192 ));
 NAND2xp5_ASAP7_75t_SL \i45/i373  (.A(\i45/n61 ),
    .B(\i45/n104 ),
    .Y(\i45/n191 ));
 NAND2xp33_ASAP7_75t_SL \i45/i374  (.A(\i45/n79 ),
    .B(\i45/n73 ),
    .Y(\i45/n190 ));
 NAND2xp5_ASAP7_75t_SL \i45/i375  (.A(\i45/n72 ),
    .B(\i45/n78 ),
    .Y(\i45/n189 ));
 NAND2xp5_ASAP7_75t_SL \i45/i376  (.A(\i45/n72 ),
    .B(\i45/n81 ),
    .Y(\i45/n231 ));
 NAND2xp5_ASAP7_75t_SL \i45/i377  (.A(\i45/n78 ),
    .B(\i45/n89 ),
    .Y(\i45/n230 ));
 NAND2xp5_ASAP7_75t_SL \i45/i378  (.A(\i45/n81 ),
    .B(\i45/n102 ),
    .Y(\i45/n188 ));
 NAND2xp5_ASAP7_75t_SL \i45/i379  (.A(\i45/n4 ),
    .B(\i45/n78 ),
    .Y(\i45/n187 ));
 NOR2xp33_ASAP7_75t_SL \i45/i38  (.A(\i45/n509 ),
    .B(\i45/n34 ),
    .Y(\i45/n543 ));
 NAND2xp5_ASAP7_75t_SL \i45/i380  (.A(\i45/n85 ),
    .B(\i45/n19 ),
    .Y(\i45/n186 ));
 NAND2xp5_ASAP7_75t_SL \i45/i381  (.A(\i45/n101 ),
    .B(\i45/n569 ),
    .Y(\i45/n185 ));
 NAND2xp5_ASAP7_75t_SL \i45/i382  (.A(\i45/n84 ),
    .B(\i45/n4 ),
    .Y(\i45/n184 ));
 NAND2xp5_ASAP7_75t_SL \i45/i383  (.A(\i45/n571 ),
    .B(\i45/n87 ),
    .Y(\i45/n183 ));
 NAND2xp5_ASAP7_75t_SL \i45/i384  (.A(\i45/n81 ),
    .B(\i45/n571 ),
    .Y(\i45/n182 ));
 NAND2xp5_ASAP7_75t_SL \i45/i385  (.A(\i45/n58 ),
    .B(\i45/n67 ),
    .Y(\i45/n181 ));
 NAND2xp5_ASAP7_75t_SL \i45/i386  (.A(\i45/n67 ),
    .B(\i45/n89 ),
    .Y(\i45/n180 ));
 NAND2xp5_ASAP7_75t_SL \i45/i387  (.A(\i45/n84 ),
    .B(\i45/n569 ),
    .Y(\i45/n179 ));
 NAND2xp5_ASAP7_75t_SL \i45/i388  (.A(\i45/n58 ),
    .B(\i45/n95 ),
    .Y(\i45/n229 ));
 AND2x2_ASAP7_75t_SL \i45/i389  (.A(\i45/n67 ),
    .B(\i45/n91 ),
    .Y(\i45/n228 ));
 NOR3xp33_ASAP7_75t_SL \i45/i39  (.A(\i45/n488 ),
    .B(\i45/n483 ),
    .C(\i45/n11 ),
    .Y(\i45/n542 ));
 AND2x2_ASAP7_75t_SL \i45/i390  (.A(\i45/n101 ),
    .B(\i45/n89 ),
    .Y(\i45/n226 ));
 AND2x2_ASAP7_75t_SL \i45/i391  (.A(\i45/n568 ),
    .B(\i45/n571 ),
    .Y(\i45/n224 ));
 NAND2xp5_ASAP7_75t_SL \i45/i392  (.A(\i45/n571 ),
    .B(\i45/n7 ),
    .Y(\i45/n29 ));
 NAND2xp5_ASAP7_75t_SL \i45/i393  (.A(\i45/n95 ),
    .B(\i45/n569 ),
    .Y(\i45/n222 ));
 NAND2xp5_ASAP7_75t_SL \i45/i394  (.A(\i45/n107 ),
    .B(\i45/n65 ),
    .Y(\i45/n220 ));
 NAND2xp5_ASAP7_75t_SL \i45/i395  (.A(\i45/n80 ),
    .B(\i45/n89 ),
    .Y(\i45/n218 ));
 AND2x2_ASAP7_75t_SL \i45/i396  (.A(\i45/n84 ),
    .B(\i45/n75 ),
    .Y(\i45/n217 ));
 NOR2xp33_ASAP7_75t_SL \i45/i397  (.A(\i45/n82 ),
    .B(\i45/n88 ),
    .Y(\i45/n28 ));
 NOR2xp33_ASAP7_75t_SL \i45/i398  (.A(\i45/n70 ),
    .B(\i45/n82 ),
    .Y(\i45/n215 ));
 NAND2xp5_ASAP7_75t_SL \i45/i399  (.A(\i45/n83 ),
    .B(\i45/n4 ),
    .Y(\i45/n178 ));
 INVx2_ASAP7_75t_SL \i45/i4  (.A(\i45/n12 ),
    .Y(\i45/n4 ));
 NAND4xp25_ASAP7_75t_SL \i45/i40  (.A(\i45/n470 ),
    .B(\i45/n464 ),
    .C(\i45/n463 ),
    .D(\i45/n496 ),
    .Y(\i45/n541 ));
 NAND2xp5_ASAP7_75t_SL \i45/i400  (.A(\i45/n93 ),
    .B(\i45/n83 ),
    .Y(\i45/n214 ));
 NOR2xp33_ASAP7_75t_SL \i45/i401  (.A(\i45/n86 ),
    .B(\i45/n96 ),
    .Y(\i45/n177 ));
 NAND2xp5_ASAP7_75t_SL \i45/i402  (.A(\i45/n80 ),
    .B(\i45/n72 ),
    .Y(\i45/n213 ));
 NAND2xp5_ASAP7_75t_SL \i45/i403  (.A(\i45/n75 ),
    .B(\i45/n78 ),
    .Y(\i45/n176 ));
 NOR2xp33_ASAP7_75t_SL \i45/i404  (.A(\i45/n77 ),
    .B(\i45/n96 ),
    .Y(\i45/n212 ));
 AND2x2_ASAP7_75t_SL \i45/i405  (.A(\i45/n81 ),
    .B(\i45/n4 ),
    .Y(\i45/n211 ));
 NOR2xp33_ASAP7_75t_SL \i45/i406  (.A(\i45/n20 ),
    .B(\i45/n18 ),
    .Y(\i45/n175 ));
 NAND2xp5_ASAP7_75t_SL \i45/i407  (.A(\i45/n83 ),
    .B(\i45/n65 ),
    .Y(\i45/n209 ));
 NOR2xp33_ASAP7_75t_SL \i45/i408  (.A(\i45/n80 ),
    .B(\i45/n101 ),
    .Y(\i45/n174 ));
 NOR2xp33_ASAP7_75t_SL \i45/i409  (.A(\i45/n77 ),
    .B(\i45/n566 ),
    .Y(\i45/n173 ));
 NAND3xp33_ASAP7_75t_L \i45/i41  (.A(\i45/n446 ),
    .B(\i45/n464 ),
    .C(\i45/n513 ),
    .Y(\i45/n540 ));
 NAND2xp5_ASAP7_75t_SL \i45/i410  (.A(\i45/n4 ),
    .B(\i45/n101 ),
    .Y(\i45/n207 ));
 NOR2xp33_ASAP7_75t_L \i45/i411  (.A(\i45/n107 ),
    .B(\i45/n63 ),
    .Y(\i45/n206 ));
 NAND2xp5_ASAP7_75t_SL \i45/i412  (.A(\i45/n80 ),
    .B(\i45/n97 ),
    .Y(\i45/n27 ));
 NAND2xp5_ASAP7_75t_SL \i45/i413  (.A(\i45/n107 ),
    .B(\i45/n68 ),
    .Y(\i45/n204 ));
 NAND2xp5_ASAP7_75t_SL \i45/i414  (.A(\i45/n569 ),
    .B(\i45/n81 ),
    .Y(\i45/n202 ));
 NAND2xp5_ASAP7_75t_SL \i45/i415  (.A(\i45/n107 ),
    .B(\i45/n571 ),
    .Y(\i45/n200 ));
 NAND2xp5_ASAP7_75t_SL \i45/i416  (.A(\i45/n84 ),
    .B(\i45/n93 ),
    .Y(\i45/n172 ));
 NOR2xp67_ASAP7_75t_SL \i45/i417  (.A(\i45/n101 ),
    .B(\i45/n84 ),
    .Y(\i45/n198 ));
 NOR2xp33_ASAP7_75t_SL \i45/i418  (.A(\i45/n71 ),
    .B(\i45/n100 ),
    .Y(\i45/n171 ));
 NOR2x1_ASAP7_75t_SL \i45/i419  (.A(\i45/n80 ),
    .B(\i45/n570 ),
    .Y(\i45/n26 ));
 NAND3xp33_ASAP7_75t_SL \i45/i42  (.A(\i45/n450 ),
    .B(\i45/n497 ),
    .C(\i45/n484 ),
    .Y(\i45/n539 ));
 OR2x2_ASAP7_75t_SL \i45/i420  (.A(\i45/n63 ),
    .B(\i45/n83 ),
    .Y(\i45/n196 ));
 INVxp67_ASAP7_75t_SL \i45/i421  (.A(\i45/n169 ),
    .Y(\i45/n170 ));
 INVxp67_ASAP7_75t_SL \i45/i422  (.A(\i45/n164 ),
    .Y(\i45/n165 ));
 INVx1_ASAP7_75t_SL \i45/i423  (.A(\i45/n162 ),
    .Y(\i45/n163 ));
 INVxp67_ASAP7_75t_SL \i45/i424  (.A(\i45/n156 ),
    .Y(\i45/n157 ));
 INVxp67_ASAP7_75t_SL \i45/i425  (.A(\i45/n154 ),
    .Y(\i45/n155 ));
 INVxp67_ASAP7_75t_SL \i45/i426  (.A(\i45/n152 ),
    .Y(\i45/n153 ));
 INVxp67_ASAP7_75t_SL \i45/i427  (.A(\i45/n150 ),
    .Y(\i45/n151 ));
 INVxp67_ASAP7_75t_SL \i45/i428  (.A(\i45/n148 ),
    .Y(\i45/n149 ));
 INVxp67_ASAP7_75t_SL \i45/i429  (.A(\i45/n146 ),
    .Y(\i45/n147 ));
 NAND2xp5_ASAP7_75t_L \i45/i43  (.A(\i45/n576 ),
    .B(\i45/n529 ),
    .Y(\i45/n538 ));
 INVxp67_ASAP7_75t_SL \i45/i430  (.A(\i45/n138 ),
    .Y(\i45/n139 ));
 INVx1_ASAP7_75t_SL \i45/i431  (.A(\i45/n134 ),
    .Y(\i45/n135 ));
 INVx1_ASAP7_75t_SL \i45/i432  (.A(\i45/n22 ),
    .Y(\i45/n23 ));
 NAND2xp5_ASAP7_75t_SL \i45/i433  (.A(\i45/n570 ),
    .B(\i45/n91 ),
    .Y(\i45/n133 ));
 NAND2xp5_ASAP7_75t_SL \i45/i434  (.A(\i45/n63 ),
    .B(\i45/n93 ),
    .Y(\i45/n132 ));
 NAND2xp5_ASAP7_75t_SL \i45/i435  (.A(\i45/n74 ),
    .B(\i45/n91 ),
    .Y(\i45/n25 ));
 NAND2xp5_ASAP7_75t_SL \i45/i436  (.A(\i45/n94 ),
    .B(\i45/n86 ),
    .Y(\i45/n131 ));
 NAND2xp5_ASAP7_75t_SL \i45/i437  (.A(\i45/n74 ),
    .B(\i45/n93 ),
    .Y(\i45/n130 ));
 NAND2xp5_ASAP7_75t_SL \i45/i438  (.A(\i45/n93 ),
    .B(\i45/n61 ),
    .Y(\i45/n129 ));
 NAND2xp5_ASAP7_75t_SL \i45/i439  (.A(\i45/n95 ),
    .B(\i45/n75 ),
    .Y(\i45/n128 ));
 NAND2xp33_ASAP7_75t_SL \i45/i44  (.A(\i45/n494 ),
    .B(\i45/n511 ),
    .Y(\i45/n537 ));
 NOR2xp33_ASAP7_75t_SL \i45/i440  (.A(\i45/n569 ),
    .B(\i45/n4 ),
    .Y(\i45/n127 ));
 NAND2xp5_ASAP7_75t_SL \i45/i441  (.A(\i45/n87 ),
    .B(\i45/n68 ),
    .Y(\i45/n126 ));
 NAND2xp5_ASAP7_75t_SL \i45/i442  (.A(\i45/n61 ),
    .B(\i45/n89 ),
    .Y(\i45/n125 ));
 NAND2xp5_ASAP7_75t_L \i45/i443  (.A(\i45/n21 ),
    .B(\i45/n59 ),
    .Y(\i45/n124 ));
 NAND2xp33_ASAP7_75t_SL \i45/i444  (.A(\i45/n76 ),
    .B(\i45/n12 ),
    .Y(\i45/n123 ));
 NAND2xp5_ASAP7_75t_SL \i45/i445  (.A(\i45/n7 ),
    .B(\i45/n72 ),
    .Y(\i45/n122 ));
 NAND2xp5_ASAP7_75t_SL \i45/i446  (.A(\i45/n568 ),
    .B(\i45/n69 ),
    .Y(\i45/n169 ));
 NAND2xp5_ASAP7_75t_SL \i45/i447  (.A(\i45/n570 ),
    .B(\i45/n72 ),
    .Y(\i45/n121 ));
 NOR2xp33_ASAP7_75t_SL \i45/i448  (.A(\i45/n71 ),
    .B(\i45/n73 ),
    .Y(\i45/n120 ));
 NAND2xp5_ASAP7_75t_SL \i45/i449  (.A(\i45/n568 ),
    .B(\i45/n4 ),
    .Y(\i45/n168 ));
 NOR2x1_ASAP7_75t_SL \i45/i45  (.A(\i45/n510 ),
    .B(\i45/n519 ),
    .Y(\i45/n545 ));
 AND2x2_ASAP7_75t_SL \i45/i450  (.A(\i45/n7 ),
    .B(\i45/n93 ),
    .Y(\i45/n167 ));
 NOR2xp33_ASAP7_75t_SL \i45/i451  (.A(\i45/n569 ),
    .B(\i45/n97 ),
    .Y(\i45/n166 ));
 NAND2xp5_ASAP7_75t_SL \i45/i452  (.A(\i45/n101 ),
    .B(\i45/n75 ),
    .Y(\i45/n164 ));
 NOR2x1_ASAP7_75t_SL \i45/i453  (.A(\i45/n89 ),
    .B(\i45/n99 ),
    .Y(\i45/n162 ));
 NAND2xp5_ASAP7_75t_SL \i45/i454  (.A(\i45/n7 ),
    .B(\i45/n97 ),
    .Y(\i45/n161 ));
 NAND2xp5_ASAP7_75t_SL \i45/i455  (.A(\i45/n95 ),
    .B(\i45/n68 ),
    .Y(\i45/n160 ));
 NAND2xp5_ASAP7_75t_SL \i45/i456  (.A(\i45/n61 ),
    .B(\i45/n91 ),
    .Y(\i45/n119 ));
 NAND2xp5_ASAP7_75t_SL \i45/i457  (.A(\i45/n67 ),
    .B(\i45/n72 ),
    .Y(\i45/n159 ));
 AND2x2_ASAP7_75t_SL \i45/i458  (.A(\i45/n7 ),
    .B(\i45/n65 ),
    .Y(\i45/n158 ));
 NOR2xp33_ASAP7_75t_SL \i45/i459  (.A(\i45/n89 ),
    .B(\i45/n72 ),
    .Y(\i45/n118 ));
 NAND2xp33_ASAP7_75t_L \i45/i46  (.A(\i45/n499 ),
    .B(\i45/n472 ),
    .Y(\i45/n534 ));
 NAND2xp5_ASAP7_75t_SL \i45/i460  (.A(\i45/n570 ),
    .B(\i45/n569 ),
    .Y(\i45/n156 ));
 NAND2xp5_ASAP7_75t_SL \i45/i461  (.A(\i45/n65 ),
    .B(\i45/n570 ),
    .Y(\i45/n154 ));
 NOR2xp67_ASAP7_75t_SL \i45/i462  (.A(\i45/n66 ),
    .B(\i45/n103 ),
    .Y(\i45/n152 ));
 NAND2xp5_ASAP7_75t_SL \i45/i463  (.A(\i45/n61 ),
    .B(\i45/n65 ),
    .Y(\i45/n150 ));
 NAND2xp33_ASAP7_75t_L \i45/i464  (.A(\i45/n64 ),
    .B(\i45/n567 ),
    .Y(\i45/n117 ));
 NAND2xp5_ASAP7_75t_SL \i45/i465  (.A(\i45/n58 ),
    .B(\i45/n568 ),
    .Y(\i45/n148 ));
 NOR2xp67_ASAP7_75t_R \i45/i466  (.A(\i45/n59 ),
    .B(\i45/n73 ),
    .Y(\i45/n146 ));
 NAND2xp5_ASAP7_75t_SL \i45/i467  (.A(\i45/n63 ),
    .B(\i45/n97 ),
    .Y(\i45/n24 ));
 NAND2xp5_ASAP7_75t_SL \i45/i468  (.A(\i45/n63 ),
    .B(\i45/n99 ),
    .Y(\i45/n145 ));
 AND2x2_ASAP7_75t_SL \i45/i469  (.A(\i45/n568 ),
    .B(\i45/n99 ),
    .Y(\i45/n144 ));
 NAND2xp33_ASAP7_75t_SL \i45/i47  (.A(\i45/n576 ),
    .B(\i45/n478 ),
    .Y(\i45/n533 ));
 NAND2xp5_ASAP7_75t_SL \i45/i470  (.A(\i45/n4 ),
    .B(\i45/n74 ),
    .Y(\i45/n143 ));
 NAND2xp5_ASAP7_75t_L \i45/i471  (.A(\i45/n18 ),
    .B(\i45/n21 ),
    .Y(\i45/n142 ));
 NAND2xp33_ASAP7_75t_L \i45/i472  (.A(\i45/n4 ),
    .B(\i45/n95 ),
    .Y(\i45/n116 ));
 AND2x2_ASAP7_75t_SL \i45/i473  (.A(\i45/n568 ),
    .B(\i45/n75 ),
    .Y(\i45/n141 ));
 NOR2xp33_ASAP7_75t_SL \i45/i474  (.A(\i45/n76 ),
    .B(\i45/n60 ),
    .Y(\i45/n115 ));
 NOR2xp33_ASAP7_75t_SL \i45/i475  (.A(\i45/n70 ),
    .B(\i45/n62 ),
    .Y(\i45/n114 ));
 NOR2xp67_ASAP7_75t_SL \i45/i476  (.A(\i45/n69 ),
    .B(\i45/n91 ),
    .Y(\i45/n140 ));
 NAND2xp5_ASAP7_75t_SL \i45/i477  (.A(\i45/n7 ),
    .B(\i45/n99 ),
    .Y(\i45/n113 ));
 NAND2xp5_ASAP7_75t_SL \i45/i478  (.A(\i45/n74 ),
    .B(\i45/n68 ),
    .Y(\i45/n138 ));
 NAND2xp5_ASAP7_75t_SL \i45/i479  (.A(\i45/n61 ),
    .B(\i45/n4 ),
    .Y(\i45/n112 ));
 NOR2xp33_ASAP7_75t_SL \i45/i48  (.A(\i45/n477 ),
    .B(\i45/n501 ),
    .Y(\i45/n532 ));
 NAND2xp5_ASAP7_75t_SL \i45/i480  (.A(\i45/n95 ),
    .B(\i45/n99 ),
    .Y(\i45/n137 ));
 NAND2xp5_ASAP7_75t_SL \i45/i481  (.A(\i45/n74 ),
    .B(\i45/n97 ),
    .Y(\i45/n111 ));
 NAND2xp5_ASAP7_75t_SL \i45/i482  (.A(\i45/n568 ),
    .B(\i45/n93 ),
    .Y(\i45/n136 ));
 NOR2xp33_ASAP7_75t_SL \i45/i483  (.A(\i45/n108 ),
    .B(\i45/n18 ),
    .Y(\i45/n110 ));
 NOR2xp33_ASAP7_75t_SL \i45/i484  (.A(\i45/n108 ),
    .B(\i45/n71 ),
    .Y(\i45/n109 ));
 NAND2xp5_ASAP7_75t_SL \i45/i485  (.A(\i45/n74 ),
    .B(\i45/n102 ),
    .Y(\i45/n134 ));
 NAND2x1_ASAP7_75t_SL \i45/i486  (.A(\i45/n7 ),
    .B(\i45/n68 ),
    .Y(\i45/n22 ));
 INVx2_ASAP7_75t_SL \i45/i487  (.A(\i45/n568 ),
    .Y(\i45/n108 ));
 INVx1_ASAP7_75t_SL \i45/i488  (.A(\i45/n107 ),
    .Y(\i45/n106 ));
 INVx3_ASAP7_75t_SL \i45/i489  (.A(\i45/n105 ),
    .Y(\i45/n104 ));
 NAND3xp33_ASAP7_75t_SL \i45/i49  (.A(\i45/n467 ),
    .B(\i45/n475 ),
    .C(\i45/n441 ),
    .Y(\i45/n531 ));
 INVx4_ASAP7_75t_SL \i45/i490  (.A(\i45/n103 ),
    .Y(\i45/n102 ));
 INVx3_ASAP7_75t_SL \i45/i491  (.A(\i45/n101 ),
    .Y(\i45/n100 ));
 INVx2_ASAP7_75t_SL \i45/i492  (.A(\i45/n570 ),
    .Y(\i45/n98 ));
 INVx4_ASAP7_75t_SL \i45/i493  (.A(\i45/n97 ),
    .Y(\i45/n96 ));
 INVx2_ASAP7_75t_SL \i45/i494  (.A(\i45/n95 ),
    .Y(\i45/n94 ));
 INVx3_ASAP7_75t_SL \i45/i495  (.A(\i45/n93 ),
    .Y(\i45/n92 ));
 INVx2_ASAP7_75t_SL \i45/i496  (.A(\i45/n571 ),
    .Y(\i45/n90 ));
 INVx4_ASAP7_75t_SL \i45/i497  (.A(\i45/n89 ),
    .Y(\i45/n88 ));
 INVx3_ASAP7_75t_SL \i45/i498  (.A(\i45/n87 ),
    .Y(\i45/n86 ));
 INVx3_ASAP7_75t_SL \i45/i499  (.A(\i45/n85 ),
    .Y(\i45/n84 ));
 INVx2_ASAP7_75t_SL \i45/i5  (.A(\i45/n40 ),
    .Y(\i45/n5 ));
 NOR2x1_ASAP7_75t_SL \i45/i50  (.A(\i45/n422 ),
    .B(\i45/n486 ),
    .Y(\i45/n530 ));
 AND2x4_ASAP7_75t_SL \i45/i500  (.A(\i45/n52 ),
    .B(\i45/n49 ),
    .Y(\i45/n107 ));
 OR2x2_ASAP7_75t_SL \i45/i501  (.A(\i45/n39 ),
    .B(\i45/n9 ),
    .Y(\i45/n105 ));
 OR2x6_ASAP7_75t_SL \i45/i502  (.A(\i45/n44 ),
    .B(\i45/n57 ),
    .Y(\i45/n103 ));
 AND2x4_ASAP7_75t_SL \i45/i503  (.A(\i45/n38 ),
    .B(\i45/n55 ),
    .Y(\i45/n101 ));
 AND2x4_ASAP7_75t_SL \i45/i504  (.A(\i45/n43 ),
    .B(\i45/n47 ),
    .Y(\i45/n99 ));
 NAND2x1_ASAP7_75t_SL \i45/i505  (.A(\i45/n43 ),
    .B(\i45/n47 ),
    .Y(\i45/n21 ));
 AND2x4_ASAP7_75t_SL \i45/i506  (.A(\i45/n56 ),
    .B(\i45/n42 ),
    .Y(\i45/n97 ));
 AND2x4_ASAP7_75t_SL \i45/i507  (.A(\i45/n38 ),
    .B(\i45/n51 ),
    .Y(\i45/n95 ));
 AND2x4_ASAP7_75t_SL \i45/i508  (.A(\i45/n43 ),
    .B(\i45/n45 ),
    .Y(\i45/n93 ));
 AND2x4_ASAP7_75t_SL \i45/i509  (.A(\i45/n46 ),
    .B(\i45/n6 ),
    .Y(\i45/n91 ));
 NOR2xp33_ASAP7_75t_SL \i45/i51  (.A(\i45/n574 ),
    .B(\i45/n400 ),
    .Y(\i45/n529 ));
 AND2x4_ASAP7_75t_SL \i45/i510  (.A(\i45/n43 ),
    .B(\i45/n42 ),
    .Y(\i45/n89 ));
 AND2x4_ASAP7_75t_SL \i45/i511  (.A(\i45/n52 ),
    .B(\i45/n50 ),
    .Y(\i45/n87 ));
 OR2x6_ASAP7_75t_SL \i45/i512  (.A(\i45/n53 ),
    .B(\i45/n37 ),
    .Y(\i45/n85 ));
 INVx2_ASAP7_75t_SL \i45/i513  (.A(\i45/n83 ),
    .Y(\i45/n82 ));
 INVx3_ASAP7_75t_SL \i45/i514  (.A(\i45/n81 ),
    .Y(\i45/n20 ));
 INVx3_ASAP7_75t_SL \i45/i515  (.A(\i45/n80 ),
    .Y(\i45/n79 ));
 INVx3_ASAP7_75t_SL \i45/i516  (.A(\i45/n78 ),
    .Y(\i45/n77 ));
 INVx4_ASAP7_75t_SL \i45/i517  (.A(\i45/n76 ),
    .Y(\i45/n75 ));
 INVx4_ASAP7_75t_SL \i45/i518  (.A(\i45/n74 ),
    .Y(\i45/n73 ));
 INVx3_ASAP7_75t_SL \i45/i519  (.A(\i45/n72 ),
    .Y(\i45/n71 ));
 NAND2xp33_ASAP7_75t_SL \i45/i52  (.A(\i45/n499 ),
    .B(\i45/n495 ),
    .Y(\i45/n528 ));
 INVx4_ASAP7_75t_SL \i45/i520  (.A(\i45/n70 ),
    .Y(\i45/n69 ));
 INVx4_ASAP7_75t_SL \i45/i521  (.A(\i45/n68 ),
    .Y(\i45/n18 ));
 INVx4_ASAP7_75t_SL \i45/i522  (.A(\i45/n67 ),
    .Y(\i45/n66 ));
 INVx2_ASAP7_75t_SL \i45/i523  (.A(\i45/n63 ),
    .Y(\i45/n62 ));
 INVx4_ASAP7_75t_SL \i45/i524  (.A(\i45/n61 ),
    .Y(\i45/n60 ));
 INVx3_ASAP7_75t_SL \i45/i525  (.A(\i45/n59 ),
    .Y(\i45/n58 ));
 AND2x4_ASAP7_75t_SL \i45/i526  (.A(\i45/n15 ),
    .B(\i45/n52 ),
    .Y(\i45/n83 ));
 AND2x4_ASAP7_75t_SL \i45/i527  (.A(\i45/n49 ),
    .B(\i45/n55 ),
    .Y(\i45/n81 ));
 AND2x4_ASAP7_75t_SL \i45/i528  (.A(\i45/n8 ),
    .B(\i45/n50 ),
    .Y(\i45/n80 ));
 OR2x2_ASAP7_75t_SL \i45/i529  (.A(\i45/n14 ),
    .B(\i45/n54 ),
    .Y(\i45/n19 ));
 NOR2x1_ASAP7_75t_SL \i45/i53  (.A(\i45/n404 ),
    .B(\i45/n501 ),
    .Y(\i45/n527 ));
 AND2x4_ASAP7_75t_SL \i45/i530  (.A(\i45/n51 ),
    .B(\i45/n49 ),
    .Y(\i45/n78 ));
 NAND2x1p5_ASAP7_75t_SL \i45/i531  (.A(\i45/n46 ),
    .B(\i45/n56 ),
    .Y(\i45/n76 ));
 NAND2x1p5_ASAP7_75t_SL \i45/i532  (.A(\i45/n5 ),
    .B(\i45/n45 ),
    .Y(\i45/n12 ));
 AND2x4_ASAP7_75t_SL \i45/i533  (.A(\i45/n51 ),
    .B(\i45/n15 ),
    .Y(\i45/n74 ));
 AND2x4_ASAP7_75t_SL \i45/i534  (.A(\i45/n45 ),
    .B(\i45/n6 ),
    .Y(\i45/n72 ));
 OR2x4_ASAP7_75t_SL \i45/i535  (.A(\i45/n40 ),
    .B(\i45/n41 ),
    .Y(\i45/n70 ));
 AND2x4_ASAP7_75t_SL \i45/i536  (.A(\i45/n42 ),
    .B(\i45/n6 ),
    .Y(\i45/n68 ));
 AND2x4_ASAP7_75t_SL \i45/i537  (.A(\i45/n8 ),
    .B(\i45/n15 ),
    .Y(\i45/n67 ));
 AND2x4_ASAP7_75t_SL \i45/i538  (.A(\i45/n5 ),
    .B(\i45/n47 ),
    .Y(\i45/n65 ));
 NAND2x1_ASAP7_75t_SL \i45/i539  (.A(\i45/n5 ),
    .B(\i45/n47 ),
    .Y(\i45/n64 ));
 NOR2x1_ASAP7_75t_SL \i45/i54  (.A(\i45/n476 ),
    .B(\i45/n487 ),
    .Y(\i45/n526 ));
 AND2x4_ASAP7_75t_SL \i45/i540  (.A(\i45/n51 ),
    .B(\i45/n50 ),
    .Y(\i45/n63 ));
 AND2x4_ASAP7_75t_SL \i45/i541  (.A(\i45/n55 ),
    .B(\i45/n50 ),
    .Y(\i45/n61 ));
 OR2x6_ASAP7_75t_SL \i45/i542  (.A(\i45/n36 ),
    .B(\i45/n48 ),
    .Y(\i45/n59 ));
 INVx2_ASAP7_75t_SL \i45/i543  (.A(\i45/n56 ),
    .Y(\i45/n57 ));
 INVx2_ASAP7_75t_SL \i45/i544  (.A(\i45/n54 ),
    .Y(\i45/n55 ));
 NAND2xp5_ASAP7_75t_SL \i45/i545  (.A(\i45/n16 ),
    .B(\i45/n2 ),
    .Y(\i45/n48 ));
 AND2x2_ASAP7_75t_SL \i45/i546  (.A(\i45/n16 ),
    .B(\i45/n2 ),
    .Y(\i45/n56 ));
 NAND2xp5_ASAP7_75t_SL \i45/i547  (.A(\i45/n13 ),
    .B(n31[5]),
    .Y(\i45/n54 ));
 NAND2x1p5_ASAP7_75t_SL \i45/i548  (.A(n31[4]),
    .B(n31[5]),
    .Y(\i45/n53 ));
 AND2x2_ASAP7_75t_SL \i45/i549  (.A(\i45/n1 ),
    .B(\i45/n13 ),
    .Y(\i45/n52 ));
 NAND2xp5_ASAP7_75t_SL \i45/i55  (.A(\i45/n440 ),
    .B(\i45/n481 ),
    .Y(\i45/n525 ));
 AND2x2_ASAP7_75t_SL \i45/i550  (.A(n31[4]),
    .B(\i45/n1 ),
    .Y(\i45/n51 ));
 AND2x4_ASAP7_75t_SL \i45/i551  (.A(n31[7]),
    .B(\i45/n17 ),
    .Y(\i45/n50 ));
 AND2x4_ASAP7_75t_SL \i45/i552  (.A(\i45/n17 ),
    .B(\i45/n0 ),
    .Y(\i45/n49 ));
 INVx2_ASAP7_75t_SL \i45/i553  (.A(\i45/n9 ),
    .Y(\i45/n47 ));
 INVx1_ASAP7_75t_SL \i45/i554  (.A(\i45/n45 ),
    .Y(\i45/n44 ));
 INVx2_ASAP7_75t_SL \i45/i555  (.A(\i45/n41 ),
    .Y(\i45/n42 ));
 INVx2_ASAP7_75t_SL \i45/i556  (.A(\i45/n38 ),
    .Y(\i45/n37 ));
 NAND2xp5_ASAP7_75t_SL \i45/i557  (.A(\i45/n35 ),
    .B(\i45/n3 ),
    .Y(\i45/n36 ));
 AND2x2_ASAP7_75t_SL \i45/i558  (.A(n31[0]),
    .B(n31[1]),
    .Y(\i45/n46 ));
 AND2x4_ASAP7_75t_SL \i45/i559  (.A(n31[0]),
    .B(\i45/n35 ),
    .Y(\i45/n45 ));
 NOR5xp2_ASAP7_75t_SL \i45/i56  (.A(\i45/n356 ),
    .B(\i45/n33 ),
    .C(\i45/n371 ),
    .D(\i45/n573 ),
    .E(\i45/n331 ),
    .Y(\i45/n524 ));
 AND2x4_ASAP7_75t_SL \i45/i560  (.A(n31[2]),
    .B(n31[3]),
    .Y(\i45/n43 ));
 NAND2xp5_ASAP7_75t_SL \i45/i561  (.A(\i45/n3 ),
    .B(n31[1]),
    .Y(\i45/n41 ));
 OR2x2_ASAP7_75t_SL \i45/i562  (.A(\i45/n2 ),
    .B(n31[3]),
    .Y(\i45/n40 ));
 NAND2x1_ASAP7_75t_SL \i45/i563  (.A(n31[3]),
    .B(\i45/n2 ),
    .Y(\i45/n39 ));
 AND2x2_ASAP7_75t_SL \i45/i564  (.A(n31[7]),
    .B(n31[6]),
    .Y(\i45/n38 ));
 INVx1_ASAP7_75t_SL \i45/i565  (.A(n31[1]),
    .Y(\i45/n35 ));
 INVx2_ASAP7_75t_SL \i45/i566  (.A(n31[6]),
    .Y(\i45/n17 ));
 INVx2_ASAP7_75t_SL \i45/i567  (.A(n31[3]),
    .Y(\i45/n16 ));
 INVx1_ASAP7_75t_SL \i45/i568  (.A(\i45/n497 ),
    .Y(\i45/n11 ));
 AND2x2_ASAP7_75t_L \i45/i569  (.A(n31[6]),
    .B(\i45/n0 ),
    .Y(\i45/n15 ));
 NOR2x1_ASAP7_75t_SL \i45/i57  (.A(\i45/n11 ),
    .B(\i45/n488 ),
    .Y(\i45/n523 ));
 NAND2xp5_ASAP7_75t_SL \i45/i570  (.A(\i45/n0 ),
    .B(n31[6]),
    .Y(\i45/n14 ));
 INVx2_ASAP7_75t_SL \i45/i571  (.A(n31[4]),
    .Y(\i45/n13 ));
 OR2x2_ASAP7_75t_SL \i45/i572  (.A(\i45/n158 ),
    .B(\i45/n271 ),
    .Y(\i45/n10 ));
 OR2x2_ASAP7_75t_SL \i45/i573  (.A(n31[0]),
    .B(n31[1]),
    .Y(\i45/n9 ));
 INVx3_ASAP7_75t_SL \i45/i574  (.A(\i45/n569 ),
    .Y(\i45/n566 ));
 INVx2_ASAP7_75t_SL \i45/i575  (.A(\i45/n91 ),
    .Y(\i45/n567 ));
 AND2x4_ASAP7_75t_SL \i45/i576  (.A(\i45/n49 ),
    .B(\i45/n8 ),
    .Y(\i45/n568 ));
 AND2x4_ASAP7_75t_SL \i45/i577  (.A(\i45/n46 ),
    .B(\i45/n5 ),
    .Y(\i45/n569 ));
 AND2x4_ASAP7_75t_SL \i45/i578  (.A(\i45/n38 ),
    .B(\i45/n52 ),
    .Y(\i45/n570 ));
 AND2x4_ASAP7_75t_SL \i45/i579  (.A(\i45/n46 ),
    .B(\i45/n43 ),
    .Y(\i45/n571 ));
 NAND2xp5_ASAP7_75t_SL \i45/i58  (.A(\i45/n485 ),
    .B(\i45/n465 ),
    .Y(\i45/n536 ));
 NAND2xp5_ASAP7_75t_SL \i45/i580  (.A(\i45/n297 ),
    .B(\i45/n572 ),
    .Y(\i45/n573 ));
 AOI22xp5_ASAP7_75t_SL \i45/i581  (.A1(\i45/n568 ),
    .A2(\i45/n569 ),
    .B1(\i45/n570 ),
    .B2(\i45/n571 ),
    .Y(\i45/n572 ));
 NAND3xp33_ASAP7_75t_SL \i45/i582  (.A(\i45/n365 ),
    .B(\i45/n395 ),
    .C(\i45/n572 ),
    .Y(\i45/n574 ));
 AND4x1_ASAP7_75t_SL \i45/i583  (.A(\i45/n355 ),
    .B(\i45/n402 ),
    .C(\i45/n416 ),
    .D(\i45/n325 ),
    .Y(\i45/n575 ));
 AND4x1_ASAP7_75t_SL \i45/i584  (.A(\i45/n343 ),
    .B(\i45/n405 ),
    .C(\i45/n370 ),
    .D(\i45/n355 ),
    .Y(\i45/n576 ));
 AND2x2_ASAP7_75t_SL \i45/i585  (.A(\i45/n577 ),
    .B(\i45/n498 ),
    .Y(\i45/n578 ));
 AOI21xp33_ASAP7_75t_SL \i45/i586  (.A1(\i45/n58 ),
    .A2(\i45/n87 ),
    .B(\i45/n144 ),
    .Y(\i45/n577 ));
 NAND3xp33_ASAP7_75t_SL \i45/i587  (.A(\i45/n579 ),
    .B(\i45/n317 ),
    .C(\i45/n393 ),
    .Y(\i45/n580 ));
 AO21x1_ASAP7_75t_SL \i45/i588  (.A1(\i45/n82 ),
    .A2(\i45/n66 ),
    .B(\i45/n566 ),
    .Y(\i45/n579 ));
 NOR3xp33_ASAP7_75t_SL \i45/i589  (.A(\i45/n581 ),
    .B(\i45/n391 ),
    .C(\i45/n259 ),
    .Y(\i45/n582 ));
 NOR2x1_ASAP7_75t_SL \i45/i59  (.A(\i45/n502 ),
    .B(\i45/n487 ),
    .Y(\i45/n522 ));
 OAI21xp5_ASAP7_75t_SL \i45/i590  (.A1(\i45/n85 ),
    .A2(\i45/n21 ),
    .B(\i45/n143 ),
    .Y(\i45/n581 ));
 INVx1_ASAP7_75t_SL \i45/i6  (.A(\i45/n39 ),
    .Y(\i45/n6 ));
 NOR2x1_ASAP7_75t_SL \i45/i60  (.A(\i45/n421 ),
    .B(\i45/n486 ),
    .Y(\i45/n535 ));
 INVxp67_ASAP7_75t_SL \i45/i61  (.A(\i45/n520 ),
    .Y(\i45/n521 ));
 INVxp67_ASAP7_75t_SL \i45/i62  (.A(\i45/n516 ),
    .Y(\i45/n517 ));
 AND5x1_ASAP7_75t_SL \i45/i63  (.A(\i45/n435 ),
    .B(\i45/n416 ),
    .C(\i45/n427 ),
    .D(\i45/n341 ),
    .E(\i45/n310 ),
    .Y(\i45/n515 ));
 NOR3xp33_ASAP7_75t_SL \i45/i64  (.A(\i45/n447 ),
    .B(\i45/n426 ),
    .C(\i45/n406 ),
    .Y(\i45/n514 ));
 NOR3xp33_ASAP7_75t_SL \i45/i65  (.A(\i45/n473 ),
    .B(\i45/n407 ),
    .C(\i45/n353 ),
    .Y(\i45/n513 ));
 AND5x1_ASAP7_75t_SL \i45/i66  (.A(\i45/n396 ),
    .B(\i45/n410 ),
    .C(\i45/n389 ),
    .D(\i45/n399 ),
    .E(\i45/n319 ),
    .Y(\i45/n512 ));
 NOR2xp33_ASAP7_75t_SL \i45/i67  (.A(\i45/n474 ),
    .B(\i45/n479 ),
    .Y(\i45/n511 ));
 NAND4xp25_ASAP7_75t_SL \i45/i68  (.A(\i45/n456 ),
    .B(\i45/n464 ),
    .C(\i45/n469 ),
    .D(\i45/n452 ),
    .Y(\i45/n510 ));
 NAND5xp2_ASAP7_75t_SL \i45/i69  (.A(\i45/n434 ),
    .B(\i45/n277 ),
    .C(\i45/n387 ),
    .D(\i45/n262 ),
    .E(\i45/n366 ),
    .Y(\i45/n509 ));
 INVx2_ASAP7_75t_SL \i45/i7  (.A(\i45/n19 ),
    .Y(\i45/n7 ));
 NOR4xp25_ASAP7_75t_SL \i45/i70  (.A(\i45/n424 ),
    .B(\i45/n33 ),
    .C(\i45/n372 ),
    .D(\i45/n345 ),
    .Y(\i45/n508 ));
 NAND4xp25_ASAP7_75t_SL \i45/i71  (.A(\i45/n444 ),
    .B(\i45/n458 ),
    .C(\i45/n461 ),
    .D(\i45/n463 ),
    .Y(\i45/n507 ));
 NAND4xp25_ASAP7_75t_SL \i45/i72  (.A(\i45/n471 ),
    .B(\i45/n469 ),
    .C(\i45/n235 ),
    .D(\i45/n309 ),
    .Y(\i45/n506 ));
 NAND3xp33_ASAP7_75t_SL \i45/i73  (.A(\i45/n463 ),
    .B(\i45/n433 ),
    .C(\i45/n24 ),
    .Y(\i45/n520 ));
 NAND4xp75_ASAP7_75t_SL \i45/i74  (.A(\i45/n362 ),
    .B(\i45/n330 ),
    .C(\i45/n420 ),
    .D(\i45/n29 ),
    .Y(\i45/n519 ));
 NAND2xp33_ASAP7_75t_L \i45/i75  (.A(\i45/n443 ),
    .B(\i45/n503 ),
    .Y(\i45/n505 ));
 AND2x2_ASAP7_75t_SL \i45/i76  (.A(\i45/n446 ),
    .B(\i45/n493 ),
    .Y(\i45/n518 ));
 NAND2xp5_ASAP7_75t_SL \i45/i77  (.A(\i45/n500 ),
    .B(\i45/n457 ),
    .Y(\i45/n516 ));
 INVxp67_ASAP7_75t_SL \i45/i78  (.A(\i45/n503 ),
    .Y(\i45/n504 ));
 NOR5xp2_ASAP7_75t_SL \i45/i79  (.A(\i45/n382 ),
    .B(\i45/n352 ),
    .C(\i45/n269 ),
    .D(\i45/n224 ),
    .E(\i45/n114 ),
    .Y(\i45/n496 ));
 INVx2_ASAP7_75t_SL \i45/i8  (.A(\i45/n53 ),
    .Y(\i45/n8 ));
 NOR3xp33_ASAP7_75t_SL \i45/i80  (.A(\i45/n468 ),
    .B(\i45/n377 ),
    .C(\i45/n369 ),
    .Y(\i45/n495 ));
 NOR2xp33_ASAP7_75t_SL \i45/i81  (.A(\i45/n423 ),
    .B(\i45/n445 ),
    .Y(\i45/n494 ));
 NOR2xp33_ASAP7_75t_SL \i45/i82  (.A(\i45/n466 ),
    .B(\i45/n412 ),
    .Y(\i45/n493 ));
 NOR2x1_ASAP7_75t_SL \i45/i83  (.A(\i45/n428 ),
    .B(\i45/n397 ),
    .Y(\i45/n503 ));
 NAND2xp5_ASAP7_75t_L \i45/i84  (.A(\i45/n465 ),
    .B(\i45/n432 ),
    .Y(\i45/n492 ));
 NAND2xp5_ASAP7_75t_SL \i45/i85  (.A(\i45/n455 ),
    .B(\i45/n411 ),
    .Y(\i45/n491 ));
 NAND3xp33_ASAP7_75t_SL \i45/i86  (.A(\i45/n416 ),
    .B(\i45/n347 ),
    .C(\i45/n325 ),
    .Y(\i45/n502 ));
 NOR3xp33_ASAP7_75t_SL \i45/i87  (.A(\i45/n436 ),
    .B(\i45/n10 ),
    .C(\i45/n327 ),
    .Y(\i45/n490 ));
 NAND2xp5_ASAP7_75t_SL \i45/i88  (.A(\i45/n27 ),
    .B(\i45/n444 ),
    .Y(\i45/n501 ));
 OR3x1_ASAP7_75t_SL \i45/i89  (.A(\i45/n356 ),
    .B(\i45/n371 ),
    .C(\i45/n573 ),
    .Y(\i45/n489 ));
 NOR2x2_ASAP7_75t_SL \i45/i9  (.A(\i45/n561 ),
    .B(\i45/n560 ),
    .Y(n30[4]));
 NOR2x1_ASAP7_75t_SL \i45/i90  (.A(\i45/n369 ),
    .B(\i45/n468 ),
    .Y(\i45/n500 ));
 NOR2xp33_ASAP7_75t_SL \i45/i91  (.A(\i45/n425 ),
    .B(\i45/n409 ),
    .Y(\i45/n499 ));
 NOR2xp33_ASAP7_75t_SL \i45/i92  (.A(\i45/n357 ),
    .B(\i45/n454 ),
    .Y(\i45/n498 ));
 NOR3x1_ASAP7_75t_SL \i45/i93  (.A(\i45/n364 ),
    .B(\i45/n240 ),
    .C(\i45/n417 ),
    .Y(\i45/n497 ));
 NOR3xp33_ASAP7_75t_SL \i45/i94  (.A(\i45/n373 ),
    .B(\i45/n276 ),
    .C(\i45/n360 ),
    .Y(\i45/n485 ));
 NOR2xp33_ASAP7_75t_SL \i45/i95  (.A(\i45/n580 ),
    .B(\i45/n439 ),
    .Y(\i45/n484 ));
 NAND3xp33_ASAP7_75t_SL \i45/i96  (.A(\i45/n355 ),
    .B(\i45/n430 ),
    .C(\i45/n370 ),
    .Y(\i45/n483 ));
 NAND4xp25_ASAP7_75t_SL \i45/i97  (.A(\i45/n336 ),
    .B(\i45/n351 ),
    .C(\i45/n383 ),
    .D(\i45/n346 ),
    .Y(\i45/n482 ));
 NAND2x1_ASAP7_75t_SL \i45/i98  (.A(\i45/n453 ),
    .B(\i45/n467 ),
    .Y(\i45/n488 ));
 NOR5xp2_ASAP7_75t_SL \i45/i99  (.A(\i45/n462 ),
    .B(\i45/n375 ),
    .C(\i45/n157 ),
    .D(\i45/n293 ),
    .E(\i45/n203 ),
    .Y(\i45/n481 ));
 XOR2xp5_ASAP7_75t_SL i450 (.A(n621),
    .B(n620),
    .Y(n1022));
 AOI22xp5_ASAP7_75t_SL i451 (.A1(n860),
    .A2(n1177),
    .B1(n861),
    .B2(n769),
    .Y(n1021));
 OAI22xp5_ASAP7_75t_SL i452 (.A1(n859),
    .A2(n815),
    .B1(n814),
    .B2(n858),
    .Y(n1020));
 XNOR2xp5_ASAP7_75t_SL i453 (.A(n614),
    .B(n775),
    .Y(n1019));
 XNOR2xp5_ASAP7_75t_SL i454 (.A(n613),
    .B(n770),
    .Y(n1018));
 AOI22xp5_ASAP7_75t_SL i455 (.A1(n854),
    .A2(n1153),
    .B1(n219),
    .B2(n227),
    .Y(n1017));
 OAI22xp5_ASAP7_75t_SL i456 (.A1(n853),
    .A2(n483),
    .B1(n852),
    .B2(n482),
    .Y(n1016));
 OAI22xp5_ASAP7_75t_SL i457 (.A1(n851),
    .A2(n782),
    .B1(n850),
    .B2(n781),
    .Y(n1015));
 OAI22xp5_ASAP7_75t_SL i458 (.A1(n849),
    .A2(n510),
    .B1(n848),
    .B2(n511),
    .Y(n1014));
 AOI22xp5_ASAP7_75t_SL i459 (.A1(n846),
    .A2(n223),
    .B1(n847),
    .B2(n778),
    .Y(n1013));
 INVx2_ASAP7_75t_SL \i46/i0  (.A(n29[7]),
    .Y(\i46/n0 ));
 INVx2_ASAP7_75t_SL \i46/i1  (.A(n29[5]),
    .Y(\i46/n1 ));
 INVx2_ASAP7_75t_SL \i46/i10  (.A(\i46/n440 ),
    .Y(\i46/n10 ));
 NAND3xp33_ASAP7_75t_SL \i46/i100  (.A(\i46/n496 ),
    .B(\i46/n306 ),
    .C(\i46/n572 ),
    .Y(\i46/n355 ));
 NAND4xp25_ASAP7_75t_SL \i46/i101  (.A(\i46/n228 ),
    .B(\i46/n574 ),
    .C(\i46/n264 ),
    .D(\i46/n235 ),
    .Y(\i46/n354 ));
 NAND2x1_ASAP7_75t_SL \i46/i102  (.A(\i46/n326 ),
    .B(\i46/n340 ),
    .Y(\i46/n360 ));
 NOR5xp2_ASAP7_75t_SL \i46/i103  (.A(\i46/n335 ),
    .B(\i46/n257 ),
    .C(\i46/n112 ),
    .D(\i46/n195 ),
    .E(\i46/n144 ),
    .Y(\i46/n353 ));
 NAND3xp33_ASAP7_75t_SL \i46/i104  (.A(\i46/n292 ),
    .B(\i46/n313 ),
    .C(\i46/n478 ),
    .Y(\i46/n352 ));
 NAND2xp33_ASAP7_75t_SL \i46/i105  (.A(\i46/n573 ),
    .B(\i46/n332 ),
    .Y(\i46/n351 ));
 NOR5xp2_ASAP7_75t_SL \i46/i106  (.A(\i46/n277 ),
    .B(\i46/n242 ),
    .C(\i46/n262 ),
    .D(\i46/n215 ),
    .E(\i46/n180 ),
    .Y(\i46/n350 ));
 NAND5xp2_ASAP7_75t_SL \i46/i107  (.A(\i46/n495 ),
    .B(\i46/n291 ),
    .C(\i46/n479 ),
    .D(\i46/n446 ),
    .E(\i46/n538 ),
    .Y(\i46/n349 ));
 NAND3xp33_ASAP7_75t_L \i46/i108  (.A(\i46/n220 ),
    .B(\i46/n247 ),
    .C(\i46/n316 ),
    .Y(\i46/n348 ));
 NOR5xp2_ASAP7_75t_SL \i46/i109  (.A(\i46/n218 ),
    .B(\i46/n230 ),
    .C(\i46/n212 ),
    .D(\i46/n100 ),
    .E(\i46/n84 ),
    .Y(\i46/n347 ));
 NOR2x2_ASAP7_75t_SL \i46/i11  (.A(\i46/n435 ),
    .B(\i46/n434 ),
    .Y(n28[4]));
 NAND5xp2_ASAP7_75t_SL \i46/i110  (.A(\i46/n25 ),
    .B(\i46/n525 ),
    .C(\i46/n479 ),
    .D(\i46/n503 ),
    .E(\i46/n159 ),
    .Y(\i46/n346 ));
 NOR5xp2_ASAP7_75t_SL \i46/i111  (.A(\i46/n188 ),
    .B(\i46/n526 ),
    .C(\i46/n179 ),
    .D(\i46/n156 ),
    .E(\i46/n154 ),
    .Y(\i46/n345 ));
 NOR2xp33_ASAP7_75t_SL \i46/i112  (.A(\i46/n307 ),
    .B(\i46/n339 ),
    .Y(\i46/n344 ));
 NOR2xp33_ASAP7_75t_SL \i46/i113  (.A(\i46/n295 ),
    .B(\i46/n324 ),
    .Y(\i46/n343 ));
 NAND3x2_ASAP7_75t_SL \i46/i114  (.B(\i46/n322 ),
    .C(\i46/n291 ),
    .Y(\i46/n359 ),
    .A(\i46/n487 ));
 NAND3x1_ASAP7_75t_SL \i46/i115  (.A(\i46/n286 ),
    .B(\i46/n266 ),
    .C(\i46/n237 ),
    .Y(\i46/n358 ));
 AOI21xp5_ASAP7_75t_L \i46/i116  (.A1(\i46/n62 ),
    .A2(\i46/n564 ),
    .B(\i46/n138 ),
    .Y(\i46/n335 ));
 NOR2xp33_ASAP7_75t_SL \i46/i117  (.A(\i46/n522 ),
    .B(\i46/n277 ),
    .Y(\i46/n334 ));
 NAND2xp5_ASAP7_75t_SL \i46/i118  (.A(\i46/n265 ),
    .B(\i46/n294 ),
    .Y(\i46/n333 ));
 NOR2xp33_ASAP7_75t_SL \i46/i119  (.A(\i46/n293 ),
    .B(\i46/n26 ),
    .Y(\i46/n332 ));
 NOR2x2_ASAP7_75t_SL \i46/i12  (.A(\i46/n430 ),
    .B(\i46/n436 ),
    .Y(n28[3]));
 NOR2xp33_ASAP7_75t_SL \i46/i120  (.A(\i46/n272 ),
    .B(\i46/n282 ),
    .Y(\i46/n331 ));
 NOR2xp67_ASAP7_75t_SL \i46/i121  (.A(\i46/n146 ),
    .B(\i46/n279 ),
    .Y(\i46/n330 ));
 NOR2xp33_ASAP7_75t_SL \i46/i122  (.A(\i46/n22 ),
    .B(\i46/n277 ),
    .Y(\i46/n329 ));
 NOR4xp25_ASAP7_75t_SL \i46/i123  (.A(\i46/n251 ),
    .B(\i46/n458 ),
    .C(\i46/n22 ),
    .D(\i46/n531 ),
    .Y(\i46/n328 ));
 NAND2xp5_ASAP7_75t_SL \i46/i124  (.A(\i46/n209 ),
    .B(\i46/n258 ),
    .Y(\i46/n327 ));
 NOR4xp25_ASAP7_75t_SL \i46/i125  (.A(\i46/n97 ),
    .B(\i46/n201 ),
    .C(\i46/n181 ),
    .D(\i46/n190 ),
    .Y(\i46/n326 ));
 NOR3xp33_ASAP7_75t_SL \i46/i126  (.A(\i46/n206 ),
    .B(\i46/n175 ),
    .C(\i46/n205 ),
    .Y(\i46/n325 ));
 NAND2xp33_ASAP7_75t_SL \i46/i127  (.A(\i46/n246 ),
    .B(\i46/n23 ),
    .Y(\i46/n324 ));
 NOR2xp33_ASAP7_75t_SL \i46/i128  (.A(\i46/n522 ),
    .B(\i46/n241 ),
    .Y(\i46/n323 ));
 NOR2x1p5_ASAP7_75t_SL \i46/i129  (.A(\i46/n226 ),
    .B(\i46/n556 ),
    .Y(\i46/n322 ));
 AND5x2_ASAP7_75t_SL \i46/i13  (.A(\i46/n428 ),
    .B(\i46/n419 ),
    .C(\i46/n421 ),
    .D(\i46/n406 ),
    .E(\i46/n398 ),
    .Y(n28[6]));
 NAND2xp33_ASAP7_75t_SL \i46/i130  (.A(\i46/n292 ),
    .B(\i46/n275 ),
    .Y(\i46/n321 ));
 NAND3xp33_ASAP7_75t_SL \i46/i131  (.A(\i46/n24 ),
    .B(\i46/n174 ),
    .C(\i46/n447 ),
    .Y(\i46/n320 ));
 NOR3xp33_ASAP7_75t_SL \i46/i132  (.A(\i46/n457 ),
    .B(\i46/n185 ),
    .C(\i46/n164 ),
    .Y(\i46/n342 ));
 NAND2xp5_ASAP7_75t_SL \i46/i133  (.A(\i46/n250 ),
    .B(\i46/n490 ),
    .Y(\i46/n341 ));
 NOR2x1_ASAP7_75t_SL \i46/i134  (.A(\i46/n225 ),
    .B(\i46/n244 ),
    .Y(\i46/n340 ));
 NAND2xp67_ASAP7_75t_SL \i46/i135  (.A(\i46/n479 ),
    .B(\i46/n252 ),
    .Y(\i46/n339 ));
 NOR2x1_ASAP7_75t_SL \i46/i136  (.A(\i46/n227 ),
    .B(\i46/n280 ),
    .Y(\i46/n338 ));
 NOR2x1_ASAP7_75t_SL \i46/i137  (.A(\i46/n458 ),
    .B(\i46/n522 ),
    .Y(\i46/n337 ));
 NOR3x1_ASAP7_75t_SL \i46/i138  (.A(\i46/n179 ),
    .B(\i46/n173 ),
    .C(\i46/n153 ),
    .Y(\i46/n336 ));
 INVx1_ASAP7_75t_SL \i46/i139  (.A(\i46/n27 ),
    .Y(\i46/n317 ));
 AND3x4_ASAP7_75t_SL \i46/i14  (.A(\i46/n428 ),
    .B(\i46/n437 ),
    .C(\i46/n416 ),
    .Y(n28[1]));
 NOR4xp25_ASAP7_75t_SL \i46/i140  (.A(\i46/n167 ),
    .B(\i46/n192 ),
    .C(\i46/n184 ),
    .D(\i46/n162 ),
    .Y(\i46/n316 ));
 NAND2xp33_ASAP7_75t_L \i46/i141  (.A(\i46/n238 ),
    .B(\i46/n260 ),
    .Y(\i46/n315 ));
 NAND5xp2_ASAP7_75t_SL \i46/i142  (.A(\i46/n542 ),
    .B(\i46/n200 ),
    .C(\i46/n211 ),
    .D(\i46/n545 ),
    .E(\i46/n484 ),
    .Y(\i46/n314 ));
 NOR4xp25_ASAP7_75t_SL \i46/i143  (.A(\i46/n268 ),
    .B(\i46/n124 ),
    .C(\i46/n459 ),
    .D(\i46/n143 ),
    .Y(\i46/n313 ));
 OAI221xp5_ASAP7_75t_SL \i46/i144  (.A1(\i46/n101 ),
    .A2(\i46/n79 ),
    .B1(\i46/n101 ),
    .B2(\i46/n18 ),
    .C(\i46/n246 ),
    .Y(\i46/n312 ));
 NOR2xp33_ASAP7_75t_SL \i46/i145  (.A(\i46/n231 ),
    .B(\i46/n449 ),
    .Y(\i46/n311 ));
 AOI211xp5_ASAP7_75t_SL \i46/i146  (.A1(\i46/n141 ),
    .A2(\i46/n63 ),
    .B(\i46/n217 ),
    .C(\i46/n157 ),
    .Y(\i46/n310 ));
 OA21x2_ASAP7_75t_SL \i46/i147  (.A1(\i46/n47 ),
    .A2(\i46/n62 ),
    .B(\i46/n525 ),
    .Y(\i46/n309 ));
 NOR4xp25_ASAP7_75t_SL \i46/i148  (.A(\i46/n454 ),
    .B(\i46/n149 ),
    .C(\i46/n455 ),
    .D(\i46/n153 ),
    .Y(\i46/n308 ));
 NAND5xp2_ASAP7_75t_SL \i46/i149  (.A(\i46/n125 ),
    .B(\i46/n546 ),
    .C(\i46/n133 ),
    .D(\i46/n569 ),
    .E(\i46/n83 ),
    .Y(\i46/n307 ));
 NOR2x1p5_ASAP7_75t_SL \i46/i15  (.A(\i46/n438 ),
    .B(\i46/n429 ),
    .Y(n28[5]));
 NOR3xp33_ASAP7_75t_SL \i46/i150  (.A(\i46/n245 ),
    .B(\i46/n460 ),
    .C(\i46/n82 ),
    .Y(\i46/n306 ));
 NAND2xp5_ASAP7_75t_SL \i46/i151  (.A(\i46/n229 ),
    .B(\i46/n25 ),
    .Y(\i46/n305 ));
 NAND5xp2_ASAP7_75t_SL \i46/i152  (.A(\i46/n537 ),
    .B(\i46/n92 ),
    .C(\i46/n170 ),
    .D(\i46/n161 ),
    .E(\i46/n544 ),
    .Y(\i46/n304 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i46/i153  (.A1(\i46/n67 ),
    .A2(\i46/n85 ),
    .B(\i46/n69 ),
    .C(\i46/n222 ),
    .Y(\i46/n303 ));
 NOR4xp25_ASAP7_75t_SL \i46/i154  (.A(\i46/n271 ),
    .B(\i46/n176 ),
    .C(\i46/n127 ),
    .D(\i46/n102 ),
    .Y(\i46/n302 ));
 NAND4xp25_ASAP7_75t_SL \i46/i155  (.A(\i46/n256 ),
    .B(\i46/n536 ),
    .C(\i46/n98 ),
    .D(\i46/n151 ),
    .Y(\i46/n301 ));
 NAND5xp2_ASAP7_75t_SL \i46/i156  (.A(\i46/n142 ),
    .B(\i46/n126 ),
    .C(\i46/n194 ),
    .D(\i46/n473 ),
    .E(\i46/n90 ),
    .Y(\i46/n300 ));
 NAND2xp5_ASAP7_75t_SL \i46/i157  (.A(\i46/n463 ),
    .B(\i46/n249 ),
    .Y(\i46/n299 ));
 NAND2xp5_ASAP7_75t_SL \i46/i158  (.A(\i46/n487 ),
    .B(\i46/n291 ),
    .Y(\i46/n298 ));
 NOR2xp33_ASAP7_75t_L \i46/i159  (.A(\i46/n270 ),
    .B(\i46/n282 ),
    .Y(\i46/n319 ));
 AND2x2_ASAP7_75t_SL \i46/i16  (.A(\i46/n439 ),
    .B(\i46/n422 ),
    .Y(n28[0]));
 NAND2xp5_ASAP7_75t_SL \i46/i160  (.A(\i46/n478 ),
    .B(\i46/n292 ),
    .Y(\i46/n297 ));
 NOR2x1_ASAP7_75t_SL \i46/i161  (.A(\i46/n232 ),
    .B(\i46/n274 ),
    .Y(\i46/n318 ));
 NAND3x1_ASAP7_75t_SL \i46/i162  (.A(\i46/n214 ),
    .B(\i46/n481 ),
    .C(\i46/n128 ),
    .Y(\i46/n27 ));
 INVxp67_ASAP7_75t_SL \i46/i163  (.A(\i46/n295 ),
    .Y(\i46/n296 ));
 INVxp67_ASAP7_75t_SL \i46/i164  (.A(\i46/n12 ),
    .Y(\i46/n294 ));
 INVxp67_ASAP7_75t_SL \i46/i165  (.A(\i46/n289 ),
    .Y(\i46/n290 ));
 INVxp67_ASAP7_75t_SL \i46/i166  (.A(\i46/n287 ),
    .Y(\i46/n288 ));
 INVx2_ASAP7_75t_SL \i46/i167  (.A(\i46/n285 ),
    .Y(\i46/n286 ));
 INVxp67_ASAP7_75t_SL \i46/i168  (.A(\i46/n283 ),
    .Y(\i46/n284 ));
 INVxp67_ASAP7_75t_SL \i46/i169  (.A(\i46/n280 ),
    .Y(\i46/n281 ));
 NOR3xp33_ASAP7_75t_SL \i46/i17  (.A(\i46/n411 ),
    .B(\i46/n407 ),
    .C(\i46/n414 ),
    .Y(\i46/n439 ));
 INVxp67_ASAP7_75t_SL \i46/i170  (.A(\i46/n524 ),
    .Y(\i46/n278 ));
 INVx1_ASAP7_75t_SL \i46/i171  (.A(\i46/n275 ),
    .Y(\i46/n276 ));
 NAND2x1_ASAP7_75t_SL \i46/i172  (.A(\i46/n470 ),
    .B(\i46/n183 ),
    .Y(\i46/n274 ));
 NOR2xp33_ASAP7_75t_SL \i46/i173  (.A(\i46/n444 ),
    .B(\i46/n206 ),
    .Y(\i46/n273 ));
 NAND2xp33_ASAP7_75t_SL \i46/i174  (.A(\i46/n174 ),
    .B(\i46/n479 ),
    .Y(\i46/n272 ));
 OAI21xp33_ASAP7_75t_SL \i46/i175  (.A1(\i46/n45 ),
    .A2(\i46/n562 ),
    .B(\i46/n491 ),
    .Y(\i46/n271 ));
 NAND2xp5_ASAP7_75t_SL \i46/i176  (.A(\i46/n152 ),
    .B(\i46/n174 ),
    .Y(\i46/n270 ));
 AOI211xp5_ASAP7_75t_SL \i46/i177  (.A1(\i46/n77 ),
    .A2(\i46/n31 ),
    .B(\i46/n482 ),
    .C(\i46/n107 ),
    .Y(\i46/n269 ));
 AOI31xp33_ASAP7_75t_SL \i46/i178  (.A1(\i46/n45 ),
    .A2(\i46/n19 ),
    .A3(\i46/n53 ),
    .B(\i46/n485 ),
    .Y(\i46/n268 ));
 NOR3xp33_ASAP7_75t_SL \i46/i179  (.A(\i46/n175 ),
    .B(\i46/n117 ),
    .C(\i46/n105 ),
    .Y(\i46/n267 ));
 NOR2x2_ASAP7_75t_SL \i46/i18  (.A(\i46/n431 ),
    .B(\i46/n432 ),
    .Y(n28[2]));
 NOR3xp33_ASAP7_75t_SL \i46/i180  (.A(\i46/n483 ),
    .B(\i46/n113 ),
    .C(\i46/n444 ),
    .Y(\i46/n266 ));
 AOI221xp5_ASAP7_75t_SL \i46/i181  (.A1(\i46/n67 ),
    .A2(\i46/n80 ),
    .B1(\i46/n523 ),
    .B2(\i46/n55 ),
    .C(\i46/n163 ),
    .Y(\i46/n265 ));
 OAI31xp33_ASAP7_75t_R \i46/i182  (.A1(\i46/n63 ),
    .A2(\i46/n65 ),
    .A3(\i46/n67 ),
    .B(\i46/n61 ),
    .Y(\i46/n264 ));
 AOI21xp5_ASAP7_75t_SL \i46/i183  (.A1(\i46/n138 ),
    .A2(\i46/n53 ),
    .B(\i46/n575 ),
    .Y(\i46/n295 ));
 AOI21xp5_ASAP7_75t_R \i46/i184  (.A1(\i46/n53 ),
    .A2(\i46/n471 ),
    .B(\i46/n76 ),
    .Y(\i46/n263 ));
 OAI221xp5_ASAP7_75t_SL \i46/i185  (.A1(\i46/n461 ),
    .A2(\i46/n79 ),
    .B1(\i46/n468 ),
    .B2(\i46/n539 ),
    .C(\i46/n565 ),
    .Y(\i46/n262 ));
 AOI21xp33_ASAP7_75t_SL \i46/i186  (.A1(\i46/n471 ),
    .A2(\i46/n41 ),
    .B(\i46/n66 ),
    .Y(\i46/n261 ));
 NOR3xp33_ASAP7_75t_SL \i46/i187  (.A(\i46/n189 ),
    .B(\i46/n483 ),
    .C(\i46/n122 ),
    .Y(\i46/n260 ));
 NAND3xp33_ASAP7_75t_SL \i46/i188  (.A(\i46/n499 ),
    .B(\i46/n501 ),
    .C(\i46/n145 ),
    .Y(\i46/n259 ));
 AOI22xp5_ASAP7_75t_SL \i46/i189  (.A1(\i46/n49 ),
    .A2(\i46/n134 ),
    .B1(\i46/n55 ),
    .B2(\i46/n440 ),
    .Y(\i46/n258 ));
 NAND4xp75_ASAP7_75t_SL \i46/i19  (.A(\i46/n397 ),
    .B(\i46/n417 ),
    .C(\i46/n395 ),
    .D(\i46/n577 ),
    .Y(\i46/n438 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i46/i190  (.A1(\i46/n76 ),
    .A2(\i46/n43 ),
    .B(\i46/n60 ),
    .C(\i46/n474 ),
    .Y(\i46/n257 ));
 OAI21xp5_ASAP7_75t_SL \i46/i191  (.A1(\i46/n52 ),
    .A2(\i46/n139 ),
    .B(\i46/n63 ),
    .Y(\i46/n256 ));
 NAND4xp25_ASAP7_75t_SL \i46/i192  (.A(\i46/n155 ),
    .B(\i46/n151 ),
    .C(\i46/n513 ),
    .D(\i46/n129 ),
    .Y(\i46/n255 ));
 NAND2xp33_ASAP7_75t_SL \i46/i193  (.A(\i46/n196 ),
    .B(\i46/n121 ),
    .Y(\i46/n254 ));
 OAI211xp5_ASAP7_75t_SL \i46/i194  (.A1(\i46/n59 ),
    .A2(\i46/n66 ),
    .B(\i46/n570 ),
    .C(\i46/n543 ),
    .Y(\i46/n293 ));
 NOR2xp67_ASAP7_75t_SL \i46/i195  (.A(\i46/n527 ),
    .B(\i46/n212 ),
    .Y(\i46/n292 ));
 AOI21x1_ASAP7_75t_SL \i46/i196  (.A1(\i46/n440 ),
    .A2(\i46/n52 ),
    .B(\i46/n217 ),
    .Y(\i46/n291 ));
 NAND2xp5_ASAP7_75t_SL \i46/i197  (.A(\i46/n541 ),
    .B(\i46/n563 ),
    .Y(\i46/n26 ));
 NOR2xp33_ASAP7_75t_SL \i46/i198  (.A(\i46/n198 ),
    .B(\i46/n454 ),
    .Y(\i46/n289 ));
 OAI211xp5_ASAP7_75t_SL \i46/i199  (.A1(\i46/n53 ),
    .A2(\i46/n66 ),
    .B(\i46/n491 ),
    .C(\i46/n512 ),
    .Y(\i46/n287 ));
 INVxp67_ASAP7_75t_SL \i46/i2  (.A(n29[4]),
    .Y(\i46/n2 ));
 NOR3xp33_ASAP7_75t_SL \i46/i20  (.A(\i46/n415 ),
    .B(\i46/n380 ),
    .C(\i46/n425 ),
    .Y(\i46/n437 ));
 OR2x2_ASAP7_75t_SL \i46/i200  (.A(\i46/n168 ),
    .B(\i46/n521 ),
    .Y(\i46/n285 ));
 AOI21xp5_ASAP7_75t_SL \i46/i201  (.A1(\i46/n65 ),
    .A2(\i46/n54 ),
    .B(\i46/n210 ),
    .Y(\i46/n283 ));
 NAND2xp5_ASAP7_75t_SL \i46/i202  (.A(\i46/n538 ),
    .B(\i46/n213 ),
    .Y(\i46/n282 ));
 NAND2xp5_ASAP7_75t_SL \i46/i203  (.A(\i46/n24 ),
    .B(\i46/n500 ),
    .Y(\i46/n280 ));
 NAND2xp5_ASAP7_75t_SL \i46/i204  (.A(\i46/n494 ),
    .B(\i46/n550 ),
    .Y(\i46/n279 ));
 NAND2xp5_ASAP7_75t_SL \i46/i205  (.A(\i46/n568 ),
    .B(\i46/n553 ),
    .Y(\i46/n277 ));
 NOR2x1_ASAP7_75t_SL \i46/i206  (.A(\i46/n197 ),
    .B(\i46/n180 ),
    .Y(\i46/n275 ));
 INVxp67_ASAP7_75t_SL \i46/i207  (.A(\i46/n251 ),
    .Y(\i46/n252 ));
 INVx1_ASAP7_75t_SL \i46/i208  (.A(\i46/n247 ),
    .Y(\i46/n248 ));
 INVx1_ASAP7_75t_SL \i46/i209  (.A(\i46/n243 ),
    .Y(\i46/n244 ));
 NAND4xp75_ASAP7_75t_SL \i46/i21  (.A(\i46/n396 ),
    .B(\i46/n427 ),
    .C(\i46/n401 ),
    .D(\i46/n391 ),
    .Y(\i46/n436 ));
 NAND4xp25_ASAP7_75t_SL \i46/i210  (.A(\i46/n99 ),
    .B(\i46/n502 ),
    .C(\i46/n474 ),
    .D(\i46/n557 ),
    .Y(\i46/n240 ));
 AOI31xp33_ASAP7_75t_SL \i46/i211  (.A1(\i46/n517 ),
    .A2(\i46/n62 ),
    .A3(\i46/n485 ),
    .B(\i46/n41 ),
    .Y(\i46/n239 ));
 NOR4xp25_ASAP7_75t_SL \i46/i212  (.A(\i46/n97 ),
    .B(\i46/n108 ),
    .C(\i46/n160 ),
    .D(\i46/n81 ),
    .Y(\i46/n238 ));
 AOI211xp5_ASAP7_75t_SL \i46/i213  (.A1(\i46/n115 ),
    .A2(\i46/n71 ),
    .B(\i46/n460 ),
    .C(\i46/n87 ),
    .Y(\i46/n237 ));
 NOR2xp33_ASAP7_75t_L \i46/i214  (.A(\i46/n528 ),
    .B(\i46/n207 ),
    .Y(\i46/n236 ));
 OAI31xp33_ASAP7_75t_SL \i46/i215  (.A1(\i46/n49 ),
    .A2(\i46/n523 ),
    .A3(\i46/n77 ),
    .B(\i46/n54 ),
    .Y(\i46/n235 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i46/i216  (.A1(\i46/n66 ),
    .A2(\i46/n43 ),
    .B(\i46/n73 ),
    .C(\i46/n510 ),
    .Y(\i46/n234 ));
 NOR2xp33_ASAP7_75t_SL \i46/i217  (.A(\i46/n448 ),
    .B(\i46/n165 ),
    .Y(\i46/n233 ));
 OAI222xp33_ASAP7_75t_SL \i46/i218  (.A1(\i46/n76 ),
    .A2(\i46/n41 ),
    .B1(\i46/n43 ),
    .B2(\i46/n19 ),
    .C1(\i46/n62 ),
    .C2(\i46/n59 ),
    .Y(\i46/n232 ));
 NAND2xp33_ASAP7_75t_L \i46/i219  (.A(\i46/n96 ),
    .B(\i46/n172 ),
    .Y(\i46/n231 ));
 AND3x4_ASAP7_75t_SL \i46/i22  (.A(\i46/n418 ),
    .B(\i46/n433 ),
    .C(\i46/n423 ),
    .Y(n28[7]));
 NAND2xp33_ASAP7_75t_SL \i46/i220  (.A(\i46/n203 ),
    .B(\i46/n548 ),
    .Y(\i46/n230 ));
 AOI22xp5_ASAP7_75t_SL \i46/i221  (.A1(\i46/n65 ),
    .A2(\i46/n94 ),
    .B1(\i46/n71 ),
    .B2(\i46/n67 ),
    .Y(\i46/n229 ));
 OA21x2_ASAP7_75t_SL \i46/i222  (.A1(\i46/n41 ),
    .A2(\i46/n562 ),
    .B(\i46/n110 ),
    .Y(\i46/n228 ));
 NAND2xp5_ASAP7_75t_SL \i46/i223  (.A(\i46/n169 ),
    .B(\i46/n216 ),
    .Y(\i46/n227 ));
 NAND4xp25_ASAP7_75t_SL \i46/i224  (.A(\i46/n566 ),
    .B(\i46/n130 ),
    .C(\i46/n91 ),
    .D(\i46/n516 ),
    .Y(\i46/n226 ));
 OAI221xp5_ASAP7_75t_SL \i46/i225  (.A1(\i46/n78 ),
    .A2(\i46/n73 ),
    .B1(\i46/n507 ),
    .B2(\i46/n18 ),
    .C(\i46/n95 ),
    .Y(\i46/n253 ));
 OAI222xp33_ASAP7_75t_SL \i46/i226  (.A1(\i46/n549 ),
    .A2(\i46/n45 ),
    .B1(\i46/n539 ),
    .B2(\i46/n59 ),
    .C1(\i46/n507 ),
    .C2(\i46/n68 ),
    .Y(\i46/n225 ));
 OAI221xp5_ASAP7_75t_SL \i46/i227  (.A1(\i46/n76 ),
    .A2(\i46/n68 ),
    .B1(\i46/n507 ),
    .B2(\i46/n60 ),
    .C(\i46/n178 ),
    .Y(\i46/n224 ));
 AND3x1_ASAP7_75t_SL \i46/i228  (.A(\i46/n109 ),
    .B(\i46/n502 ),
    .C(\i46/n509 ),
    .Y(\i46/n223 ));
 NAND2xp33_ASAP7_75t_SL \i46/i229  (.A(\i46/n489 ),
    .B(\i46/n193 ),
    .Y(\i46/n222 ));
 NAND4xp75_ASAP7_75t_SL \i46/i23  (.A(\i46/n400 ),
    .B(\i46/n379 ),
    .C(\i46/n409 ),
    .D(\i46/n426 ),
    .Y(\i46/n435 ));
 OAI221xp5_ASAP7_75t_SL \i46/i230  (.A1(\i46/n76 ),
    .A2(\i46/n70 ),
    .B1(\i46/n461 ),
    .B2(\i46/n19 ),
    .C(\i46/n202 ),
    .Y(\i46/n221 ));
 NAND3x1_ASAP7_75t_SL \i46/i231  (.A(\i46/n511 ),
    .B(\i46/n132 ),
    .C(\i46/n492 ),
    .Y(\i46/n251 ));
 AOI22xp5_ASAP7_75t_SL \i46/i232  (.A1(\i46/n131 ),
    .A2(\i46/n77 ),
    .B1(\i46/n523 ),
    .B2(\i46/n61 ),
    .Y(\i46/n250 ));
 AOI22xp5_ASAP7_75t_SL \i46/i233  (.A1(\i46/n80 ),
    .A2(\i46/n88 ),
    .B1(\i46/n42 ),
    .B2(\i46/n63 ),
    .Y(\i46/n249 ));
 AOI221x1_ASAP7_75t_SL \i46/i234  (.A1(\i46/n77 ),
    .A2(\i46/n61 ),
    .B1(\i46/n67 ),
    .B2(\i46/n69 ),
    .C(\i46/n571 ),
    .Y(\i46/n247 ));
 AOI211x1_ASAP7_75t_SL \i46/i235  (.A1(\i46/n89 ),
    .A2(\i46/n57 ),
    .B(\i46/n514 ),
    .C(\i46/n160 ),
    .Y(\i46/n246 ));
 OAI21xp5_ASAP7_75t_SL \i46/i236  (.A1(\i46/n485 ),
    .A2(\i46/n73 ),
    .B(\i46/n199 ),
    .Y(\i46/n245 ));
 NOR2x1_ASAP7_75t_SL \i46/i237  (.A(\i46/n111 ),
    .B(\i46/n456 ),
    .Y(\i46/n243 ));
 OAI221xp5_ASAP7_75t_SL \i46/i238  (.A1(\i46/n21 ),
    .A2(\i46/n78 ),
    .B1(\i46/n50 ),
    .B2(\i46/n60 ),
    .C(\i46/n567 ),
    .Y(\i46/n242 ));
 OAI211xp5_ASAP7_75t_SL \i46/i239  (.A1(\i46/n561 ),
    .A2(\i46/n60 ),
    .B(\i46/n98 ),
    .C(\i46/n551 ),
    .Y(\i46/n241 ));
 NAND2x1_ASAP7_75t_SL \i46/i24  (.A(\i46/n388 ),
    .B(\i46/n419 ),
    .Y(\i46/n434 ));
 NOR2xp33_ASAP7_75t_L \i46/i240  (.A(\i46/n118 ),
    .B(\i46/n171 ),
    .Y(\i46/n25 ));
 NOR2xp33_ASAP7_75t_SL \i46/i241  (.A(\i46/n119 ),
    .B(\i46/n453 ),
    .Y(\i46/n220 ));
 INVx1_ASAP7_75t_SL \i46/i242  (.A(\i46/n550 ),
    .Y(\i46/n218 ));
 INVx1_ASAP7_75t_SL \i46/i243  (.A(\i46/n215 ),
    .Y(\i46/n216 ));
 INVx1_ASAP7_75t_SL \i46/i244  (.A(\i46/n453 ),
    .Y(\i46/n214 ));
 INVxp67_ASAP7_75t_SL \i46/i245  (.A(\i46/n210 ),
    .Y(\i46/n211 ));
 INVx1_ASAP7_75t_SL \i46/i246  (.A(\i46/n207 ),
    .Y(\i46/n208 ));
 OAI21xp33_ASAP7_75t_SL \i46/i247  (.A1(\i46/n64 ),
    .A2(\i46/n51 ),
    .B(\i46/n515 ),
    .Y(\i46/n205 ));
 NAND2xp5_ASAP7_75t_SL \i46/i248  (.A(\i46/n555 ),
    .B(\i46/n114 ),
    .Y(\i46/n204 ));
 OAI21xp5_ASAP7_75t_SL \i46/i249  (.A1(\i46/n523 ),
    .A2(\i46/n440 ),
    .B(\i46/n74 ),
    .Y(\i46/n203 ));
 NOR2xp67_ASAP7_75t_SL \i46/i25  (.A(\i46/n420 ),
    .B(\i46/n381 ),
    .Y(\i46/n433 ));
 NOR2xp33_ASAP7_75t_SL \i46/i250  (.A(\i46/n120 ),
    .B(\i46/n150 ),
    .Y(\i46/n202 ));
 NAND2xp33_ASAP7_75t_L \i46/i251  (.A(\i46/n558 ),
    .B(\i46/n547 ),
    .Y(\i46/n201 ));
 NOR2xp33_ASAP7_75t_SL \i46/i252  (.A(\i46/n443 ),
    .B(\i46/n103 ),
    .Y(\i46/n200 ));
 OAI21xp5_ASAP7_75t_SL \i46/i253  (.A1(\i46/n65 ),
    .A2(\i46/n72 ),
    .B(\i46/n55 ),
    .Y(\i46/n199 ));
 OAI21xp5_ASAP7_75t_SL \i46/i254  (.A1(\i46/n47 ),
    .A2(\i46/n575 ),
    .B(\i46/n148 ),
    .Y(\i46/n198 ));
 OAI21xp5_ASAP7_75t_SL \i46/i255  (.A1(\i46/n19 ),
    .A2(\i46/n507 ),
    .B(\i46/n116 ),
    .Y(\i46/n197 ));
 OAI21xp5_ASAP7_75t_SL \i46/i256  (.A1(\i46/n65 ),
    .A2(\i46/n440 ),
    .B(\i46/n58 ),
    .Y(\i46/n196 ));
 OA21x2_ASAP7_75t_SL \i46/i257  (.A1(\i46/n56 ),
    .A2(\i46/n10 ),
    .B(\i46/n545 ),
    .Y(\i46/n219 ));
 AOI21xp33_ASAP7_75t_SL \i46/i258  (.A1(\i46/n59 ),
    .A2(\i46/n56 ),
    .B(\i46/n485 ),
    .Y(\i46/n195 ));
 OAI21xp5_ASAP7_75t_SL \i46/i259  (.A1(\i46/n69 ),
    .A2(\i46/n80 ),
    .B(\i46/n75 ),
    .Y(\i46/n194 ));
 NAND4xp75_ASAP7_75t_SL \i46/i26  (.A(\i46/n392 ),
    .B(\i46/n404 ),
    .C(\i46/n386 ),
    .D(\i46/n389 ),
    .Y(\i46/n432 ));
 OAI21xp5_ASAP7_75t_SL \i46/i260  (.A1(\i46/n58 ),
    .A2(\i46/n42 ),
    .B(\i46/n75 ),
    .Y(\i46/n193 ));
 AOI21xp33_ASAP7_75t_SL \i46/i261  (.A1(\i46/n53 ),
    .A2(\i46/n73 ),
    .B(\i46/n485 ),
    .Y(\i46/n192 ));
 OAI21xp5_ASAP7_75t_SL \i46/i262  (.A1(\i46/n47 ),
    .A2(\i46/n507 ),
    .B(\i46/n23 ),
    .Y(\i46/n191 ));
 AOI21xp33_ASAP7_75t_SL \i46/i263  (.A1(\i46/n66 ),
    .A2(\i46/n485 ),
    .B(\i46/n60 ),
    .Y(\i46/n190 ));
 NAND2xp5_ASAP7_75t_SL \i46/i264  (.A(\i46/n75 ),
    .B(\i46/n472 ),
    .Y(\i46/n24 ));
 NAND2xp5_ASAP7_75t_L \i46/i265  (.A(\i46/n491 ),
    .B(\i46/n512 ),
    .Y(\i46/n189 ));
 OAI22xp5_ASAP7_75t_SL \i46/i266  (.A1(\i46/n51 ),
    .A2(\i46/n76 ),
    .B1(\i46/n477 ),
    .B2(\i46/n10 ),
    .Y(\i46/n217 ));
 OAI22xp5_ASAP7_75t_SL \i46/i267  (.A1(\i46/n477 ),
    .A2(\i46/n507 ),
    .B1(\i46/n461 ),
    .B2(\i46/n59 ),
    .Y(\i46/n215 ));
 AOI22xp5_ASAP7_75t_SL \i46/i268  (.A1(\i46/n57 ),
    .A2(\i46/n77 ),
    .B1(\i46/n8 ),
    .B2(\i46/n72 ),
    .Y(\i46/n213 ));
 OAI22xp33_ASAP7_75t_SL \i46/i269  (.A1(\i46/n477 ),
    .A2(\i46/n78 ),
    .B1(\i46/n41 ),
    .B2(\i46/n549 ),
    .Y(\i46/n212 ));
 OR3x1_ASAP7_75t_SL \i46/i27  (.A(\i46/n412 ),
    .B(\i46/n410 ),
    .C(\i46/n393 ),
    .Y(\i46/n431 ));
 OAI22xp5_ASAP7_75t_SL \i46/i270  (.A1(\i46/n47 ),
    .A2(\i46/n78 ),
    .B1(\i46/n59 ),
    .B2(\i46/n575 ),
    .Y(\i46/n210 ));
 OAI21xp5_ASAP7_75t_SL \i46/i271  (.A1(\i46/n65 ),
    .A2(\i46/n44 ),
    .B(\i46/n74 ),
    .Y(\i46/n209 ));
 NOR2xp33_ASAP7_75t_L \i46/i272  (.A(\i46/n10 ),
    .B(\i46/n21 ),
    .Y(\i46/n207 ));
 NAND2xp33_ASAP7_75t_L \i46/i273  (.A(\i46/n98 ),
    .B(\i46/n551 ),
    .Y(\i46/n188 ));
 OAI21xp5_ASAP7_75t_SL \i46/i274  (.A1(\i46/n60 ),
    .A2(\i46/n539 ),
    .B(\i46/n484 ),
    .Y(\i46/n206 ));
 INVxp67_ASAP7_75t_SL \i46/i275  (.A(\i46/n186 ),
    .Y(\i46/n187 ));
 INVxp67_ASAP7_75t_SL \i46/i276  (.A(\i46/n493 ),
    .Y(\i46/n185 ));
 INVx1_ASAP7_75t_SL \i46/i277  (.A(\i46/n470 ),
    .Y(\i46/n184 ));
 INVx1_ASAP7_75t_SL \i46/i278  (.A(\i46/n182 ),
    .Y(\i46/n183 ));
 INVxp67_ASAP7_75t_SL \i46/i279  (.A(\i46/n565 ),
    .Y(\i46/n181 ));
 OR3x1_ASAP7_75t_SL \i46/i28  (.A(\i46/n413 ),
    .B(\i46/n378 ),
    .C(\i46/n352 ),
    .Y(\i46/n430 ));
 INVxp67_ASAP7_75t_SL \i46/i280  (.A(\i46/n448 ),
    .Y(\i46/n178 ));
 INVxp67_ASAP7_75t_SL \i46/i281  (.A(\i46/n457 ),
    .Y(\i46/n177 ));
 OAI21xp5_ASAP7_75t_SL \i46/i282  (.A1(\i46/n18 ),
    .A2(\i46/n549 ),
    .B(\i46/n106 ),
    .Y(\i46/n173 ));
 OAI21xp33_ASAP7_75t_SL \i46/i283  (.A1(\i46/n523 ),
    .A2(\i46/n44 ),
    .B(\i46/n48 ),
    .Y(\i46/n172 ));
 OAI22xp5_ASAP7_75t_SL \i46/i284  (.A1(\i46/n78 ),
    .A2(\i46/n45 ),
    .B1(\i46/n468 ),
    .B2(\i46/n10 ),
    .Y(\i46/n171 ));
 OAI21xp33_ASAP7_75t_SL \i46/i285  (.A1(\i46/n48 ),
    .A2(\i46/n71 ),
    .B(\i46/n523 ),
    .Y(\i46/n170 ));
 AOI22xp33_ASAP7_75t_SL \i46/i286  (.A1(\i46/n57 ),
    .A2(\i46/n65 ),
    .B1(\i46/n8 ),
    .B2(\i46/n523 ),
    .Y(\i46/n169 ));
 OAI22xp33_ASAP7_75t_SL \i46/i287  (.A1(\i46/n51 ),
    .A2(\i46/n485 ),
    .B1(\i46/n76 ),
    .B2(\i46/n53 ),
    .Y(\i46/n168 ));
 OAI22xp5_ASAP7_75t_SL \i46/i288  (.A1(\i46/n79 ),
    .A2(\i46/n549 ),
    .B1(\i46/n18 ),
    .B2(\i46/n76 ),
    .Y(\i46/n167 ));
 OAI22xp5_ASAP7_75t_SL \i46/i289  (.A1(\i46/n53 ),
    .A2(\i46/n549 ),
    .B1(\i46/n73 ),
    .B2(\i46/n66 ),
    .Y(\i46/n166 ));
 NAND3xp33_ASAP7_75t_SL \i46/i29  (.A(\i46/n424 ),
    .B(\i46/n392 ),
    .C(\i46/n409 ),
    .Y(\i46/n429 ));
 OAI22xp33_ASAP7_75t_SL \i46/i290  (.A1(\i46/n43 ),
    .A2(\i46/n51 ),
    .B1(\i46/n10 ),
    .B2(\i46/n45 ),
    .Y(\i46/n165 ));
 OAI22xp5_ASAP7_75t_SL \i46/i291  (.A1(\i46/n51 ),
    .A2(\i46/n78 ),
    .B1(\i46/n59 ),
    .B2(\i46/n10 ),
    .Y(\i46/n164 ));
 OAI21xp5_ASAP7_75t_SL \i46/i292  (.A1(\i46/n41 ),
    .A2(\i46/n539 ),
    .B(\i46/n104 ),
    .Y(\i46/n186 ));
 OAI22xp5_ASAP7_75t_SL \i46/i293  (.A1(\i46/n485 ),
    .A2(\i46/n18 ),
    .B1(\i46/n51 ),
    .B2(\i46/n62 ),
    .Y(\i46/n163 ));
 NAND2xp33_ASAP7_75t_SL \i46/i294  (.A(\i46/n544 ),
    .B(\i46/n161 ),
    .Y(\i46/n162 ));
 OAI22x1_ASAP7_75t_SL \i46/i295  (.A1(\i46/n19 ),
    .A2(\i46/n78 ),
    .B1(\i46/n468 ),
    .B2(\i46/n64 ),
    .Y(\i46/n182 ));
 AO22x2_ASAP7_75t_SL \i46/i296  (.A1(\i46/n80 ),
    .A2(\i46/n77 ),
    .B1(\i46/n46 ),
    .B2(\i46/n72 ),
    .Y(\i46/n180 ));
 OAI21xp5_ASAP7_75t_SL \i46/i297  (.A1(\i46/n68 ),
    .A2(\i46/n43 ),
    .B(\i46/n93 ),
    .Y(\i46/n179 ));
 OAI22xp5_ASAP7_75t_SL \i46/i298  (.A1(\i46/n66 ),
    .A2(\i46/n51 ),
    .B1(\i46/n62 ),
    .B2(\i46/n56 ),
    .Y(\i46/n176 ));
 OAI22xp5_ASAP7_75t_SL \i46/i299  (.A1(\i46/n45 ),
    .A2(\i46/n50 ),
    .B1(\i46/n59 ),
    .B2(\i46/n64 ),
    .Y(\i46/n175 ));
 INVx2_ASAP7_75t_SL \i46/i3  (.A(n29[2]),
    .Y(\i46/n3 ));
 NOR2x1_ASAP7_75t_SL \i46/i30  (.A(\i46/n333 ),
    .B(\i46/n410 ),
    .Y(\i46/n427 ));
 AOI22xp5_ASAP7_75t_SL \i46/i300  (.A1(\i46/n48 ),
    .A2(\i46/n72 ),
    .B1(\i46/n42 ),
    .B2(\i46/n49 ),
    .Y(\i46/n174 ));
 INVxp67_ASAP7_75t_SL \i46/i301  (.A(\i46/n514 ),
    .Y(\i46/n159 ));
 INVx1_ASAP7_75t_SL \i46/i302  (.A(\i46/n480 ),
    .Y(\i46/n158 ));
 INVxp67_ASAP7_75t_SL \i46/i303  (.A(\i46/n568 ),
    .Y(\i46/n157 ));
 INVxp67_ASAP7_75t_SL \i46/i304  (.A(\i46/n155 ),
    .Y(\i46/n156 ));
 INVxp67_ASAP7_75t_SL \i46/i305  (.A(\i46/n515 ),
    .Y(\i46/n154 ));
 INVxp67_ASAP7_75t_SL \i46/i306  (.A(\i46/n531 ),
    .Y(\i46/n152 ));
 INVxp67_ASAP7_75t_SL \i46/i307  (.A(\i46/n148 ),
    .Y(\i46/n149 ));
 INVxp67_ASAP7_75t_SL \i46/i308  (.A(\i46/n558 ),
    .Y(\i46/n147 ));
 INVxp67_ASAP7_75t_SL \i46/i309  (.A(\i46/n145 ),
    .Y(\i46/n146 ));
 NOR2x1_ASAP7_75t_SL \i46/i31  (.A(\i46/n394 ),
    .B(\i46/n390 ),
    .Y(\i46/n426 ));
 INVxp67_ASAP7_75t_SL \i46/i310  (.A(\i46/n567 ),
    .Y(\i46/n144 ));
 INVxp67_ASAP7_75t_SL \i46/i311  (.A(\i46/n142 ),
    .Y(\i46/n143 ));
 INVxp67_ASAP7_75t_SL \i46/i312  (.A(\i46/n140 ),
    .Y(\i46/n141 ));
 INVxp67_ASAP7_75t_SL \i46/i313  (.A(\i46/n21 ),
    .Y(\i46/n139 ));
 INVx2_ASAP7_75t_SL \i46/i314  (.A(\i46/n472 ),
    .Y(\i46/n138 ));
 NAND2xp5_ASAP7_75t_SL \i46/i315  (.A(\i46/n58 ),
    .B(\i46/n75 ),
    .Y(\i46/n161 ));
 NAND2xp5_ASAP7_75t_SL \i46/i316  (.A(\i46/n74 ),
    .B(\i46/n72 ),
    .Y(\i46/n137 ));
 NAND2xp5_ASAP7_75t_SL \i46/i317  (.A(\i46/n73 ),
    .B(\i46/n70 ),
    .Y(\i46/n136 ));
 NAND2xp5_ASAP7_75t_SL \i46/i318  (.A(\i46/n42 ),
    .B(\i46/n77 ),
    .Y(\i46/n135 ));
 NAND2xp33_ASAP7_75t_SL \i46/i319  (.A(\i46/n53 ),
    .B(\i46/n47 ),
    .Y(\i46/n134 ));
 NAND3xp33_ASAP7_75t_SL \i46/i32  (.A(\i46/n373 ),
    .B(\i46/n302 ),
    .C(\i46/n370 ),
    .Y(\i46/n425 ));
 NAND2xp5_ASAP7_75t_SL \i46/i320  (.A(\i46/n55 ),
    .B(\i46/n75 ),
    .Y(\i46/n133 ));
 NAND2xp5_ASAP7_75t_SL \i46/i321  (.A(\i46/n7 ),
    .B(\i46/n52 ),
    .Y(\i46/n132 ));
 NAND2xp5_ASAP7_75t_SL \i46/i322  (.A(\i46/n59 ),
    .B(\i46/n18 ),
    .Y(\i46/n131 ));
 NAND2xp5_ASAP7_75t_SL \i46/i323  (.A(\i46/n58 ),
    .B(\i46/n7 ),
    .Y(\i46/n130 ));
 NAND2xp5_ASAP7_75t_SL \i46/i324  (.A(\i46/n63 ),
    .B(\i46/n61 ),
    .Y(\i46/n129 ));
 NAND2xp5_ASAP7_75t_SL \i46/i325  (.A(\i46/n55 ),
    .B(\i46/n63 ),
    .Y(\i46/n128 ));
 AND2x2_ASAP7_75t_SL \i46/i326  (.A(\i46/n46 ),
    .B(\i46/n65 ),
    .Y(\i46/n160 ));
 NAND2xp5_ASAP7_75t_SL \i46/i327  (.A(\i46/n63 ),
    .B(\i46/n8 ),
    .Y(\i46/n23 ));
 NAND2xp5_ASAP7_75t_SL \i46/i328  (.A(\i46/n80 ),
    .B(\i46/n44 ),
    .Y(\i46/n155 ));
 NOR2xp33_ASAP7_75t_SL \i46/i329  (.A(\i46/n59 ),
    .B(\i46/n461 ),
    .Y(\i46/n127 ));
 NOR2x1_ASAP7_75t_SL \i46/i33  (.A(\i46/n399 ),
    .B(\i46/n361 ),
    .Y(\i46/n424 ));
 AND2x2_ASAP7_75t_SL \i46/i330  (.A(\i46/n58 ),
    .B(\i46/n49 ),
    .Y(\i46/n153 ));
 NOR2xp67_ASAP7_75t_SL \i46/i331  (.A(\i46/n56 ),
    .B(\i46/n507 ),
    .Y(\i46/n22 ));
 NAND2xp5_ASAP7_75t_SL \i46/i332  (.A(\i46/n57 ),
    .B(\i46/n7 ),
    .Y(\i46/n126 ));
 NAND2xp5_ASAP7_75t_SL \i46/i333  (.A(\i46/n67 ),
    .B(\i46/n57 ),
    .Y(\i46/n151 ));
 NAND2xp5_ASAP7_75t_SL \i46/i334  (.A(\i46/n49 ),
    .B(\i46/n52 ),
    .Y(\i46/n125 ));
 AND2x2_ASAP7_75t_SL \i46/i335  (.A(\i46/n55 ),
    .B(\i46/n7 ),
    .Y(\i46/n150 ));
 NOR2xp33_ASAP7_75t_SL \i46/i336  (.A(\i46/n19 ),
    .B(\i46/n10 ),
    .Y(\i46/n124 ));
 NAND2xp5_ASAP7_75t_SL \i46/i337  (.A(\i46/n57 ),
    .B(\i46/n44 ),
    .Y(\i46/n148 ));
 NOR2xp33_ASAP7_75t_SL \i46/i338  (.A(\i46/n54 ),
    .B(\i46/n74 ),
    .Y(\i46/n123 ));
 NOR2xp33_ASAP7_75t_SL \i46/i339  (.A(\i46/n51 ),
    .B(\i46/n575 ),
    .Y(\i46/n122 ));
 NOR5xp2_ASAP7_75t_SL \i46/i34  (.A(\i46/n363 ),
    .B(\i46/n314 ),
    .C(\i46/n354 ),
    .D(\i46/n279 ),
    .E(\i46/n451 ),
    .Y(\i46/n423 ));
 NAND2xp5_ASAP7_75t_SL \i46/i340  (.A(\i46/n80 ),
    .B(\i46/n440 ),
    .Y(\i46/n145 ));
 NAND2xp5_ASAP7_75t_SL \i46/i341  (.A(\i46/n80 ),
    .B(\i46/n63 ),
    .Y(\i46/n142 ));
 NAND2xp5_ASAP7_75t_SL \i46/i342  (.A(\i46/n58 ),
    .B(\i46/n67 ),
    .Y(\i46/n121 ));
 NOR2xp67_ASAP7_75t_SL \i46/i343  (.A(\i46/n74 ),
    .B(\i46/n58 ),
    .Y(\i46/n140 ));
 NOR2xp33_ASAP7_75t_SL \i46/i344  (.A(\i46/n539 ),
    .B(\i46/n73 ),
    .Y(\i46/n120 ));
 NOR2x1_ASAP7_75t_SL \i46/i345  (.A(\i46/n54 ),
    .B(\i46/n71 ),
    .Y(\i46/n21 ));
 INVxp67_ASAP7_75t_SL \i46/i346  (.A(\i46/n481 ),
    .Y(\i46/n119 ));
 INVxp67_ASAP7_75t_SL \i46/i347  (.A(\i46/n116 ),
    .Y(\i46/n117 ));
 INVx1_ASAP7_75t_SL \i46/i348  (.A(\i46/n517 ),
    .Y(\i46/n115 ));
 INVxp67_ASAP7_75t_SL \i46/i349  (.A(\i46/n566 ),
    .Y(\i46/n112 ));
 NOR3xp33_ASAP7_75t_SL \i46/i35  (.A(\i46/n359 ),
    .B(\i46/n375 ),
    .C(\i46/n408 ),
    .Y(\i46/n422 ));
 INVxp67_ASAP7_75t_SL \i46/i350  (.A(\i46/n110 ),
    .Y(\i46/n111 ));
 INVxp67_ASAP7_75t_SL \i46/i351  (.A(\i46/n108 ),
    .Y(\i46/n109 ));
 INVxp67_ASAP7_75t_SL \i46/i352  (.A(\i46/n106 ),
    .Y(\i46/n107 ));
 INVxp67_ASAP7_75t_R \i46/i353  (.A(\i46/n488 ),
    .Y(\i46/n105 ));
 INVxp67_ASAP7_75t_SL \i46/i354  (.A(\i46/n103 ),
    .Y(\i46/n104 ));
 INVxp67_ASAP7_75t_SL \i46/i355  (.A(\i46/n557 ),
    .Y(\i46/n102 ));
 INVxp67_ASAP7_75t_SL \i46/i356  (.A(\i46/n99 ),
    .Y(\i46/n100 ));
 INVx1_ASAP7_75t_SL \i46/i357  (.A(\i46/n96 ),
    .Y(\i46/n97 ));
 NAND2xp5_ASAP7_75t_SL \i46/i358  (.A(\i46/n71 ),
    .B(\i46/n65 ),
    .Y(\i46/n95 ));
 NAND2xp5_ASAP7_75t_SL \i46/i359  (.A(\i46/n48 ),
    .B(\i46/n65 ),
    .Y(\i46/n20 ));
 NOR2x1_ASAP7_75t_SL \i46/i36  (.A(\i46/n405 ),
    .B(\i46/n364 ),
    .Y(\i46/n421 ));
 NAND2xp5_ASAP7_75t_SL \i46/i360  (.A(\i46/n68 ),
    .B(\i46/n60 ),
    .Y(\i46/n94 ));
 NAND2xp5_ASAP7_75t_SL \i46/i361  (.A(\i46/n48 ),
    .B(\i46/n67 ),
    .Y(\i46/n93 ));
 NAND2xp5_ASAP7_75t_SL \i46/i362  (.A(\i46/n67 ),
    .B(\i46/n42 ),
    .Y(\i46/n92 ));
 NAND2xp5_ASAP7_75t_SL \i46/i363  (.A(\i46/n69 ),
    .B(\i46/n49 ),
    .Y(\i46/n91 ));
 NAND2xp5_ASAP7_75t_R \i46/i364  (.A(\i46/n61 ),
    .B(\i46/n440 ),
    .Y(\i46/n90 ));
 NAND2xp5_ASAP7_75t_L \i46/i365  (.A(\i46/n461 ),
    .B(\i46/n485 ),
    .Y(\i46/n89 ));
 NAND2xp33_ASAP7_75t_SL \i46/i366  (.A(\i46/n50 ),
    .B(\i46/n549 ),
    .Y(\i46/n88 ));
 NOR2xp33_ASAP7_75t_SL \i46/i367  (.A(\i46/n539 ),
    .B(\i46/n47 ),
    .Y(\i46/n87 ));
 AND2x2_ASAP7_75t_SL \i46/i368  (.A(\i46/n8 ),
    .B(\i46/n67 ),
    .Y(\i46/n118 ));
 NAND2xp5_ASAP7_75t_SL \i46/i369  (.A(\i46/n74 ),
    .B(\i46/n49 ),
    .Y(\i46/n116 ));
 NAND2xp5_ASAP7_75t_SL \i46/i37  (.A(\i46/n362 ),
    .B(\i46/n382 ),
    .Y(\i46/n420 ));
 NAND2xp5_ASAP7_75t_SL \i46/i370  (.A(\i46/n69 ),
    .B(\i46/n440 ),
    .Y(\i46/n114 ));
 NAND2xp5_ASAP7_75t_SL \i46/i371  (.A(\i46/n42 ),
    .B(\i46/n65 ),
    .Y(\i46/n86 ));
 AND2x2_ASAP7_75t_SL \i46/i372  (.A(\i46/n8 ),
    .B(\i46/n44 ),
    .Y(\i46/n113 ));
 NAND2xp5_ASAP7_75t_SL \i46/i373  (.A(\i46/n71 ),
    .B(\i46/n44 ),
    .Y(\i46/n110 ));
 NOR2xp67_ASAP7_75t_SL \i46/i374  (.A(\i46/n45 ),
    .B(\i46/n76 ),
    .Y(\i46/n108 ));
 NAND2xp5_ASAP7_75t_SL \i46/i375  (.A(\i46/n42 ),
    .B(\i46/n44 ),
    .Y(\i46/n106 ));
 NAND2xp33_ASAP7_75t_L \i46/i376  (.A(\i46/n43 ),
    .B(\i46/n64 ),
    .Y(\i46/n85 ));
 NOR2xp67_ASAP7_75t_R \i46/i377  (.A(\i46/n485 ),
    .B(\i46/n47 ),
    .Y(\i46/n103 ));
 NOR2xp33_ASAP7_75t_SL \i46/i378  (.A(\i46/n50 ),
    .B(\i46/n41 ),
    .Y(\i46/n84 ));
 NOR2xp67_ASAP7_75t_SL \i46/i379  (.A(\i46/n523 ),
    .B(\i46/n65 ),
    .Y(\i46/n101 ));
 NOR3x1_ASAP7_75t_SL \i46/i38  (.A(\i46/n27 ),
    .B(\i46/n377 ),
    .C(\i46/n305 ),
    .Y(\i46/n428 ));
 NAND2xp5_ASAP7_75t_SL \i46/i380  (.A(\i46/n8 ),
    .B(\i46/n72 ),
    .Y(\i46/n83 ));
 NAND2xp5_ASAP7_75t_SL \i46/i381  (.A(\i46/n48 ),
    .B(\i46/n440 ),
    .Y(\i46/n99 ));
 NAND2xp5_ASAP7_75t_SL \i46/i382  (.A(\i46/n69 ),
    .B(\i46/n72 ),
    .Y(\i46/n98 ));
 NOR2xp33_ASAP7_75t_SL \i46/i383  (.A(\i46/n477 ),
    .B(\i46/n10 ),
    .Y(\i46/n82 ));
 NOR2xp33_ASAP7_75t_SL \i46/i384  (.A(\i46/n477 ),
    .B(\i46/n539 ),
    .Y(\i46/n81 ));
 NAND2xp5_ASAP7_75t_SL \i46/i385  (.A(\i46/n48 ),
    .B(\i46/n75 ),
    .Y(\i46/n96 ));
 INVx1_ASAP7_75t_SL \i46/i386  (.A(\i46/n80 ),
    .Y(\i46/n79 ));
 INVx3_ASAP7_75t_SL \i46/i387  (.A(\i46/n78 ),
    .Y(\i46/n77 ));
 INVx4_ASAP7_75t_SL \i46/i388  (.A(\i46/n76 ),
    .Y(\i46/n75 ));
 INVx2_ASAP7_75t_SL \i46/i389  (.A(\i46/n74 ),
    .Y(\i46/n73 ));
 NOR3xp33_ASAP7_75t_SL \i46/i39  (.A(\i46/n321 ),
    .B(\i46/n27 ),
    .C(\i46/n402 ),
    .Y(\i46/n418 ));
 INVx2_ASAP7_75t_SL \i46/i390  (.A(\i46/n71 ),
    .Y(\i46/n70 ));
 INVx2_ASAP7_75t_SL \i46/i391  (.A(\i46/n69 ),
    .Y(\i46/n68 ));
 INVx3_ASAP7_75t_SL \i46/i392  (.A(\i46/n67 ),
    .Y(\i46/n66 ));
 INVx2_ASAP7_75t_SL \i46/i393  (.A(\i46/n65 ),
    .Y(\i46/n64 ));
 INVx2_ASAP7_75t_SL \i46/i394  (.A(\i46/n63 ),
    .Y(\i46/n62 ));
 INVx3_ASAP7_75t_SL \i46/i395  (.A(\i46/n61 ),
    .Y(\i46/n60 ));
 INVx3_ASAP7_75t_SL \i46/i396  (.A(\i46/n59 ),
    .Y(\i46/n58 ));
 AND2x4_ASAP7_75t_SL \i46/i397  (.A(\i46/n36 ),
    .B(\i46/n475 ),
    .Y(\i46/n80 ));
 OR2x4_ASAP7_75t_SL \i46/i398  (.A(\i46/n32 ),
    .B(\i46/n11 ),
    .Y(\i46/n78 ));
 OR2x6_ASAP7_75t_SL \i46/i399  (.A(\i46/n33 ),
    .B(\i46/n40 ),
    .Y(\i46/n76 ));
 INVx2_ASAP7_75t_SL \i46/i4  (.A(n29[0]),
    .Y(\i46/n4 ));
 NOR2xp67_ASAP7_75t_SL \i46/i40  (.A(\i46/n383 ),
    .B(\i46/n27 ),
    .Y(\i46/n417 ));
 AND2x4_ASAP7_75t_SL \i46/i400  (.A(\i46/n31 ),
    .B(\i46/n39 ),
    .Y(\i46/n74 ));
 AND2x4_ASAP7_75t_SL \i46/i401  (.A(\i46/n504 ),
    .B(\i46/n34 ),
    .Y(\i46/n72 ));
 AND2x4_ASAP7_75t_SL \i46/i402  (.A(\i46/n31 ),
    .B(\i46/n36 ),
    .Y(\i46/n71 ));
 AND2x4_ASAP7_75t_SL \i46/i403  (.A(\i46/n31 ),
    .B(\i46/n465 ),
    .Y(\i46/n69 ));
 AND2x4_ASAP7_75t_SL \i46/i404  (.A(\i46/n504 ),
    .B(\i46/n533 ),
    .Y(\i46/n67 ));
 AND2x4_ASAP7_75t_SL \i46/i405  (.A(\i46/n559 ),
    .B(\i46/n6 ),
    .Y(\i46/n65 ));
 AND2x4_ASAP7_75t_SL \i46/i406  (.A(\i46/n559 ),
    .B(\i46/n504 ),
    .Y(\i46/n63 ));
 AND2x4_ASAP7_75t_SL \i46/i407  (.A(\i46/n36 ),
    .B(\i46/n466 ),
    .Y(\i46/n61 ));
 OR2x6_ASAP7_75t_SL \i46/i408  (.A(\i46/n37 ),
    .B(\i46/n30 ),
    .Y(\i46/n59 ));
 INVx3_ASAP7_75t_SL \i46/i409  (.A(\i46/n57 ),
    .Y(\i46/n56 ));
 NOR3xp33_ASAP7_75t_SL \i46/i41  (.A(\i46/n360 ),
    .B(\i46/n355 ),
    .C(\i46/n13 ),
    .Y(\i46/n416 ));
 INVx3_ASAP7_75t_SL \i46/i410  (.A(\i46/n55 ),
    .Y(\i46/n19 ));
 INVx3_ASAP7_75t_SL \i46/i411  (.A(\i46/n54 ),
    .Y(\i46/n53 ));
 INVx3_ASAP7_75t_SL \i46/i412  (.A(\i46/n52 ),
    .Y(\i46/n51 ));
 INVx3_ASAP7_75t_SL \i46/i413  (.A(\i46/n50 ),
    .Y(\i46/n49 ));
 INVx5_ASAP7_75t_SL \i46/i414  (.A(\i46/n48 ),
    .Y(\i46/n47 ));
 INVx4_ASAP7_75t_SL \i46/i415  (.A(\i46/n46 ),
    .Y(\i46/n45 ));
 INVx3_ASAP7_75t_SL \i46/i416  (.A(\i46/n42 ),
    .Y(\i46/n41 ));
 AND2x4_ASAP7_75t_SL \i46/i417  (.A(\i46/n36 ),
    .B(\i46/n15 ),
    .Y(\i46/n57 ));
 AND2x4_ASAP7_75t_SL \i46/i418  (.A(\i46/n475 ),
    .B(\i46/n39 ),
    .Y(\i46/n55 ));
 AND2x4_ASAP7_75t_SL \i46/i419  (.A(\i46/n9 ),
    .B(\i46/n466 ),
    .Y(\i46/n54 ));
 NAND4xp25_ASAP7_75t_SL \i46/i42  (.A(\i46/n343 ),
    .B(\i46/n337 ),
    .C(\i46/n336 ),
    .D(\i46/n368 ),
    .Y(\i46/n415 ));
 OR2x2_ASAP7_75t_SL \i46/i420  (.A(\i46/n38 ),
    .B(\i46/n14 ),
    .Y(\i46/n18 ));
 AND2x4_ASAP7_75t_SL \i46/i421  (.A(\i46/n465 ),
    .B(\i46/n475 ),
    .Y(\i46/n52 ));
 NAND2x1p5_ASAP7_75t_SL \i46/i422  (.A(\i46/n559 ),
    .B(\i46/n497 ),
    .Y(\i46/n50 ));
 AND2x4_ASAP7_75t_SL \i46/i423  (.A(\i46/n465 ),
    .B(\i46/n15 ),
    .Y(\i46/n48 ));
 AND2x4_ASAP7_75t_SL \i46/i424  (.A(\i46/n9 ),
    .B(\i46/n15 ),
    .Y(\i46/n46 ));
 AND2x4_ASAP7_75t_SL \i46/i425  (.A(\i46/n5 ),
    .B(\i46/n34 ),
    .Y(\i46/n44 ));
 NAND2x1_ASAP7_75t_SL \i46/i426  (.A(\i46/n5 ),
    .B(\i46/n34 ),
    .Y(\i46/n43 ));
 AND2x4_ASAP7_75t_SL \i46/i427  (.A(\i46/n39 ),
    .B(\i46/n466 ),
    .Y(\i46/n42 ));
 INVx2_ASAP7_75t_SL \i46/i428  (.A(\i46/n497 ),
    .Y(\i46/n40 ));
 INVx2_ASAP7_75t_SL \i46/i429  (.A(\i46/n38 ),
    .Y(\i46/n39 ));
 NAND3xp33_ASAP7_75t_L \i46/i43  (.A(\i46/n319 ),
    .B(\i46/n337 ),
    .C(\i46/n387 ),
    .Y(\i46/n414 ));
 NAND2xp5_ASAP7_75t_SL \i46/i430  (.A(\i46/n16 ),
    .B(\i46/n3 ),
    .Y(\i46/n35 ));
 NAND2xp5_ASAP7_75t_SL \i46/i431  (.A(\i46/n2 ),
    .B(n29[5]),
    .Y(\i46/n38 ));
 NAND2x1p5_ASAP7_75t_SL \i46/i432  (.A(n29[4]),
    .B(n29[5]),
    .Y(\i46/n37 ));
 AND2x4_ASAP7_75t_SL \i46/i433  (.A(\i46/n1 ),
    .B(\i46/n2 ),
    .Y(\i46/n36 ));
 INVx2_ASAP7_75t_SL \i46/i434  (.A(\i46/n11 ),
    .Y(\i46/n34 ));
 INVx1_ASAP7_75t_SL \i46/i435  (.A(\i46/n533 ),
    .Y(\i46/n33 ));
 INVx2_ASAP7_75t_SL \i46/i436  (.A(\i46/n31 ),
    .Y(\i46/n30 ));
 NAND2xp5_ASAP7_75t_SL \i46/i437  (.A(\i46/n28 ),
    .B(\i46/n4 ),
    .Y(\i46/n29 ));
 NAND2x1_ASAP7_75t_SL \i46/i438  (.A(n29[3]),
    .B(\i46/n3 ),
    .Y(\i46/n32 ));
 AND2x2_ASAP7_75t_SL \i46/i439  (.A(n29[7]),
    .B(n29[6]),
    .Y(\i46/n31 ));
 NAND3xp33_ASAP7_75t_SL \i46/i44  (.A(\i46/n323 ),
    .B(\i46/n369 ),
    .C(\i46/n356 ),
    .Y(\i46/n413 ));
 INVx1_ASAP7_75t_SL \i46/i440  (.A(n29[1]),
    .Y(\i46/n28 ));
 INVx2_ASAP7_75t_SL \i46/i441  (.A(n29[6]),
    .Y(\i46/n17 ));
 INVx2_ASAP7_75t_SL \i46/i442  (.A(n29[3]),
    .Y(\i46/n16 ));
 INVx1_ASAP7_75t_SL \i46/i443  (.A(\i46/n369 ),
    .Y(\i46/n13 ));
 AND2x2_ASAP7_75t_L \i46/i444  (.A(\i46/n0 ),
    .B(n29[6]),
    .Y(\i46/n15 ));
 NAND2xp5_ASAP7_75t_SL \i46/i445  (.A(\i46/n0 ),
    .B(n29[6]),
    .Y(\i46/n14 ));
 OR2x2_ASAP7_75t_SL \i46/i446  (.A(\i46/n113 ),
    .B(\i46/n521 ),
    .Y(\i46/n12 ));
 OR2x2_ASAP7_75t_SL \i46/i447  (.A(n29[0]),
    .B(n29[1]),
    .Y(\i46/n11 ));
 AND2x4_ASAP7_75t_SL \i46/i448  (.A(\i46/n505 ),
    .B(\i46/n6 ),
    .Y(\i46/n440 ));
 NAND4xp25_ASAP7_75t_SL \i46/i449  (.A(\i46/n490 ),
    .B(\i46/n493 ),
    .C(\i46/n469 ),
    .D(\i46/n441 ),
    .Y(\i46/n442 ));
 NAND2xp5_ASAP7_75t_L \i46/i45  (.A(\i46/n578 ),
    .B(\i46/n403 ),
    .Y(\i46/n412 ));
 NAND2xp5_ASAP7_75t_SL \i46/i450  (.A(\i46/n8 ),
    .B(\i46/n440 ),
    .Y(\i46/n441 ));
 INVx1_ASAP7_75t_SL \i46/i451  (.A(\i46/n441 ),
    .Y(\i46/n443 ));
 NAND2xp5_ASAP7_75t_L \i46/i452  (.A(\i46/n441 ),
    .B(\i46/n135 ),
    .Y(\i46/n444 ));
 AO21x1_ASAP7_75t_SL \i46/i453  (.A1(\i46/n486 ),
    .A2(\i46/n61 ),
    .B(\i46/n482 ),
    .Y(\i46/n445 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i46/i454  (.A1(\i46/n74 ),
    .A2(\i46/n8 ),
    .B(\i46/n560 ),
    .C(\i46/n443 ),
    .Y(\i46/n446 ));
 AOI22xp33_ASAP7_75t_SL \i46/i455  (.A1(\i46/n80 ),
    .A2(\i46/n523 ),
    .B1(\i46/n57 ),
    .B2(\i46/n7 ),
    .Y(\i46/n447 ));
 OAI22xp5_ASAP7_75t_L \i46/i456  (.A1(\i46/n70 ),
    .A2(\i46/n485 ),
    .B1(\i46/n41 ),
    .B2(\i46/n450 ),
    .Y(\i46/n448 ));
 OAI22xp5_ASAP7_75t_SL \i46/i457  (.A1(\i46/n450 ),
    .A2(\i46/n140 ),
    .B1(\i46/n59 ),
    .B2(\i46/n535 ),
    .Y(\i46/n449 ));
 OAI211xp5_ASAP7_75t_SL \i46/i458  (.A1(\i46/n79 ),
    .A2(\i46/n450 ),
    .B(\i46/n158 ),
    .C(\i46/n114 ),
    .Y(\i46/n451 ));
 OAI222xp33_ASAP7_75t_SL \i46/i459  (.A1(\i46/n450 ),
    .A2(\i46/n70 ),
    .B1(\i46/n78 ),
    .B2(\i46/n68 ),
    .C1(\i46/n461 ),
    .C2(\i46/n53 ),
    .Y(\i46/n452 ));
 NAND2xp5_ASAP7_75t_L \i46/i46  (.A(\i46/n576 ),
    .B(\i46/n385 ),
    .Y(\i46/n411 ));
 OAI22xp5_ASAP7_75t_SL \i46/i460  (.A1(\i46/n79 ),
    .A2(\i46/n539 ),
    .B1(\i46/n47 ),
    .B2(\i46/n450 ),
    .Y(\i46/n453 ));
 OAI22xp5_ASAP7_75t_SL \i46/i461  (.A1(\i46/n60 ),
    .A2(\i46/n450 ),
    .B1(\i46/n507 ),
    .B2(\i46/n468 ),
    .Y(\i46/n454 ));
 AOI21xp33_ASAP7_75t_SL \i46/i462  (.A1(\i46/n507 ),
    .A2(\i46/n450 ),
    .B(\i46/n70 ),
    .Y(\i46/n455 ));
 OAI22xp33_ASAP7_75t_SL \i46/i463  (.A1(\i46/n461 ),
    .A2(\i46/n51 ),
    .B1(\i46/n450 ),
    .B2(\i46/n73 ),
    .Y(\i46/n456 ));
 OAI22xp5_ASAP7_75t_SL \i46/i464  (.A1(\i46/n53 ),
    .A2(\i46/n43 ),
    .B1(\i46/n59 ),
    .B2(\i46/n450 ),
    .Y(\i46/n457 ));
 OAI22x1_ASAP7_75t_L \i46/i465  (.A1(\i46/n56 ),
    .A2(\i46/n450 ),
    .B1(\i46/n60 ),
    .B2(\i46/n76 ),
    .Y(\i46/n458 ));
 NOR2xp33_ASAP7_75t_SL \i46/i466  (.A(\i46/n60 ),
    .B(\i46/n450 ),
    .Y(\i46/n459 ));
 NOR2xp33_ASAP7_75t_SL \i46/i467  (.A(\i46/n51 ),
    .B(\i46/n450 ),
    .Y(\i46/n460 ));
 NAND2x1_ASAP7_75t_SL \i46/i468  (.A(\i46/n504 ),
    .B(\i46/n34 ),
    .Y(\i46/n461 ));
 OAI21xp33_ASAP7_75t_L \i46/i469  (.A1(\i46/n462 ),
    .A2(\i46/n65 ),
    .B(\i46/n71 ),
    .Y(\i46/n463 ));
 NOR2x1_ASAP7_75t_SL \i46/i47  (.A(\i46/n393 ),
    .B(\i46/n384 ),
    .Y(\i46/n419 ));
 NAND2xp5_ASAP7_75t_SL \i46/i470  (.A(\i46/n10 ),
    .B(\i46/n461 ),
    .Y(\i46/n462 ));
 AOI211xp5_ASAP7_75t_SL \i46/i471  (.A1(\i46/n462 ),
    .A2(\i46/n46 ),
    .B(\i46/n261 ),
    .C(\i46/n204 ),
    .Y(\i46/n464 ));
 AND2x2_ASAP7_75t_SL \i46/i472  (.A(n29[4]),
    .B(\i46/n1 ),
    .Y(\i46/n465 ));
 AND2x4_ASAP7_75t_SL \i46/i473  (.A(n29[7]),
    .B(\i46/n17 ),
    .Y(\i46/n466 ));
 AND2x4_ASAP7_75t_SL \i46/i474  (.A(\i46/n465 ),
    .B(\i46/n466 ),
    .Y(\i46/n467 ));
 INVx2_ASAP7_75t_SL \i46/i475  (.A(\i46/n467 ),
    .Y(\i46/n468 ));
 OAI31xp33_ASAP7_75t_SL \i46/i476  (.A1(\i46/n42 ),
    .A2(\i46/n467 ),
    .A3(\i46/n61 ),
    .B(\i46/n77 ),
    .Y(\i46/n469 ));
 AOI22xp5_ASAP7_75t_SL \i46/i477  (.A1(\i46/n467 ),
    .A2(\i46/n44 ),
    .B1(\i46/n49 ),
    .B2(\i46/n55 ),
    .Y(\i46/n470 ));
 NOR2xp33_ASAP7_75t_L \i46/i478  (.A(\i46/n80 ),
    .B(\i46/n467 ),
    .Y(\i46/n471 ));
 OR2x2_ASAP7_75t_SL \i46/i479  (.A(\i46/n467 ),
    .B(\i46/n57 ),
    .Y(\i46/n472 ));
 NAND2xp33_ASAP7_75t_L \i46/i48  (.A(\i46/n372 ),
    .B(\i46/n345 ),
    .Y(\i46/n408 ));
 NAND2xp5_ASAP7_75t_SL \i46/i480  (.A(\i46/n467 ),
    .B(\i46/n67 ),
    .Y(\i46/n473 ));
 NAND2xp5_ASAP7_75t_SL \i46/i481  (.A(\i46/n467 ),
    .B(\i46/n72 ),
    .Y(\i46/n474 ));
 AND2x2_ASAP7_75t_SL \i46/i482  (.A(\i46/n0 ),
    .B(\i46/n17 ),
    .Y(\i46/n475 ));
 AND2x4_ASAP7_75t_SL \i46/i483  (.A(\i46/n475 ),
    .B(\i46/n9 ),
    .Y(\i46/n476 ));
 INVx2_ASAP7_75t_SL \i46/i484  (.A(\i46/n476 ),
    .Y(\i46/n477 ));
 AOI22xp5_ASAP7_75t_SL \i46/i485  (.A1(\i46/n476 ),
    .A2(\i46/n75 ),
    .B1(\i46/n74 ),
    .B2(\i46/n440 ),
    .Y(\i46/n478 ));
 AOI22xp5_ASAP7_75t_SL \i46/i486  (.A1(\i46/n476 ),
    .A2(\i46/n44 ),
    .B1(\i46/n54 ),
    .B2(\i46/n63 ),
    .Y(\i46/n479 ));
 AND2x2_ASAP7_75t_SL \i46/i487  (.A(\i46/n476 ),
    .B(\i46/n63 ),
    .Y(\i46/n480 ));
 NAND2xp5_ASAP7_75t_SL \i46/i488  (.A(\i46/n476 ),
    .B(\i46/n523 ),
    .Y(\i46/n481 ));
 AND2x2_ASAP7_75t_SL \i46/i489  (.A(\i46/n476 ),
    .B(\i46/n72 ),
    .Y(\i46/n482 ));
 NAND2xp33_ASAP7_75t_L \i46/i49  (.A(\i46/n578 ),
    .B(\i46/n350 ),
    .Y(\i46/n407 ));
 AND2x2_ASAP7_75t_SL \i46/i490  (.A(\i46/n476 ),
    .B(\i46/n49 ),
    .Y(\i46/n483 ));
 NAND2xp5_ASAP7_75t_SL \i46/i491  (.A(\i46/n476 ),
    .B(\i46/n67 ),
    .Y(\i46/n484 ));
 OR2x6_ASAP7_75t_SL \i46/i492  (.A(\i46/n29 ),
    .B(\i46/n35 ),
    .Y(\i46/n485 ));
 AOI22xp5_ASAP7_75t_R \i46/i493  (.A1(\i46/n486 ),
    .A2(\i46/n42 ),
    .B1(\i46/n476 ),
    .B2(\i46/n65 ),
    .Y(\i46/n487 ));
 INVx4_ASAP7_75t_SL \i46/i494  (.A(\i46/n485 ),
    .Y(\i46/n486 ));
 NAND2xp5_ASAP7_75t_SL \i46/i495  (.A(\i46/n486 ),
    .B(\i46/n476 ),
    .Y(\i46/n488 ));
 OAI21xp5_ASAP7_75t_SL \i46/i496  (.A1(\i46/n486 ),
    .A2(\i46/n44 ),
    .B(\i46/n467 ),
    .Y(\i46/n489 ));
 AOI22xp5_ASAP7_75t_SL \i46/i497  (.A1(\i46/n486 ),
    .A2(\i46/n467 ),
    .B1(\i46/n61 ),
    .B2(\i46/n72 ),
    .Y(\i46/n490 ));
 NAND2xp5_ASAP7_75t_SL \i46/i498  (.A(\i46/n486 ),
    .B(\i46/n69 ),
    .Y(\i46/n491 ));
 NAND2xp5_ASAP7_75t_SL \i46/i499  (.A(\i46/n486 ),
    .B(\i46/n46 ),
    .Y(\i46/n492 ));
 INVx2_ASAP7_75t_SL \i46/i5  (.A(\i46/n518 ),
    .Y(\i46/n5 ));
 NOR2xp33_ASAP7_75t_SL \i46/i50  (.A(\i46/n349 ),
    .B(\i46/n374 ),
    .Y(\i46/n406 ));
 AOI22xp5_ASAP7_75t_SL \i46/i500  (.A1(\i46/n486 ),
    .A2(\i46/n58 ),
    .B1(\i46/n42 ),
    .B2(\i46/n440 ),
    .Y(\i46/n493 ));
 AOI22xp5_ASAP7_75t_SL \i46/i501  (.A1(\i46/n486 ),
    .A2(\i46/n80 ),
    .B1(\i46/n42 ),
    .B2(\i46/n65 ),
    .Y(\i46/n494 ));
 AOI221xp5_ASAP7_75t_SL \i46/i502  (.A1(\i46/n55 ),
    .A2(\i46/n486 ),
    .B1(\i46/n44 ),
    .B2(\i46/n58 ),
    .C(\i46/n530 ),
    .Y(\i46/n495 ));
 AOI222xp33_ASAP7_75t_SL \i46/i503  (.A1(\i46/n67 ),
    .A2(\i46/n55 ),
    .B1(\i46/n8 ),
    .B2(\i46/n486 ),
    .C1(\i46/n63 ),
    .C2(\i46/n52 ),
    .Y(\i46/n496 ));
 AND2x2_ASAP7_75t_SL \i46/i504  (.A(\i46/n16 ),
    .B(\i46/n3 ),
    .Y(\i46/n497 ));
 AND2x4_ASAP7_75t_SL \i46/i505  (.A(\i46/n497 ),
    .B(\i46/n505 ),
    .Y(\i46/n498 ));
 NAND2xp5_ASAP7_75t_SL \i46/i506  (.A(\i46/n467 ),
    .B(\i46/n498 ),
    .Y(\i46/n499 ));
 INVx5_ASAP7_75t_SL \i46/i507  (.A(\i46/n498 ),
    .Y(\i46/n450 ));
 AOI22xp5_ASAP7_75t_SL \i46/i508  (.A1(\i46/n55 ),
    .A2(\i46/n498 ),
    .B1(\i46/n42 ),
    .B2(\i46/n72 ),
    .Y(\i46/n500 ));
 NAND2xp5_ASAP7_75t_SL \i46/i509  (.A(\i46/n54 ),
    .B(\i46/n498 ),
    .Y(\i46/n501 ));
 NAND3xp33_ASAP7_75t_SL \i46/i51  (.A(\i46/n340 ),
    .B(\i46/n347 ),
    .C(\i46/n508 ),
    .Y(\i46/n405 ));
 NAND2xp5_ASAP7_75t_SL \i46/i510  (.A(\i46/n8 ),
    .B(\i46/n498 ),
    .Y(\i46/n502 ));
 NAND2xp5_ASAP7_75t_SL \i46/i511  (.A(\i46/n48 ),
    .B(\i46/n498 ),
    .Y(\i46/n503 ));
 AND2x4_ASAP7_75t_SL \i46/i512  (.A(n29[2]),
    .B(n29[3]),
    .Y(\i46/n504 ));
 INVx2_ASAP7_75t_SL \i46/i513  (.A(\i46/n519 ),
    .Y(\i46/n505 ));
 AND2x4_ASAP7_75t_SL \i46/i514  (.A(\i46/n504 ),
    .B(\i46/n505 ),
    .Y(\i46/n506 ));
 INVx4_ASAP7_75t_SL \i46/i515  (.A(\i46/n506 ),
    .Y(\i46/n507 ));
 AOI211xp5_ASAP7_75t_SL \i46/i516  (.A1(\i46/n506 ),
    .A2(\i46/n58 ),
    .B(\i46/n556 ),
    .C(\i46/n150 ),
    .Y(\i46/n508 ));
 OAI21xp5_ASAP7_75t_SL \i46/i517  (.A1(\i46/n65 ),
    .A2(\i46/n506 ),
    .B(\i46/n80 ),
    .Y(\i46/n509 ));
 OAI21xp5_ASAP7_75t_SL \i46/i518  (.A1(\i46/n506 ),
    .A2(\i46/n49 ),
    .B(\i46/n69 ),
    .Y(\i46/n510 ));
 OAI21xp5_ASAP7_75t_SL \i46/i519  (.A1(\i46/n48 ),
    .A2(\i46/n61 ),
    .B(\i46/n506 ),
    .Y(\i46/n511 ));
 NOR2x1_ASAP7_75t_SL \i46/i52  (.A(\i46/n298 ),
    .B(\i46/n358 ),
    .Y(\i46/n404 ));
 NAND2xp5_ASAP7_75t_SL \i46/i520  (.A(\i46/n52 ),
    .B(\i46/n506 ),
    .Y(\i46/n512 ));
 NAND2xp5_ASAP7_75t_SL \i46/i521  (.A(\i46/n46 ),
    .B(\i46/n506 ),
    .Y(\i46/n513 ));
 AND2x2_ASAP7_75t_SL \i46/i522  (.A(\i46/n74 ),
    .B(\i46/n506 ),
    .Y(\i46/n514 ));
 NAND2xp5_ASAP7_75t_SL \i46/i523  (.A(\i46/n54 ),
    .B(\i46/n506 ),
    .Y(\i46/n515 ));
 NAND2xp5_ASAP7_75t_SL \i46/i524  (.A(\i46/n42 ),
    .B(\i46/n506 ),
    .Y(\i46/n516 ));
 NOR2x1_ASAP7_75t_SL \i46/i525  (.A(\i46/n506 ),
    .B(\i46/n72 ),
    .Y(\i46/n517 ));
 OR2x2_ASAP7_75t_SL \i46/i526  (.A(\i46/n3 ),
    .B(n29[3]),
    .Y(\i46/n518 ));
 NAND2xp5_ASAP7_75t_SL \i46/i527  (.A(\i46/n4 ),
    .B(n29[1]),
    .Y(\i46/n519 ));
 OAI22xp5_ASAP7_75t_SL \i46/i528  (.A1(\i46/n45 ),
    .A2(\i46/n450 ),
    .B1(\i46/n59 ),
    .B2(\i46/n520 ),
    .Y(\i46/n521 ));
 OR2x4_ASAP7_75t_SL \i46/i529  (.A(\i46/n518 ),
    .B(\i46/n519 ),
    .Y(\i46/n520 ));
 NOR2xp33_ASAP7_75t_SL \i46/i53  (.A(\i46/n365 ),
    .B(\i46/n279 ),
    .Y(\i46/n403 ));
 OAI221xp5_ASAP7_75t_SL \i46/i530  (.A1(\i46/n47 ),
    .A2(\i46/n43 ),
    .B1(\i46/n520 ),
    .B2(\i46/n41 ),
    .C(\i46/n488 ),
    .Y(\i46/n522 ));
 INVx4_ASAP7_75t_SL \i46/i531  (.A(\i46/n520 ),
    .Y(\i46/n523 ));
 OAI221xp5_ASAP7_75t_SL \i46/i532  (.A1(\i46/n539 ),
    .A2(\i46/n56 ),
    .B1(\i46/n45 ),
    .B2(\i46/n520 ),
    .C(\i46/n20 ),
    .Y(\i46/n524 ));
 AO21x1_ASAP7_75t_SL \i46/i533  (.A1(\i46/n520 ),
    .A2(\i46/n137 ),
    .B(\i46/n123 ),
    .Y(\i46/n525 ));
 AOI31xp33_ASAP7_75t_SL \i46/i534  (.A1(\i46/n45 ),
    .A2(\i46/n70 ),
    .A3(\i46/n60 ),
    .B(\i46/n520 ),
    .Y(\i46/n526 ));
 OAI22xp33_ASAP7_75t_SL \i46/i535  (.A1(\i46/n468 ),
    .A2(\i46/n78 ),
    .B1(\i46/n520 ),
    .B2(\i46/n51 ),
    .Y(\i46/n527 ));
 OAI21xp5_ASAP7_75t_SL \i46/i536  (.A1(\i46/n68 ),
    .A2(\i46/n520 ),
    .B(\i46/n548 ),
    .Y(\i46/n528 ));
 OA21x2_ASAP7_75t_SL \i46/i537  (.A1(\i46/n45 ),
    .A2(\i46/n520 ),
    .B(\i46/n20 ),
    .Y(\i46/n529 ));
 OAI22xp5_ASAP7_75t_SL \i46/i538  (.A1(\i46/n45 ),
    .A2(\i46/n43 ),
    .B1(\i46/n520 ),
    .B2(\i46/n468 ),
    .Y(\i46/n530 ));
 NOR2xp33_ASAP7_75t_SL \i46/i539  (.A(\i46/n520 ),
    .B(\i46/n56 ),
    .Y(\i46/n531 ));
 NAND2xp5_ASAP7_75t_SL \i46/i54  (.A(\i46/n372 ),
    .B(\i46/n367 ),
    .Y(\i46/n402 ));
 NOR2xp33_ASAP7_75t_SL \i46/i540  (.A(\i46/n520 ),
    .B(\i46/n468 ),
    .Y(\i46/n532 ));
 AND2x4_ASAP7_75t_SL \i46/i541  (.A(n29[0]),
    .B(\i46/n28 ),
    .Y(\i46/n533 ));
 NOR2xp33_ASAP7_75t_SL \i46/i542  (.A(\i46/n506 ),
    .B(\i46/n534 ),
    .Y(\i46/n535 ));
 AND2x4_ASAP7_75t_SL \i46/i543  (.A(\i46/n533 ),
    .B(\i46/n6 ),
    .Y(\i46/n534 ));
 OAI21xp5_ASAP7_75t_SL \i46/i544  (.A1(\i46/n506 ),
    .A2(\i46/n534 ),
    .B(\i46/n467 ),
    .Y(\i46/n536 ));
 OAI21xp5_ASAP7_75t_SL \i46/i545  (.A1(\i46/n534 ),
    .A2(\i46/n498 ),
    .B(\i46/n69 ),
    .Y(\i46/n537 ));
 AOI22xp5_ASAP7_75t_SL \i46/i546  (.A1(\i46/n57 ),
    .A2(\i46/n49 ),
    .B1(\i46/n476 ),
    .B2(\i46/n534 ),
    .Y(\i46/n538 ));
 INVx4_ASAP7_75t_SL \i46/i547  (.A(\i46/n534 ),
    .Y(\i46/n539 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i46/i548  (.A1(\i46/n49 ),
    .A2(\i46/n534 ),
    .B(\i46/n8 ),
    .C(\i46/n147 ),
    .Y(\i46/n540 ));
 AOI22xp5_ASAP7_75t_SL \i46/i549  (.A1(\i46/n74 ),
    .A2(\i46/n534 ),
    .B1(\i46/n69 ),
    .B2(\i46/n63 ),
    .Y(\i46/n541 ));
 NOR2x1_ASAP7_75t_SL \i46/i55  (.A(\i46/n451 ),
    .B(\i46/n374 ),
    .Y(\i46/n401 ));
 AOI22xp5_ASAP7_75t_SL \i46/i550  (.A1(\i46/n52 ),
    .A2(\i46/n49 ),
    .B1(\i46/n69 ),
    .B2(\i46/n534 ),
    .Y(\i46/n542 ));
 NAND2xp5_ASAP7_75t_SL \i46/i551  (.A(\i46/n534 ),
    .B(\i46/n52 ),
    .Y(\i46/n543 ));
 NAND2xp5_ASAP7_75t_SL \i46/i552  (.A(\i46/n534 ),
    .B(\i46/n55 ),
    .Y(\i46/n544 ));
 NAND2xp5_ASAP7_75t_SL \i46/i553  (.A(\i46/n54 ),
    .B(\i46/n534 ),
    .Y(\i46/n545 ));
 NAND2xp5_ASAP7_75t_SL \i46/i554  (.A(\i46/n8 ),
    .B(\i46/n534 ),
    .Y(\i46/n546 ));
 NAND2xp5_ASAP7_75t_SL \i46/i555  (.A(\i46/n71 ),
    .B(\i46/n534 ),
    .Y(\i46/n547 ));
 NAND2xp5_ASAP7_75t_SL \i46/i556  (.A(\i46/n46 ),
    .B(\i46/n534 ),
    .Y(\i46/n548 ));
 NAND2x1p5_ASAP7_75t_SL \i46/i557  (.A(\i46/n5 ),
    .B(\i46/n533 ),
    .Y(\i46/n549 ));
 AOI22xp5_ASAP7_75t_SL \i46/i558  (.A1(\i46/n476 ),
    .A2(\i46/n498 ),
    .B1(\i46/n69 ),
    .B2(\i46/n7 ),
    .Y(\i46/n550 ));
 NAND2xp5_ASAP7_75t_SL \i46/i559  (.A(\i46/n476 ),
    .B(\i46/n7 ),
    .Y(\i46/n551 ));
 NOR2x1_ASAP7_75t_SL \i46/i56  (.A(\i46/n348 ),
    .B(\i46/n359 ),
    .Y(\i46/n400 ));
 OAI31xp33_ASAP7_75t_SL \i46/i560  (.A1(\i46/n63 ),
    .A2(\i46/n7 ),
    .A3(\i46/n440 ),
    .B(\i46/n467 ),
    .Y(\i46/n552 ));
 AOI22xp5_ASAP7_75t_SL \i46/i561  (.A1(\i46/n71 ),
    .A2(\i46/n49 ),
    .B1(\i46/n467 ),
    .B2(\i46/n7 ),
    .Y(\i46/n553 ));
 NAND2xp5_ASAP7_75t_SL \i46/i562  (.A(\i46/n42 ),
    .B(\i46/n7 ),
    .Y(\i46/n554 ));
 NAND2xp33_ASAP7_75t_L \i46/i563  (.A(\i46/n7 ),
    .B(\i46/n69 ),
    .Y(\i46/n555 ));
 AO21x2_ASAP7_75t_SL \i46/i564  (.A1(\i46/n71 ),
    .A2(\i46/n7 ),
    .B(\i46/n176 ),
    .Y(\i46/n556 ));
 NAND2xp5_ASAP7_75t_SL \i46/i565  (.A(\i46/n7 ),
    .B(\i46/n48 ),
    .Y(\i46/n557 ));
 NAND2xp5_ASAP7_75t_SL \i46/i566  (.A(\i46/n74 ),
    .B(\i46/n7 ),
    .Y(\i46/n558 ));
 AND2x2_ASAP7_75t_SL \i46/i567  (.A(n29[0]),
    .B(n29[1]),
    .Y(\i46/n559 ));
 NOR2xp33_ASAP7_75t_SL \i46/i568  (.A(\i46/n560 ),
    .B(\i46/n7 ),
    .Y(\i46/n561 ));
 AND2x4_ASAP7_75t_SL \i46/i569  (.A(\i46/n559 ),
    .B(\i46/n5 ),
    .Y(\i46/n560 ));
 NAND2xp5_ASAP7_75t_SL \i46/i57  (.A(\i46/n464 ),
    .B(\i46/n353 ),
    .Y(\i46/n399 ));
 NOR2xp33_ASAP7_75t_SL \i46/i570  (.A(\i46/n560 ),
    .B(\i46/n498 ),
    .Y(\i46/n562 ));
 AOI22xp5_ASAP7_75t_SL \i46/i571  (.A1(\i46/n560 ),
    .A2(\i46/n476 ),
    .B1(\i46/n71 ),
    .B2(\i46/n63 ),
    .Y(\i46/n563 ));
 OAI21xp5_ASAP7_75t_SL \i46/i572  (.A1(\i46/n560 ),
    .A2(\i46/n65 ),
    .B(\i46/n467 ),
    .Y(\i46/n564 ));
 AOI22xp5_ASAP7_75t_SL \i46/i573  (.A1(\i46/n467 ),
    .A2(\i46/n49 ),
    .B1(\i46/n42 ),
    .B2(\i46/n560 ),
    .Y(\i46/n565 ));
 NAND2xp5_ASAP7_75t_SL \i46/i574  (.A(\i46/n71 ),
    .B(\i46/n560 ),
    .Y(\i46/n566 ));
 NAND2xp5_ASAP7_75t_SL \i46/i575  (.A(\i46/n560 ),
    .B(\i46/n55 ),
    .Y(\i46/n567 ));
 NAND2xp5_ASAP7_75t_SL \i46/i576  (.A(\i46/n69 ),
    .B(\i46/n560 ),
    .Y(\i46/n568 ));
 NAND2xp5_ASAP7_75t_SL \i46/i577  (.A(\i46/n58 ),
    .B(\i46/n560 ),
    .Y(\i46/n569 ));
 NAND2xp5_ASAP7_75t_SL \i46/i578  (.A(\i46/n74 ),
    .B(\i46/n560 ),
    .Y(\i46/n570 ));
 OA21x2_ASAP7_75t_SL \i46/i579  (.A1(\i46/n8 ),
    .A2(\i46/n80 ),
    .B(\i46/n560 ),
    .Y(\i46/n571 ));
 NOR5xp2_ASAP7_75t_SL \i46/i58  (.A(\i46/n241 ),
    .B(\i46/n524 ),
    .C(\i46/n253 ),
    .D(\i46/n26 ),
    .E(\i46/n224 ),
    .Y(\i46/n398 ));
 AOI22xp5_ASAP7_75t_SL \i46/i580  (.A1(\i46/n75 ),
    .A2(\i46/n136 ),
    .B1(\i46/n52 ),
    .B2(\i46/n560 ),
    .Y(\i46/n572 ));
 AOI21xp5_ASAP7_75t_SL \i46/i581  (.A1(\i46/n472 ),
    .A2(\i46/n560 ),
    .B(\i46/n191 ),
    .Y(\i46/n573 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i46/i582  (.A1(\i46/n560 ),
    .A2(\i46/n44 ),
    .B(\i46/n61 ),
    .C(\i46/n118 ),
    .Y(\i46/n574 ));
 INVx2_ASAP7_75t_SL \i46/i583  (.A(\i46/n560 ),
    .Y(\i46/n575 ));
 AND4x1_ASAP7_75t_SL \i46/i584  (.A(\i46/n243 ),
    .B(\i46/n554 ),
    .C(\i46/n86 ),
    .D(\i46/n318 ),
    .Y(\i46/n576 ));
 AND4x1_ASAP7_75t_SL \i46/i585  (.A(\i46/n496 ),
    .B(\i46/n281 ),
    .C(\i46/n581 ),
    .D(\i46/n219 ),
    .Y(\i46/n577 ));
 AND4x1_ASAP7_75t_SL \i46/i586  (.A(\i46/n233 ),
    .B(\i46/n283 ),
    .C(\i46/n572 ),
    .D(\i46/n496 ),
    .Y(\i46/n578 ));
 NAND3xp33_ASAP7_75t_SL \i46/i587  (.A(\i46/n579 ),
    .B(\i46/n213 ),
    .C(\i46/n273 ),
    .Y(\i46/n580 ));
 AO21x1_ASAP7_75t_SL \i46/i588  (.A1(\i46/n56 ),
    .A2(\i46/n45 ),
    .B(\i46/n575 ),
    .Y(\i46/n579 ));
 AOI21xp5_ASAP7_75t_SL \i46/i589  (.A1(\i46/n46 ),
    .A2(\i46/n63 ),
    .B(\i46/n530 ),
    .Y(\i46/n581 ));
 NOR2x1_ASAP7_75t_SL \i46/i59  (.A(\i46/n13 ),
    .B(\i46/n360 ),
    .Y(\i46/n397 ));
 INVx1_ASAP7_75t_SL \i46/i6  (.A(\i46/n32 ),
    .Y(\i46/n6 ));
 NAND2xp5_ASAP7_75t_SL \i46/i60  (.A(\i46/n357 ),
    .B(\i46/n338 ),
    .Y(\i46/n410 ));
 NOR2x1_ASAP7_75t_SL \i46/i61  (.A(\i46/n375 ),
    .B(\i46/n359 ),
    .Y(\i46/n396 ));
 NOR2x1_ASAP7_75t_SL \i46/i62  (.A(\i46/n297 ),
    .B(\i46/n358 ),
    .Y(\i46/n409 ));
 INVxp67_ASAP7_75t_SL \i46/i63  (.A(\i46/n394 ),
    .Y(\i46/n395 ));
 INVxp67_ASAP7_75t_SL \i46/i64  (.A(\i46/n390 ),
    .Y(\i46/n391 ));
 AND5x1_ASAP7_75t_SL \i46/i65  (.A(\i46/n311 ),
    .B(\i46/n581 ),
    .C(\i46/n303 ),
    .D(\i46/n540 ),
    .E(\i46/n209 ),
    .Y(\i46/n389 ));
 NOR3xp33_ASAP7_75t_SL \i46/i66  (.A(\i46/n320 ),
    .B(\i46/n301 ),
    .C(\i46/n284 ),
    .Y(\i46/n388 ));
 NOR3xp33_ASAP7_75t_SL \i46/i67  (.A(\i46/n442 ),
    .B(\i46/n285 ),
    .C(\i46/n240 ),
    .Y(\i46/n387 ));
 AND5x1_ASAP7_75t_SL \i46/i68  (.A(\i46/n275 ),
    .B(\i46/n288 ),
    .C(\i46/n269 ),
    .D(\i46/n278 ),
    .E(\i46/n214 ),
    .Y(\i46/n386 ));
 NOR2xp33_ASAP7_75t_SL \i46/i69  (.A(\i46/n346 ),
    .B(\i46/n351 ),
    .Y(\i46/n385 ));
 INVx2_ASAP7_75t_SL \i46/i7  (.A(\i46/n549 ),
    .Y(\i46/n7 ));
 NAND4xp25_ASAP7_75t_SL \i46/i70  (.A(\i46/n329 ),
    .B(\i46/n337 ),
    .C(\i46/n342 ),
    .D(\i46/n325 ),
    .Y(\i46/n384 ));
 NAND5xp2_ASAP7_75t_SL \i46/i71  (.A(\i46/n310 ),
    .B(\i46/n187 ),
    .C(\i46/n267 ),
    .D(\i46/n177 ),
    .E(\i46/n250 ),
    .Y(\i46/n383 ));
 NOR4xp25_ASAP7_75t_SL \i46/i72  (.A(\i46/n299 ),
    .B(\i46/n524 ),
    .C(\i46/n254 ),
    .D(\i46/n234 ),
    .Y(\i46/n382 ));
 NAND4xp25_ASAP7_75t_SL \i46/i73  (.A(\i46/n318 ),
    .B(\i46/n331 ),
    .C(\i46/n334 ),
    .D(\i46/n336 ),
    .Y(\i46/n381 ));
 NAND4xp25_ASAP7_75t_SL \i46/i74  (.A(\i46/n344 ),
    .B(\i46/n342 ),
    .C(\i46/n529 ),
    .D(\i46/n208 ),
    .Y(\i46/n380 ));
 NOR2x1_ASAP7_75t_SL \i46/i75  (.A(\i46/n445 ),
    .B(\i46/n371 ),
    .Y(\i46/n379 ));
 NAND3xp33_ASAP7_75t_SL \i46/i76  (.A(\i46/n336 ),
    .B(\i46/n309 ),
    .C(\i46/n499 ),
    .Y(\i46/n394 ));
 NAND4xp75_ASAP7_75t_SL \i46/i77  (.A(\i46/n246 ),
    .B(\i46/n223 ),
    .C(\i46/n296 ),
    .D(\i46/n23 ),
    .Y(\i46/n393 ));
 NAND2xp33_ASAP7_75t_L \i46/i78  (.A(\i46/n317 ),
    .B(\i46/n376 ),
    .Y(\i46/n378 ));
 AND2x2_ASAP7_75t_SL \i46/i79  (.A(\i46/n319 ),
    .B(\i46/n366 ),
    .Y(\i46/n392 ));
 INVx2_ASAP7_75t_SL \i46/i8  (.A(\i46/n18 ),
    .Y(\i46/n8 ));
 NAND2x1p5_ASAP7_75t_SL \i46/i80  (.A(\i46/n373 ),
    .B(\i46/n330 ),
    .Y(\i46/n390 ));
 INVxp67_ASAP7_75t_SL \i46/i81  (.A(\i46/n376 ),
    .Y(\i46/n377 ));
 INVxp67_ASAP7_75t_SL \i46/i82  (.A(\i46/n370 ),
    .Y(\i46/n371 ));
 NOR5xp2_ASAP7_75t_SL \i46/i83  (.A(\i46/n263 ),
    .B(\i46/n239 ),
    .C(\i46/n182 ),
    .D(\i46/n480 ),
    .E(\i46/n532 ),
    .Y(\i46/n368 ));
 NOR3xp33_ASAP7_75t_SL \i46/i84  (.A(\i46/n341 ),
    .B(\i46/n259 ),
    .C(\i46/n452 ),
    .Y(\i46/n367 ));
 NOR2xp33_ASAP7_75t_SL \i46/i85  (.A(\i46/n339 ),
    .B(\i46/n290 ),
    .Y(\i46/n366 ));
 NOR2x1_ASAP7_75t_SL \i46/i86  (.A(\i46/n304 ),
    .B(\i46/n276 ),
    .Y(\i46/n376 ));
 NAND3xp33_ASAP7_75t_SL \i46/i87  (.A(\i46/n249 ),
    .B(\i46/n552 ),
    .C(\i46/n563 ),
    .Y(\i46/n365 ));
 NAND2xp5_ASAP7_75t_L \i46/i88  (.A(\i46/n338 ),
    .B(\i46/n308 ),
    .Y(\i46/n364 ));
 NAND2xp5_ASAP7_75t_SL \i46/i89  (.A(\i46/n289 ),
    .B(\i46/n328 ),
    .Y(\i46/n363 ));
 INVx2_ASAP7_75t_SL \i46/i9  (.A(\i46/n37 ),
    .Y(\i46/n9 ));
 NAND3xp33_ASAP7_75t_SL \i46/i90  (.A(\i46/n581 ),
    .B(\i46/n236 ),
    .C(\i46/n219 ),
    .Y(\i46/n375 ));
 NOR3xp33_ASAP7_75t_SL \i46/i91  (.A(\i46/n312 ),
    .B(\i46/n12 ),
    .C(\i46/n221 ),
    .Y(\i46/n362 ));
 NAND2xp5_ASAP7_75t_SL \i46/i92  (.A(\i46/n501 ),
    .B(\i46/n318 ),
    .Y(\i46/n374 ));
 OR3x1_ASAP7_75t_SL \i46/i93  (.A(\i46/n241 ),
    .B(\i46/n253 ),
    .C(\i46/n26 ),
    .Y(\i46/n361 ));
 NOR2x1_ASAP7_75t_SL \i46/i94  (.A(\i46/n452 ),
    .B(\i46/n341 ),
    .Y(\i46/n373 ));
 NOR2xp33_ASAP7_75t_L \i46/i95  (.A(\i46/n300 ),
    .B(\i46/n287 ),
    .Y(\i46/n372 ));
 NOR2xp67_ASAP7_75t_SL \i46/i96  (.A(\i46/n242 ),
    .B(\i46/n327 ),
    .Y(\i46/n370 ));
 NOR3x1_ASAP7_75t_SL \i46/i97  (.A(\i46/n248 ),
    .B(\i46/n166 ),
    .C(\i46/n293 ),
    .Y(\i46/n369 ));
 NOR3xp33_ASAP7_75t_SL \i46/i98  (.A(\i46/n255 ),
    .B(\i46/n186 ),
    .C(\i46/n245 ),
    .Y(\i46/n357 ));
 NOR2xp33_ASAP7_75t_SL \i46/i99  (.A(\i46/n580 ),
    .B(\i46/n315 ),
    .Y(\i46/n356 ));
 OAI22xp5_ASAP7_75t_SL i460 (.A1(n758),
    .A2(n270),
    .B1(n759),
    .B2(n1154),
    .Y(n1012));
 OAI22xp5_ASAP7_75t_SL i461 (.A1(n842),
    .A2(n786),
    .B1(n843),
    .B2(n785),
    .Y(n1011));
 OAI22xp5_ASAP7_75t_SL i462 (.A1(n845),
    .A2(n768),
    .B1(n767),
    .B2(n844),
    .Y(n1010));
 XNOR2xp5_ASAP7_75t_SL i463 (.A(n599),
    .B(n776),
    .Y(n1009));
 AOI22xp5_ASAP7_75t_SL i464 (.A1(n837),
    .A2(n793),
    .B1(n838),
    .B2(n794),
    .Y(n1008));
 OAI22xp5_ASAP7_75t_SL i465 (.A1(n835),
    .A2(n786),
    .B1(n834),
    .B2(n785),
    .Y(n1007));
 OAI22xp5_ASAP7_75t_SL i466 (.A1(n830),
    .A2(n805),
    .B1(n806),
    .B2(n831),
    .Y(n1006));
 OAI22xp5_ASAP7_75t_SL i467 (.A1(n829),
    .A2(n805),
    .B1(n806),
    .B2(n828),
    .Y(n1005));
 OAI22xp5_ASAP7_75t_SL i468 (.A1(n870),
    .A2(n235),
    .B1(n1151),
    .B2(n871),
    .Y(n1004));
 AOI22xp5_ASAP7_75t_SL i469 (.A1(n826),
    .A2(n1232),
    .B1(n827),
    .B2(n777),
    .Y(n1003));
 INVx2_ASAP7_75t_SL \i47/i0  (.A(n27[7]),
    .Y(\i47/n0 ));
 INVxp67_ASAP7_75t_SL \i47/i1  (.A(n27[4]),
    .Y(\i47/n1 ));
 AND5x2_ASAP7_75t_SL \i47/i10  (.A(\i47/n406 ),
    .B(\i47/n397 ),
    .C(\i47/n399 ),
    .D(\i47/n386 ),
    .E(\i47/n487 ),
    .Y(n26[6]));
 NAND3xp33_ASAP7_75t_L \i47/i100  (.A(\i47/n217 ),
    .B(\i47/n241 ),
    .C(\i47/n300 ),
    .Y(\i47/n331 ));
 NOR5xp2_ASAP7_75t_SL \i47/i101  (.A(\i47/n216 ),
    .B(\i47/n226 ),
    .C(\i47/n454 ),
    .D(\i47/n94 ),
    .E(\i47/n77 ),
    .Y(\i47/n330 ));
 NAND5xp2_ASAP7_75t_SL \i47/i102  (.A(\i47/n23 ),
    .B(\i47/n278 ),
    .C(\i47/n545 ),
    .D(\i47/n500 ),
    .E(\i47/n157 ),
    .Y(\i47/n329 ));
 NAND4xp25_ASAP7_75t_R \i47/i103  (.A(\i47/n513 ),
    .B(\i47/n179 ),
    .C(\i47/n508 ),
    .D(\i47/n18 ),
    .Y(\i47/n328 ));
 NOR5xp2_ASAP7_75t_SL \i47/i104  (.A(\i47/n185 ),
    .B(\i47/n219 ),
    .C(\i47/n174 ),
    .D(\i47/n152 ),
    .E(\i47/n151 ),
    .Y(\i47/n327 ));
 NOR2xp33_ASAP7_75t_SL \i47/i105  (.A(\i47/n292 ),
    .B(\i47/n321 ),
    .Y(\i47/n326 ));
 NOR2xp33_ASAP7_75t_SL \i47/i106  (.A(\i47/n282 ),
    .B(\i47/n307 ),
    .Y(\i47/n325 ));
 NAND3x1_ASAP7_75t_SL \i47/i107  (.A(\i47/n183 ),
    .B(\i47/n306 ),
    .C(\i47/n277 ),
    .Y(\i47/n342 ));
 NAND3x1_ASAP7_75t_SL \i47/i108  (.A(\i47/n272 ),
    .B(\i47/n255 ),
    .C(\i47/n423 ),
    .Y(\i47/n341 ));
 AOI21xp5_ASAP7_75t_L \i47/i109  (.A1(\i47/n546 ),
    .A2(\i47/n510 ),
    .B(\i47/n135 ),
    .Y(\i47/n318 ));
 AND3x4_ASAP7_75t_SL \i47/i11  (.A(\i47/n406 ),
    .B(\i47/n415 ),
    .C(\i47/n394 ),
    .Y(n26[1]));
 NOR2xp33_ASAP7_75t_SL \i47/i110  (.A(\i47/n418 ),
    .B(\i47/n263 ),
    .Y(\i47/n317 ));
 NAND2xp5_ASAP7_75t_SL \i47/i111  (.A(\i47/n254 ),
    .B(\i47/n281 ),
    .Y(\i47/n316 ));
 NOR2xp33_ASAP7_75t_SL \i47/i112  (.A(\i47/n280 ),
    .B(\i47/n24 ),
    .Y(\i47/n315 ));
 NOR2xp33_ASAP7_75t_SL \i47/i113  (.A(\i47/n259 ),
    .B(\i47/n268 ),
    .Y(\i47/n314 ));
 NOR2xp67_ASAP7_75t_SL \i47/i114  (.A(\i47/n142 ),
    .B(\i47/n265 ),
    .Y(\i47/n313 ));
 NOR2xp67_ASAP7_75t_SL \i47/i115  (.A(\i47/n479 ),
    .B(\i47/n263 ),
    .Y(\i47/n312 ));
 NOR4xp25_ASAP7_75t_SL \i47/i116  (.A(\i47/n243 ),
    .B(\i47/n520 ),
    .C(\i47/n479 ),
    .D(\i47/n480 ),
    .Y(\i47/n311 ));
 NAND2xp5_ASAP7_75t_SL \i47/i117  (.A(\i47/n446 ),
    .B(\i47/n248 ),
    .Y(\i47/n310 ));
 NOR4xp25_ASAP7_75t_SL \i47/i118  (.A(\i47/n92 ),
    .B(\i47/n202 ),
    .C(\i47/n176 ),
    .D(\i47/n188 ),
    .Y(\i47/n309 ));
 NOR3xp33_ASAP7_75t_SL \i47/i119  (.A(\i47/n206 ),
    .B(\i47/n171 ),
    .C(\i47/n569 ),
    .Y(\i47/n308 ));
 NOR2x1p5_ASAP7_75t_SL \i47/i12  (.A(\i47/n416 ),
    .B(\i47/n407 ),
    .Y(n26[5]));
 NAND2xp33_ASAP7_75t_SL \i47/i120  (.A(\i47/n539 ),
    .B(\i47/n557 ),
    .Y(\i47/n307 ));
 NOR2x1p5_ASAP7_75t_SL \i47/i121  (.A(\i47/n222 ),
    .B(\i47/n240 ),
    .Y(\i47/n306 ));
 NAND2xp33_ASAP7_75t_SL \i47/i122  (.A(\i47/n279 ),
    .B(\i47/n261 ),
    .Y(\i47/n305 ));
 NAND3xp33_ASAP7_75t_SL \i47/i123  (.A(\i47/n22 ),
    .B(\i47/n495 ),
    .C(\i47/n447 ),
    .Y(\i47/n304 ));
 NOR3xp33_ASAP7_75t_SL \i47/i124  (.A(\i47/n529 ),
    .B(\i47/n180 ),
    .C(\i47/n566 ),
    .Y(\i47/n324 ));
 NAND2xp5_ASAP7_75t_SL \i47/i125  (.A(\i47/n12 ),
    .B(\i47/n513 ),
    .Y(\i47/n323 ));
 NOR2x1_ASAP7_75t_SL \i47/i126  (.A(\i47/n221 ),
    .B(\i47/n238 ),
    .Y(\i47/n322 ));
 NAND2xp67_ASAP7_75t_SL \i47/i127  (.A(\i47/n545 ),
    .B(\i47/n244 ),
    .Y(\i47/n321 ));
 NOR2x1_ASAP7_75t_SL \i47/i128  (.A(\i47/n223 ),
    .B(\i47/n266 ),
    .Y(\i47/n320 ));
 NOR3x1_ASAP7_75t_SL \i47/i129  (.A(\i47/n174 ),
    .B(\i47/n473 ),
    .C(\i47/n149 ),
    .Y(\i47/n319 ));
 AND2x4_ASAP7_75t_SL \i47/i13  (.A(\i47/n417 ),
    .B(\i47/n400 ),
    .Y(n26[0]));
 INVx1_ASAP7_75t_SL \i47/i130  (.A(\i47/n25 ),
    .Y(\i47/n301 ));
 NOR4xp25_ASAP7_75t_SL \i47/i131  (.A(\i47/n462 ),
    .B(\i47/n191 ),
    .C(\i47/n178 ),
    .D(\i47/n163 ),
    .Y(\i47/n300 ));
 AOI211xp5_ASAP7_75t_SL \i47/i132  (.A1(\i47/n59 ),
    .A2(\i47/n55 ),
    .B(\i47/n240 ),
    .C(\i47/n146 ),
    .Y(\i47/n299 ));
 AOI211xp5_ASAP7_75t_SL \i47/i133  (.A1(\i47/n97 ),
    .A2(\i47/n44 ),
    .B(\i47/n252 ),
    .C(\i47/n205 ),
    .Y(\i47/n298 ));
 NAND2xp33_ASAP7_75t_SL \i47/i134  (.A(\i47/n234 ),
    .B(\i47/n250 ),
    .Y(\i47/n297 ));
 NAND5xp2_ASAP7_75t_SL \i47/i135  (.A(\i47/n189 ),
    .B(\i47/n201 ),
    .C(\i47/n209 ),
    .D(\i47/n147 ),
    .E(\i47/n93 ),
    .Y(\i47/n296 ));
 NOR2xp33_ASAP7_75t_SL \i47/i136  (.A(\i47/n227 ),
    .B(\i47/n524 ),
    .Y(\i47/n295 ));
 OA21x2_ASAP7_75t_SL \i47/i137  (.A1(\i47/n492 ),
    .A2(\i47/n546 ),
    .B(\i47/n278 ),
    .Y(\i47/n294 ));
 NOR4xp25_ASAP7_75t_SL \i47/i138  (.A(\i47/n526 ),
    .B(\i47/n145 ),
    .C(\i47/n527 ),
    .D(\i47/n149 ),
    .Y(\i47/n293 ));
 NAND5xp2_ASAP7_75t_SL \i47/i139  (.A(\i47/n122 ),
    .B(\i47/n83 ),
    .C(\i47/n129 ),
    .D(\i47/n123 ),
    .E(\i47/n75 ),
    .Y(\i47/n292 ));
 NOR3xp33_ASAP7_75t_SL \i47/i14  (.A(\i47/n391 ),
    .B(\i47/n387 ),
    .C(\i47/n421 ),
    .Y(\i47/n417 ));
 NAND2xp5_ASAP7_75t_SL \i47/i140  (.A(\i47/n225 ),
    .B(\i47/n23 ),
    .Y(\i47/n291 ));
 NAND5xp2_ASAP7_75t_SL \i47/i141  (.A(\i47/n169 ),
    .B(\i47/n89 ),
    .C(\i47/n494 ),
    .D(\i47/n162 ),
    .E(\i47/n161 ),
    .Y(\i47/n290 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i47/i142  (.A1(\i47/n63 ),
    .A2(\i47/n79 ),
    .B(\i47/n433 ),
    .C(\i47/n218 ),
    .Y(\i47/n289 ));
 NAND4xp25_ASAP7_75t_SL \i47/i143  (.A(\i47/n549 ),
    .B(\i47/n509 ),
    .C(\i47/n482 ),
    .D(\i47/n534 ),
    .Y(\i47/n288 ));
 NAND5xp2_ASAP7_75t_SL \i47/i144  (.A(\i47/n558 ),
    .B(\i47/n535 ),
    .C(\i47/n195 ),
    .D(\i47/n515 ),
    .E(\i47/n87 ),
    .Y(\i47/n287 ));
 NAND2xp5_ASAP7_75t_SL \i47/i145  (.A(\i47/n224 ),
    .B(\i47/n550 ),
    .Y(\i47/n286 ));
 NAND2xp5_ASAP7_75t_SL \i47/i146  (.A(\i47/n183 ),
    .B(\i47/n277 ),
    .Y(\i47/n285 ));
 NOR2xp33_ASAP7_75t_L \i47/i147  (.A(\i47/n258 ),
    .B(\i47/n268 ),
    .Y(\i47/n303 ));
 NAND2xp5_ASAP7_75t_SL \i47/i148  (.A(\i47/n184 ),
    .B(\i47/n279 ),
    .Y(\i47/n284 ));
 NOR2x1p5_ASAP7_75t_SL \i47/i149  (.A(\i47/n464 ),
    .B(\i47/n260 ),
    .Y(\i47/n302 ));
 NOR2x2_ASAP7_75t_SL \i47/i15  (.A(\i47/n409 ),
    .B(\i47/n410 ),
    .Y(n26[2]));
 NAND3x1_ASAP7_75t_SL \i47/i150  (.A(\i47/n212 ),
    .B(\i47/n116 ),
    .C(\i47/n555 ),
    .Y(\i47/n25 ));
 INVxp67_ASAP7_75t_SL \i47/i151  (.A(\i47/n282 ),
    .Y(\i47/n283 ));
 INVxp67_ASAP7_75t_SL \i47/i152  (.A(\i47/n8 ),
    .Y(\i47/n281 ));
 INVxp67_ASAP7_75t_SL \i47/i153  (.A(\i47/n275 ),
    .Y(\i47/n276 ));
 INVxp67_ASAP7_75t_SL \i47/i154  (.A(\i47/n273 ),
    .Y(\i47/n274 ));
 INVx2_ASAP7_75t_SL \i47/i155  (.A(\i47/n271 ),
    .Y(\i47/n272 ));
 INVxp67_ASAP7_75t_SL \i47/i156  (.A(\i47/n269 ),
    .Y(\i47/n270 ));
 INVxp67_ASAP7_75t_SL \i47/i157  (.A(\i47/n266 ),
    .Y(\i47/n267 ));
 INVxp67_ASAP7_75t_SL \i47/i158  (.A(\i47/n475 ),
    .Y(\i47/n264 ));
 INVx1_ASAP7_75t_SL \i47/i159  (.A(\i47/n261 ),
    .Y(\i47/n262 ));
 NAND4xp75_ASAP7_75t_SL \i47/i16  (.A(\i47/n378 ),
    .B(\i47/n395 ),
    .C(\i47/n376 ),
    .D(\i47/n570 ),
    .Y(\i47/n416 ));
 NAND2x1_ASAP7_75t_SL \i47/i160  (.A(\i47/n506 ),
    .B(\i47/n177 ),
    .Y(\i47/n260 ));
 NAND2xp33_ASAP7_75t_SL \i47/i161  (.A(\i47/n495 ),
    .B(\i47/n545 ),
    .Y(\i47/n259 ));
 NAND2xp5_ASAP7_75t_SL \i47/i162  (.A(\i47/n148 ),
    .B(\i47/n495 ),
    .Y(\i47/n258 ));
 AOI31xp33_ASAP7_75t_SL \i47/i163  (.A1(\i47/n43 ),
    .A2(\i47/n16 ),
    .A3(\i47/n52 ),
    .B(\i47/n39 ),
    .Y(\i47/n257 ));
 NOR3xp33_ASAP7_75t_SL \i47/i164  (.A(\i47/n171 ),
    .B(\i47/n114 ),
    .C(\i47/n102 ),
    .Y(\i47/n256 ));
 NOR3xp33_ASAP7_75t_SL \i47/i165  (.A(\i47/n96 ),
    .B(\i47/n441 ),
    .C(\i47/n210 ),
    .Y(\i47/n255 ));
 AOI221xp5_ASAP7_75t_SL \i47/i166  (.A1(\i47/n63 ),
    .A2(\i47/n70 ),
    .B1(\i47/n46 ),
    .B2(\i47/n54 ),
    .C(\i47/n426 ),
    .Y(\i47/n254 ));
 AOI21xp5_ASAP7_75t_SL \i47/i167  (.A1(\i47/n135 ),
    .A2(\i47/n52 ),
    .B(\i47/n68 ),
    .Y(\i47/n282 ));
 OAI221xp5_ASAP7_75t_SL \i47/i168  (.A1(\i47/n17 ),
    .A2(\i47/n69 ),
    .B1(\i47/n507 ),
    .B2(\i47/n48 ),
    .C(\i47/n512 ),
    .Y(\i47/n253 ));
 AOI21xp33_ASAP7_75t_R \i47/i169  (.A1(\i47/n514 ),
    .A2(\i47/n40 ),
    .B(\i47/n62 ),
    .Y(\i47/n252 ));
 NOR3xp33_ASAP7_75t_SL \i47/i17  (.A(\i47/n420 ),
    .B(\i47/n362 ),
    .C(\i47/n403 ),
    .Y(\i47/n415 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i47/i170  (.A1(\i47/n430 ),
    .A2(\i47/n7 ),
    .B(\i47/n434 ),
    .C(\i47/n19 ),
    .Y(\i47/n251 ));
 NOR3xp33_ASAP7_75t_SL \i47/i171  (.A(\i47/n186 ),
    .B(\i47/n96 ),
    .C(\i47/n567 ),
    .Y(\i47/n250 ));
 NAND3xp33_ASAP7_75t_SL \i47/i172  (.A(\i47/n516 ),
    .B(\i47/n21 ),
    .C(\i47/n141 ),
    .Y(\i47/n249 ));
 AOI22xp5_ASAP7_75t_SL \i47/i173  (.A1(\i47/n50 ),
    .A2(\i47/n131 ),
    .B1(\i47/n54 ),
    .B2(\i47/n45 ),
    .Y(\i47/n248 ));
 NAND4xp25_ASAP7_75t_SL \i47/i174  (.A(\i47/n443 ),
    .B(\i47/n534 ),
    .C(\i47/n124 ),
    .D(\i47/n554 ),
    .Y(\i47/n247 ));
 NAND2xp33_ASAP7_75t_SL \i47/i175  (.A(\i47/n197 ),
    .B(\i47/n119 ),
    .Y(\i47/n246 ));
 OAI211xp5_ASAP7_75t_SL \i47/i176  (.A1(\i47/n56 ),
    .A2(\i47/n62 ),
    .B(\i47/n127 ),
    .C(\i47/n130 ),
    .Y(\i47/n280 ));
 NOR2xp67_ASAP7_75t_SL \i47/i177  (.A(\i47/n565 ),
    .B(\i47/n454 ),
    .Y(\i47/n279 ));
 AO21x1_ASAP7_75t_SL \i47/i178  (.A1(\i47/n47 ),
    .A2(\i47/n134 ),
    .B(\i47/n120 ),
    .Y(\i47/n278 ));
 AOI21x1_ASAP7_75t_SL \i47/i179  (.A1(\i47/n45 ),
    .A2(\i47/n559 ),
    .B(\i47/n564 ),
    .Y(\i47/n277 ));
 NAND4xp75_ASAP7_75t_SL \i47/i18  (.A(\i47/n377 ),
    .B(\i47/n405 ),
    .C(\i47/n381 ),
    .D(\i47/n372 ),
    .Y(\i47/n414 ));
 NAND2xp5_ASAP7_75t_SL \i47/i180  (.A(\i47/n552 ),
    .B(\i47/n553 ),
    .Y(\i47/n24 ));
 NOR2xp67_ASAP7_75t_SL \i47/i181  (.A(\i47/n526 ),
    .B(\i47/n199 ),
    .Y(\i47/n275 ));
 OAI211xp5_ASAP7_75t_SL \i47/i182  (.A1(\i47/n52 ),
    .A2(\i47/n62 ),
    .B(\i47/n159 ),
    .C(\i47/n160 ),
    .Y(\i47/n273 ));
 OR2x2_ASAP7_75t_SL \i47/i183  (.A(\i47/n563 ),
    .B(\i47/n528 ),
    .Y(\i47/n271 ));
 AOI21xp5_ASAP7_75t_SL \i47/i184  (.A1(\i47/n61 ),
    .A2(\i47/n53 ),
    .B(\i47/n455 ),
    .Y(\i47/n269 ));
 NAND2xp5_ASAP7_75t_SL \i47/i185  (.A(\i47/n537 ),
    .B(\i47/n538 ),
    .Y(\i47/n268 ));
 NAND2xp5_ASAP7_75t_SL \i47/i186  (.A(\i47/n22 ),
    .B(\i47/n166 ),
    .Y(\i47/n266 ));
 NAND2xp5_ASAP7_75t_SL \i47/i187  (.A(\i47/n196 ),
    .B(\i47/n215 ),
    .Y(\i47/n265 ));
 NAND2xp5_ASAP7_75t_SL \i47/i188  (.A(\i47/n153 ),
    .B(\i47/n511 ),
    .Y(\i47/n263 ));
 NOR2x1_ASAP7_75t_SL \i47/i189  (.A(\i47/n198 ),
    .B(\i47/n175 ),
    .Y(\i47/n261 ));
 AND3x4_ASAP7_75t_SL \i47/i19  (.A(\i47/n396 ),
    .B(\i47/n411 ),
    .C(\i47/n401 ),
    .Y(n26[7]));
 INVxp67_ASAP7_75t_SL \i47/i190  (.A(\i47/n243 ),
    .Y(\i47/n244 ));
 INVx1_ASAP7_75t_SL \i47/i191  (.A(\i47/n241 ),
    .Y(\i47/n242 ));
 INVx1_ASAP7_75t_SL \i47/i192  (.A(\i47/n237 ),
    .Y(\i47/n238 ));
 NAND4xp25_ASAP7_75t_SL \i47/i193  (.A(\i47/n499 ),
    .B(\i47/n110 ),
    .C(\i47/n517 ),
    .D(\i47/n498 ),
    .Y(\i47/n236 ));
 AOI31xp33_ASAP7_75t_SL \i47/i194  (.A1(\i47/n111 ),
    .A2(\i47/n546 ),
    .A3(\i47/n39 ),
    .B(\i47/n40 ),
    .Y(\i47/n235 ));
 NOR4xp25_ASAP7_75t_SL \i47/i195  (.A(\i47/n92 ),
    .B(\i47/n461 ),
    .C(\i47/n158 ),
    .D(\i47/n73 ),
    .Y(\i47/n234 ));
 AOI21xp5_ASAP7_75t_SL \i47/i196  (.A1(\i47/n533 ),
    .A2(\i47/n434 ),
    .B(\i47/n190 ),
    .Y(\i47/n233 ));
 NOR2xp33_ASAP7_75t_L \i47/i197  (.A(\i47/n165 ),
    .B(\i47/n207 ),
    .Y(\i47/n232 ));
 OAI31xp33_ASAP7_75t_SL \i47/i198  (.A1(\i47/n50 ),
    .A2(\i47/n46 ),
    .A3(\i47/n451 ),
    .B(\i47/n53 ),
    .Y(\i47/n231 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i47/i199  (.A1(\i47/n62 ),
    .A2(\i47/n42 ),
    .B(\i47/n67 ),
    .C(\i47/n187 ),
    .Y(\i47/n230 ));
 INVx2_ASAP7_75t_SL \i47/i2  (.A(n27[2]),
    .Y(\i47/n2 ));
 NAND4xp75_ASAP7_75t_SL \i47/i20  (.A(\i47/n361 ),
    .B(\i47/n380 ),
    .C(\i47/n389 ),
    .D(\i47/n404 ),
    .Y(\i47/n413 ));
 NOR2xp33_ASAP7_75t_SL \i47/i200  (.A(\i47/n523 ),
    .B(\i47/n568 ),
    .Y(\i47/n229 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i47/i201  (.A1(\i47/n50 ),
    .A2(\i47/n49 ),
    .B(\i47/n7 ),
    .C(\i47/n144 ),
    .Y(\i47/n228 ));
 NAND2xp33_ASAP7_75t_L \i47/i202  (.A(\i47/n501 ),
    .B(\i47/n491 ),
    .Y(\i47/n227 ));
 NAND2xp33_ASAP7_75t_SL \i47/i203  (.A(\i47/n204 ),
    .B(\i47/n108 ),
    .Y(\i47/n226 ));
 AOI22xp5_ASAP7_75t_SL \i47/i204  (.A1(\i47/n61 ),
    .A2(\i47/n90 ),
    .B1(\i47/n432 ),
    .B2(\i47/n63 ),
    .Y(\i47/n225 ));
 OAI21xp33_ASAP7_75t_SL \i47/i205  (.A1(\i47/n97 ),
    .A2(\i47/n61 ),
    .B(\i47/n432 ),
    .Y(\i47/n224 ));
 NAND2xp5_ASAP7_75t_SL \i47/i206  (.A(\i47/n536 ),
    .B(\i47/n214 ),
    .Y(\i47/n223 ));
 NAND4xp25_ASAP7_75t_SL \i47/i207  (.A(\i47/n106 ),
    .B(\i47/n126 ),
    .C(\i47/n88 ),
    .D(\i47/n86 ),
    .Y(\i47/n222 ));
 OAI222xp33_ASAP7_75t_SL \i47/i208  (.A1(\i47/n10 ),
    .A2(\i47/n43 ),
    .B1(\i47/n48 ),
    .B2(\i47/n56 ),
    .C1(\i47/n58 ),
    .C2(\i47/n64 ),
    .Y(\i47/n221 ));
 AND3x1_ASAP7_75t_SL \i47/i209  (.A(\i47/n104 ),
    .B(\i47/n110 ),
    .C(\i47/n192 ),
    .Y(\i47/n220 ));
 NAND2x1_ASAP7_75t_SL \i47/i21  (.A(\i47/n369 ),
    .B(\i47/n397 ),
    .Y(\i47/n412 ));
 AOI22xp5_ASAP7_75t_SL \i47/i210  (.A1(\i47/n467 ),
    .A2(\i47/n133 ),
    .B1(\i47/n559 ),
    .B2(\i47/n434 ),
    .Y(\i47/n245 ));
 AOI31xp33_ASAP7_75t_SL \i47/i211  (.A1(\i47/n43 ),
    .A2(\i47/n65 ),
    .A3(\i47/n481 ),
    .B(\i47/n47 ),
    .Y(\i47/n219 ));
 NAND2xp33_ASAP7_75t_SL \i47/i212  (.A(\i47/n505 ),
    .B(\i47/n193 ),
    .Y(\i47/n218 ));
 NAND3x1_ASAP7_75t_SL \i47/i213  (.A(\i47/n493 ),
    .B(\i47/n128 ),
    .C(\i47/n125 ),
    .Y(\i47/n243 ));
 AOI22x1_ASAP7_75t_SL \i47/i214  (.A1(\i47/n472 ),
    .A2(\i47/n451 ),
    .B1(\i47/n46 ),
    .B2(\i47/n57 ),
    .Y(\i47/n12 ));
 AOI221x1_ASAP7_75t_SL \i47/i215  (.A1(\i47/n451 ),
    .A2(\i47/n57 ),
    .B1(\i47/n63 ),
    .B2(\i47/n433 ),
    .C(\i47/n194 ),
    .Y(\i47/n241 ));
 AO21x2_ASAP7_75t_SL \i47/i216  (.A1(\i47/n432 ),
    .A2(\i47/n4 ),
    .B(\i47/n562 ),
    .Y(\i47/n240 ));
 OAI21xp5_ASAP7_75t_SL \i47/i217  (.A1(\i47/n39 ),
    .A2(\i47/n67 ),
    .B(\i47/n200 ),
    .Y(\i47/n239 ));
 NOR2x1_ASAP7_75t_SL \i47/i218  (.A(\i47/n105 ),
    .B(\i47/n561 ),
    .Y(\i47/n237 ));
 NOR2xp33_ASAP7_75t_L \i47/i219  (.A(\i47/n115 ),
    .B(\i47/n456 ),
    .Y(\i47/n23 ));
 NOR2xp67_ASAP7_75t_SL \i47/i22  (.A(\i47/n398 ),
    .B(\i47/n363 ),
    .Y(\i47/n411 ));
 NOR2xp33_ASAP7_75t_SL \i47/i220  (.A(\i47/n117 ),
    .B(\i47/n522 ),
    .Y(\i47/n217 ));
 INVx1_ASAP7_75t_SL \i47/i221  (.A(\i47/n215 ),
    .Y(\i47/n216 ));
 INVx1_ASAP7_75t_SL \i47/i222  (.A(\i47/n213 ),
    .Y(\i47/n214 ));
 INVx1_ASAP7_75t_SL \i47/i223  (.A(\i47/n522 ),
    .Y(\i47/n212 ));
 INVxp67_ASAP7_75t_SL \i47/i224  (.A(\i47/n538 ),
    .Y(\i47/n211 ));
 INVxp67_ASAP7_75t_SL \i47/i225  (.A(\i47/n455 ),
    .Y(\i47/n209 ));
 INVx1_ASAP7_75t_SL \i47/i226  (.A(\i47/n207 ),
    .Y(\i47/n208 ));
 NAND2xp5_ASAP7_75t_SL \i47/i227  (.A(\i47/n78 ),
    .B(\i47/n109 ),
    .Y(\i47/n205 ));
 OAI21xp5_ASAP7_75t_SL \i47/i228  (.A1(\i47/n46 ),
    .A2(\i47/n45 ),
    .B(\i47/n430 ),
    .Y(\i47/n204 ));
 NOR2xp33_ASAP7_75t_SL \i47/i229  (.A(\i47/n118 ),
    .B(\i47/n146 ),
    .Y(\i47/n203 ));
 NAND4xp75_ASAP7_75t_SL \i47/i23  (.A(\i47/n373 ),
    .B(\i47/n384 ),
    .C(\i47/n367 ),
    .D(\i47/n370 ),
    .Y(\i47/n410 ));
 NAND2xp33_ASAP7_75t_L \i47/i230  (.A(\i47/n143 ),
    .B(\i47/n82 ),
    .Y(\i47/n202 ));
 NOR2xp33_ASAP7_75t_SL \i47/i231  (.A(\i47/n19 ),
    .B(\i47/n99 ),
    .Y(\i47/n201 ));
 OAI21xp5_ASAP7_75t_SL \i47/i232  (.A1(\i47/n61 ),
    .A2(\i47/n66 ),
    .B(\i47/n54 ),
    .Y(\i47/n200 ));
 OAI21xp5_ASAP7_75t_SL \i47/i233  (.A1(\i47/n492 ),
    .A2(\i47/n68 ),
    .B(\i47/n540 ),
    .Y(\i47/n199 ));
 OAI21xp5_ASAP7_75t_SL \i47/i234  (.A1(\i47/n16 ),
    .A2(\i47/n58 ),
    .B(\i47/n113 ),
    .Y(\i47/n198 ));
 OAI21xp5_ASAP7_75t_SL \i47/i235  (.A1(\i47/n61 ),
    .A2(\i47/n45 ),
    .B(\i47/n55 ),
    .Y(\i47/n197 ));
 AOI22xp5_ASAP7_75t_SL \i47/i236  (.A1(\i47/n38 ),
    .A2(\i47/n70 ),
    .B1(\i47/n41 ),
    .B2(\i47/n61 ),
    .Y(\i47/n196 ));
 OAI21xp5_ASAP7_75t_SL \i47/i237  (.A1(\i47/n433 ),
    .A2(\i47/n70 ),
    .B(\i47/n467 ),
    .Y(\i47/n195 ));
 OA21x2_ASAP7_75t_SL \i47/i238  (.A1(\i47/n7 ),
    .A2(\i47/n70 ),
    .B(\i47/n434 ),
    .Y(\i47/n194 ));
 OAI21xp5_ASAP7_75t_SL \i47/i239  (.A1(\i47/n55 ),
    .A2(\i47/n41 ),
    .B(\i47/n467 ),
    .Y(\i47/n193 ));
 OR3x1_ASAP7_75t_SL \i47/i24  (.A(\i47/n392 ),
    .B(\i47/n390 ),
    .C(\i47/n374 ),
    .Y(\i47/n409 ));
 OAI21xp5_ASAP7_75t_SL \i47/i240  (.A1(\i47/n61 ),
    .A2(\i47/n59 ),
    .B(\i47/n70 ),
    .Y(\i47/n192 ));
 AOI21xp33_ASAP7_75t_SL \i47/i241  (.A1(\i47/n52 ),
    .A2(\i47/n67 ),
    .B(\i47/n39 ),
    .Y(\i47/n191 ));
 OAI21xp5_ASAP7_75t_SL \i47/i242  (.A1(\i47/n492 ),
    .A2(\i47/n58 ),
    .B(\i47/n557 ),
    .Y(\i47/n190 ));
 AOI22xp5_ASAP7_75t_SL \i47/i243  (.A1(\i47/n559 ),
    .A2(\i47/n50 ),
    .B1(\i47/n433 ),
    .B2(\i47/n49 ),
    .Y(\i47/n189 ));
 AOI21xp33_ASAP7_75t_SL \i47/i244  (.A1(\i47/n62 ),
    .A2(\i47/n39 ),
    .B(\i47/n481 ),
    .Y(\i47/n188 ));
 OAI21xp5_ASAP7_75t_SL \i47/i245  (.A1(\i47/n59 ),
    .A2(\i47/n50 ),
    .B(\i47/n433 ),
    .Y(\i47/n187 ));
 NAND2xp5_ASAP7_75t_SL \i47/i246  (.A(\i47/n467 ),
    .B(\i47/n533 ),
    .Y(\i47/n22 ));
 AOI22xp5_ASAP7_75t_SL \i47/i247  (.A1(\i47/n72 ),
    .A2(\i47/n518 ),
    .B1(\i47/n433 ),
    .B2(\i47/n4 ),
    .Y(\i47/n215 ));
 NAND2xp5_ASAP7_75t_L \i47/i248  (.A(\i47/n159 ),
    .B(\i47/n160 ),
    .Y(\i47/n186 ));
 OAI22xp5_ASAP7_75t_SL \i47/i249  (.A1(\i47/n71 ),
    .A2(\i47/n58 ),
    .B1(\i47/n17 ),
    .B2(\i47/n56 ),
    .Y(\i47/n213 ));
 OR3x1_ASAP7_75t_SL \i47/i25  (.A(\i47/n393 ),
    .B(\i47/n360 ),
    .C(\i47/n335 ),
    .Y(\i47/n408 ));
 NAND2xp5_ASAP7_75t_L \i47/i250  (.A(\i47/n18 ),
    .B(\i47/n132 ),
    .Y(\i47/n210 ));
 NOR2xp33_ASAP7_75t_L \i47/i251  (.A(\i47/n15 ),
    .B(\i47/n20 ),
    .Y(\i47/n207 ));
 NAND2xp33_ASAP7_75t_L \i47/i252  (.A(\i47/n482 ),
    .B(\i47/n483 ),
    .Y(\i47/n185 ));
 OAI21xp5_ASAP7_75t_SL \i47/i253  (.A1(\i47/n481 ),
    .A2(\i47/n48 ),
    .B(\i47/n93 ),
    .Y(\i47/n206 ));
 INVxp67_ASAP7_75t_SL \i47/i254  (.A(\i47/n181 ),
    .Y(\i47/n182 ));
 INVxp67_ASAP7_75t_SL \i47/i255  (.A(\i47/n179 ),
    .Y(\i47/n180 ));
 INVx1_ASAP7_75t_SL \i47/i256  (.A(\i47/n506 ),
    .Y(\i47/n178 ));
 INVx1_ASAP7_75t_SL \i47/i257  (.A(\i47/n457 ),
    .Y(\i47/n177 ));
 INVxp67_ASAP7_75t_SL \i47/i258  (.A(\i47/n512 ),
    .Y(\i47/n176 ));
 INVxp67_ASAP7_75t_SL \i47/i259  (.A(\i47/n523 ),
    .Y(\i47/n173 ));
 NAND3xp33_ASAP7_75t_SL \i47/i26  (.A(\i47/n402 ),
    .B(\i47/n389 ),
    .C(\i47/n373 ),
    .Y(\i47/n407 ));
 INVxp67_ASAP7_75t_SL \i47/i260  (.A(\i47/n529 ),
    .Y(\i47/n172 ));
 OAI21xp5_ASAP7_75t_SL \i47/i261  (.A1(\i47/n49 ),
    .A2(\i47/n518 ),
    .B(\i47/n433 ),
    .Y(\i47/n169 ));
 AO21x1_ASAP7_75t_SL \i47/i262  (.A1(\i47/n38 ),
    .A2(\i47/n57 ),
    .B(\i47/n98 ),
    .Y(\i47/n168 ));
 AOI22xp5_ASAP7_75t_SL \i47/i263  (.A1(\i47/n72 ),
    .A2(\i47/n467 ),
    .B1(\i47/n430 ),
    .B2(\i47/n45 ),
    .Y(\i47/n184 ));
 OAI22xp5_ASAP7_75t_SL \i47/i264  (.A1(\i47/n52 ),
    .A2(\i47/n10 ),
    .B1(\i47/n67 ),
    .B2(\i47/n62 ),
    .Y(\i47/n167 ));
 AOI22xp5_ASAP7_75t_SL \i47/i265  (.A1(\i47/n38 ),
    .A2(\i47/n41 ),
    .B1(\i47/n72 ),
    .B2(\i47/n61 ),
    .Y(\i47/n183 ));
 AOI22xp5_ASAP7_75t_SL \i47/i266  (.A1(\i47/n54 ),
    .A2(\i47/n518 ),
    .B1(\i47/n41 ),
    .B2(\i47/n66 ),
    .Y(\i47/n166 ));
 OAI21xp5_ASAP7_75t_SL \i47/i267  (.A1(\i47/n64 ),
    .A2(\i47/n47 ),
    .B(\i47/n108 ),
    .Y(\i47/n165 ));
 OAI21xp5_ASAP7_75t_SL \i47/i268  (.A1(\i47/n40 ),
    .A2(\i47/n48 ),
    .B(\i47/n100 ),
    .Y(\i47/n181 ));
 AOI22xp5_ASAP7_75t_SL \i47/i269  (.A1(\i47/n38 ),
    .A2(\i47/n55 ),
    .B1(\i47/n41 ),
    .B2(\i47/n45 ),
    .Y(\i47/n179 ));
 NOR2x1_ASAP7_75t_SL \i47/i27  (.A(\i47/n316 ),
    .B(\i47/n390 ),
    .Y(\i47/n405 ));
 OA21x2_ASAP7_75t_SL \i47/i270  (.A1(\i47/n43 ),
    .A2(\i47/n47 ),
    .B(\i47/n496 ),
    .Y(\i47/n164 ));
 NAND2xp33_ASAP7_75t_SL \i47/i271  (.A(\i47/n161 ),
    .B(\i47/n162 ),
    .Y(\i47/n163 ));
 AO22x2_ASAP7_75t_SL \i47/i272  (.A1(\i47/n70 ),
    .A2(\i47/n451 ),
    .B1(\i47/n44 ),
    .B2(\i47/n66 ),
    .Y(\i47/n175 ));
 OAI21xp5_ASAP7_75t_SL \i47/i273  (.A1(\i47/n64 ),
    .A2(\i47/n42 ),
    .B(\i47/n497 ),
    .Y(\i47/n174 ));
 OAI22xp5_ASAP7_75t_SL \i47/i274  (.A1(\i47/n43 ),
    .A2(\i47/n51 ),
    .B1(\i47/n56 ),
    .B2(\i47/n60 ),
    .Y(\i47/n171 ));
 OAI22xp5_ASAP7_75t_SL \i47/i275  (.A1(\i47/n43 ),
    .A2(\i47/n42 ),
    .B1(\i47/n47 ),
    .B2(\i47/n507 ),
    .Y(\i47/n170 ));
 INVxp67_ASAP7_75t_SL \i47/i276  (.A(\i47/n156 ),
    .Y(\i47/n157 ));
 INVx1_ASAP7_75t_SL \i47/i277  (.A(\i47/n556 ),
    .Y(\i47/n155 ));
 INVxp67_ASAP7_75t_SL \i47/i278  (.A(\i47/n153 ),
    .Y(\i47/n154 ));
 INVxp67_ASAP7_75t_SL \i47/i279  (.A(\i47/n443 ),
    .Y(\i47/n152 ));
 NOR2x1_ASAP7_75t_SL \i47/i28  (.A(\i47/n375 ),
    .B(\i47/n371 ),
    .Y(\i47/n404 ));
 INVxp67_ASAP7_75t_SL \i47/i280  (.A(\i47/n150 ),
    .Y(\i47/n151 ));
 INVxp33_ASAP7_75t_SL \i47/i281  (.A(\i47/n480 ),
    .Y(\i47/n148 ));
 INVxp67_ASAP7_75t_SL \i47/i282  (.A(\i47/n540 ),
    .Y(\i47/n145 ));
 INVxp67_ASAP7_75t_SL \i47/i283  (.A(\i47/n143 ),
    .Y(\i47/n144 ));
 INVxp67_ASAP7_75t_SL \i47/i284  (.A(\i47/n141 ),
    .Y(\i47/n142 ));
 INVxp67_ASAP7_75t_SL \i47/i285  (.A(\i47/n139 ),
    .Y(\i47/n140 ));
 INVxp67_ASAP7_75t_SL \i47/i286  (.A(\i47/n137 ),
    .Y(\i47/n138 ));
 INVxp67_ASAP7_75t_SL \i47/i287  (.A(\i47/n20 ),
    .Y(\i47/n136 ));
 INVx2_ASAP7_75t_SL \i47/i288  (.A(\i47/n533 ),
    .Y(\i47/n135 ));
 NAND2xp5_ASAP7_75t_SL \i47/i289  (.A(\i47/n55 ),
    .B(\i47/n467 ),
    .Y(\i47/n162 ));
 NAND3xp33_ASAP7_75t_SL \i47/i29  (.A(\i47/n355 ),
    .B(\i47/n579 ),
    .C(\i47/n352 ),
    .Y(\i47/n403 ));
 NAND2xp5_ASAP7_75t_SL \i47/i290  (.A(\i47/n430 ),
    .B(\i47/n66 ),
    .Y(\i47/n134 ));
 NAND2xp5_ASAP7_75t_SL \i47/i291  (.A(\i47/n67 ),
    .B(\i47/n65 ),
    .Y(\i47/n133 ));
 NAND2xp5_ASAP7_75t_SL \i47/i292  (.A(\i47/n41 ),
    .B(\i47/n451 ),
    .Y(\i47/n132 ));
 NAND2xp33_ASAP7_75t_SL \i47/i293  (.A(\i47/n52 ),
    .B(\i47/n492 ),
    .Y(\i47/n131 ));
 NAND2xp5_ASAP7_75t_SL \i47/i294  (.A(\i47/n49 ),
    .B(\i47/n559 ),
    .Y(\i47/n130 ));
 NAND2xp5_ASAP7_75t_SL \i47/i295  (.A(\i47/n49 ),
    .B(\i47/n54 ),
    .Y(\i47/n161 ));
 NAND2xp5_ASAP7_75t_SL \i47/i296  (.A(\i47/n559 ),
    .B(\i47/n59 ),
    .Y(\i47/n160 ));
 NAND2xp5_ASAP7_75t_SL \i47/i297  (.A(\i47/n54 ),
    .B(\i47/n467 ),
    .Y(\i47/n129 ));
 NAND2xp5_ASAP7_75t_SL \i47/i298  (.A(\i47/n4 ),
    .B(\i47/n559 ),
    .Y(\i47/n128 ));
 NAND2xp5_ASAP7_75t_SL \i47/i299  (.A(\i47/n430 ),
    .B(\i47/n434 ),
    .Y(\i47/n127 ));
 INVx2_ASAP7_75t_SL \i47/i3  (.A(n27[0]),
    .Y(\i47/n3 ));
 NOR2xp33_ASAP7_75t_SL \i47/i30  (.A(\i47/n379 ),
    .B(\i47/n489 ),
    .Y(\i47/n402 ));
 NAND2xp5_ASAP7_75t_SL \i47/i300  (.A(\i47/n55 ),
    .B(\i47/n4 ),
    .Y(\i47/n126 ));
 NAND2xp67_ASAP7_75t_SL \i47/i301  (.A(\i47/n38 ),
    .B(\i47/n44 ),
    .Y(\i47/n125 ));
 NAND2xp5_ASAP7_75t_SL \i47/i302  (.A(\i47/n44 ),
    .B(\i47/n59 ),
    .Y(\i47/n124 ));
 NAND2xp5_ASAP7_75t_SL \i47/i303  (.A(\i47/n55 ),
    .B(\i47/n434 ),
    .Y(\i47/n123 ));
 NAND2xp5_ASAP7_75t_SL \i47/i304  (.A(\i47/n38 ),
    .B(\i47/n433 ),
    .Y(\i47/n159 ));
 AND2x2_ASAP7_75t_SL \i47/i305  (.A(\i47/n44 ),
    .B(\i47/n61 ),
    .Y(\i47/n158 ));
 AND2x2_ASAP7_75t_SL \i47/i306  (.A(\i47/n430 ),
    .B(\i47/n59 ),
    .Y(\i47/n156 ));
 NAND2xp5_ASAP7_75t_SL \i47/i307  (.A(\i47/n433 ),
    .B(\i47/n434 ),
    .Y(\i47/n153 ));
 NAND2xp5_ASAP7_75t_SL \i47/i308  (.A(\i47/n53 ),
    .B(\i47/n59 ),
    .Y(\i47/n150 ));
 AND2x2_ASAP7_75t_SL \i47/i309  (.A(\i47/n55 ),
    .B(\i47/n50 ),
    .Y(\i47/n149 ));
 NOR5xp2_ASAP7_75t_SL \i47/i31  (.A(\i47/n345 ),
    .B(\i47/n296 ),
    .C(\i47/n337 ),
    .D(\i47/n265 ),
    .E(\i47/n525 ),
    .Y(\i47/n401 ));
 NAND2xp5_ASAP7_75t_SL \i47/i310  (.A(\i47/n53 ),
    .B(\i47/n49 ),
    .Y(\i47/n147 ));
 NAND2xp5_ASAP7_75t_SL \i47/i311  (.A(\i47/n50 ),
    .B(\i47/n559 ),
    .Y(\i47/n122 ));
 AND2x2_ASAP7_75t_SL \i47/i312  (.A(\i47/n54 ),
    .B(\i47/n4 ),
    .Y(\i47/n146 ));
 NOR2xp33_ASAP7_75t_L \i47/i313  (.A(\i47/n16 ),
    .B(\i47/n15 ),
    .Y(\i47/n121 ));
 NOR2xp33_ASAP7_75t_SL \i47/i314  (.A(\i47/n53 ),
    .B(\i47/n430 ),
    .Y(\i47/n120 ));
 NAND2xp5_ASAP7_75t_SL \i47/i315  (.A(\i47/n430 ),
    .B(\i47/n4 ),
    .Y(\i47/n143 ));
 NAND2xp5_ASAP7_75t_SL \i47/i316  (.A(\i47/n53 ),
    .B(\i47/n518 ),
    .Y(\i47/n21 ));
 NAND2xp5_ASAP7_75t_SL \i47/i317  (.A(\i47/n70 ),
    .B(\i47/n45 ),
    .Y(\i47/n141 ));
 NAND2xp5_ASAP7_75t_SL \i47/i318  (.A(\i47/n434 ),
    .B(\i47/n54 ),
    .Y(\i47/n139 ));
 NAND2xp5_ASAP7_75t_SL \i47/i319  (.A(\i47/n55 ),
    .B(\i47/n63 ),
    .Y(\i47/n119 ));
 NOR3xp33_ASAP7_75t_SL \i47/i32  (.A(\i47/n342 ),
    .B(\i47/n357 ),
    .C(\i47/n388 ),
    .Y(\i47/n400 ));
 NOR2xp33_ASAP7_75t_SL \i47/i320  (.A(\i47/n430 ),
    .B(\i47/n55 ),
    .Y(\i47/n137 ));
 NOR2xp33_ASAP7_75t_SL \i47/i321  (.A(\i47/n48 ),
    .B(\i47/n67 ),
    .Y(\i47/n118 ));
 NOR2x1_ASAP7_75t_SL \i47/i322  (.A(\i47/n53 ),
    .B(\i47/n432 ),
    .Y(\i47/n20 ));
 INVxp67_ASAP7_75t_SL \i47/i323  (.A(\i47/n116 ),
    .Y(\i47/n117 ));
 INVxp67_ASAP7_75t_SL \i47/i324  (.A(\i47/n113 ),
    .Y(\i47/n114 ));
 INVx1_ASAP7_75t_SL \i47/i325  (.A(\i47/n111 ),
    .Y(\i47/n112 ));
 INVxp67_ASAP7_75t_SL \i47/i326  (.A(\i47/n106 ),
    .Y(\i47/n107 ));
 INVxp67_ASAP7_75t_SL \i47/i327  (.A(\i47/n445 ),
    .Y(\i47/n105 ));
 INVxp67_ASAP7_75t_SL \i47/i328  (.A(\i47/n461 ),
    .Y(\i47/n104 ));
 INVxp67_ASAP7_75t_SL \i47/i329  (.A(\i47/n442 ),
    .Y(\i47/n103 ));
 NOR2x1_ASAP7_75t_SL \i47/i33  (.A(\i47/n385 ),
    .B(\i47/n346 ),
    .Y(\i47/n399 ));
 INVxp67_ASAP7_75t_SL \i47/i330  (.A(\i47/n101 ),
    .Y(\i47/n102 ));
 INVxp67_ASAP7_75t_SL \i47/i331  (.A(\i47/n99 ),
    .Y(\i47/n100 ));
 INVxp67_ASAP7_75t_SL \i47/i332  (.A(\i47/n499 ),
    .Y(\i47/n94 ));
 INVx1_ASAP7_75t_SL \i47/i333  (.A(\i47/n501 ),
    .Y(\i47/n92 ));
 INVx1_ASAP7_75t_SL \i47/i334  (.A(\i47/n18 ),
    .Y(\i47/n19 ));
 NAND2xp5_ASAP7_75t_SL \i47/i335  (.A(\i47/n432 ),
    .B(\i47/n61 ),
    .Y(\i47/n91 ));
 NAND2xp5_ASAP7_75t_SL \i47/i336  (.A(\i47/n64 ),
    .B(\i47/n481 ),
    .Y(\i47/n90 ));
 NAND2xp5_ASAP7_75t_SL \i47/i337  (.A(\i47/n63 ),
    .B(\i47/n41 ),
    .Y(\i47/n89 ));
 NAND2xp5_ASAP7_75t_SL \i47/i338  (.A(\i47/n433 ),
    .B(\i47/n50 ),
    .Y(\i47/n88 ));
 NAND2xp5_ASAP7_75t_SL \i47/i339  (.A(\i47/n57 ),
    .B(\i47/n45 ),
    .Y(\i47/n87 ));
 NAND2xp5_ASAP7_75t_SL \i47/i34  (.A(\i47/n344 ),
    .B(\i47/n364 ),
    .Y(\i47/n398 ));
 NAND2xp5_ASAP7_75t_SL \i47/i340  (.A(\i47/n41 ),
    .B(\i47/n59 ),
    .Y(\i47/n86 ));
 NAND2xp5_ASAP7_75t_L \i47/i341  (.A(\i47/n17 ),
    .B(\i47/n39 ),
    .Y(\i47/n85 ));
 NAND2xp33_ASAP7_75t_SL \i47/i342  (.A(\i47/n51 ),
    .B(\i47/n10 ),
    .Y(\i47/n84 ));
 NAND2xp5_ASAP7_75t_SL \i47/i343  (.A(\i47/n7 ),
    .B(\i47/n49 ),
    .Y(\i47/n83 ));
 NAND2xp5_ASAP7_75t_SL \i47/i344  (.A(\i47/n72 ),
    .B(\i47/n46 ),
    .Y(\i47/n116 ));
 NAND2xp5_ASAP7_75t_SL \i47/i345  (.A(\i47/n432 ),
    .B(\i47/n49 ),
    .Y(\i47/n82 ));
 NOR2xp33_ASAP7_75t_SL \i47/i346  (.A(\i47/n48 ),
    .B(\i47/n492 ),
    .Y(\i47/n81 ));
 AND2x2_ASAP7_75t_SL \i47/i347  (.A(\i47/n7 ),
    .B(\i47/n63 ),
    .Y(\i47/n115 ));
 NAND2xp5_ASAP7_75t_SL \i47/i348  (.A(\i47/n430 ),
    .B(\i47/n50 ),
    .Y(\i47/n113 ));
 NOR2x1_ASAP7_75t_SL \i47/i349  (.A(\i47/n59 ),
    .B(\i47/n66 ),
    .Y(\i47/n111 ));
 NOR3x1_ASAP7_75t_SL \i47/i35  (.A(\i47/n25 ),
    .B(\i47/n359 ),
    .C(\i47/n291 ),
    .Y(\i47/n406 ));
 NAND2xp5_ASAP7_75t_SL \i47/i350  (.A(\i47/n7 ),
    .B(\i47/n518 ),
    .Y(\i47/n110 ));
 NAND2xp5_ASAP7_75t_SL \i47/i351  (.A(\i47/n433 ),
    .B(\i47/n45 ),
    .Y(\i47/n109 ));
 NAND2xp5_ASAP7_75t_SL \i47/i352  (.A(\i47/n44 ),
    .B(\i47/n49 ),
    .Y(\i47/n108 ));
 NOR2xp33_ASAP7_75t_SL \i47/i353  (.A(\i47/n59 ),
    .B(\i47/n49 ),
    .Y(\i47/n80 ));
 NAND2xp5_ASAP7_75t_SL \i47/i354  (.A(\i47/n432 ),
    .B(\i47/n434 ),
    .Y(\i47/n106 ));
 NAND2xp33_ASAP7_75t_L \i47/i355  (.A(\i47/n42 ),
    .B(\i47/n60 ),
    .Y(\i47/n79 ));
 NAND2xp5_ASAP7_75t_SL \i47/i356  (.A(\i47/n38 ),
    .B(\i47/n72 ),
    .Y(\i47/n101 ));
 NOR2xp67_ASAP7_75t_R \i47/i357  (.A(\i47/n39 ),
    .B(\i47/n492 ),
    .Y(\i47/n99 ));
 AND2x2_ASAP7_75t_SL \i47/i358  (.A(\i47/n72 ),
    .B(\i47/n66 ),
    .Y(\i47/n98 ));
 NAND2xp5_ASAP7_75t_L \i47/i359  (.A(\i47/n15 ),
    .B(\i47/n17 ),
    .Y(\i47/n97 ));
 NOR3xp33_ASAP7_75t_SL \i47/i36  (.A(\i47/n382 ),
    .B(\i47/n25 ),
    .C(\i47/n305 ),
    .Y(\i47/n396 ));
 NAND2xp33_ASAP7_75t_L \i47/i360  (.A(\i47/n4 ),
    .B(\i47/n433 ),
    .Y(\i47/n78 ));
 AND2x2_ASAP7_75t_SL \i47/i361  (.A(\i47/n72 ),
    .B(\i47/n50 ),
    .Y(\i47/n96 ));
 NOR2xp33_ASAP7_75t_SL \i47/i362  (.A(\i47/n51 ),
    .B(\i47/n40 ),
    .Y(\i47/n77 ));
 NOR2xp33_ASAP7_75t_SL \i47/i363  (.A(\i47/n47 ),
    .B(\i47/n507 ),
    .Y(\i47/n76 ));
 NOR2xp67_ASAP7_75t_SL \i47/i364  (.A(\i47/n46 ),
    .B(\i47/n61 ),
    .Y(\i47/n95 ));
 NAND2xp5_ASAP7_75t_SL \i47/i365  (.A(\i47/n7 ),
    .B(\i47/n66 ),
    .Y(\i47/n75 ));
 NAND2xp5_ASAP7_75t_SL \i47/i366  (.A(\i47/n72 ),
    .B(\i47/n63 ),
    .Y(\i47/n93 ));
 NOR2xp33_ASAP7_75t_SL \i47/i367  (.A(\i47/n71 ),
    .B(\i47/n15 ),
    .Y(\i47/n74 ));
 NOR2xp33_ASAP7_75t_SL \i47/i368  (.A(\i47/n71 ),
    .B(\i47/n48 ),
    .Y(\i47/n73 ));
 NAND2xp5_ASAP7_75t_SL \i47/i369  (.A(\i47/n7 ),
    .B(\i47/n45 ),
    .Y(\i47/n18 ));
 NOR2xp67_ASAP7_75t_SL \i47/i37  (.A(\i47/n365 ),
    .B(\i47/n25 ),
    .Y(\i47/n395 ));
 INVx2_ASAP7_75t_SL \i47/i370  (.A(\i47/n72 ),
    .Y(\i47/n71 ));
 INVx1_ASAP7_75t_SL \i47/i371  (.A(\i47/n70 ),
    .Y(\i47/n69 ));
 INVx3_ASAP7_75t_SL \i47/i372  (.A(\i47/n434 ),
    .Y(\i47/n68 ));
 INVx2_ASAP7_75t_SL \i47/i373  (.A(\i47/n430 ),
    .Y(\i47/n67 ));
 INVx2_ASAP7_75t_SL \i47/i374  (.A(\i47/n432 ),
    .Y(\i47/n65 ));
 INVx2_ASAP7_75t_SL \i47/i375  (.A(\i47/n433 ),
    .Y(\i47/n64 ));
 INVx3_ASAP7_75t_SL \i47/i376  (.A(\i47/n63 ),
    .Y(\i47/n62 ));
 INVx2_ASAP7_75t_SL \i47/i377  (.A(\i47/n61 ),
    .Y(\i47/n60 ));
 INVx3_ASAP7_75t_SL \i47/i378  (.A(\i47/n59 ),
    .Y(\i47/n58 ));
 INVx3_ASAP7_75t_SL \i47/i379  (.A(\i47/n56 ),
    .Y(\i47/n55 ));
 NOR3xp33_ASAP7_75t_SL \i47/i38  (.A(\i47/n343 ),
    .B(\i47/n338 ),
    .C(\i47/n9 ),
    .Y(\i47/n394 ));
 AND2x4_ASAP7_75t_SL \i47/i380  (.A(\i47/n34 ),
    .B(\i47/n6 ),
    .Y(\i47/n72 ));
 AND2x4_ASAP7_75t_SL \i47/i381  (.A(\i47/n530 ),
    .B(\i47/n34 ),
    .Y(\i47/n70 ));
 AND2x4_ASAP7_75t_SL \i47/i382  (.A(\i47/n542 ),
    .B(\i47/n438 ),
    .Y(\i47/n66 ));
 NAND2x1_ASAP7_75t_SL \i47/i383  (.A(\i47/n542 ),
    .B(\i47/n438 ),
    .Y(\i47/n17 ));
 AND2x4_ASAP7_75t_SL \i47/i384  (.A(\i47/n542 ),
    .B(\i47/n32 ),
    .Y(\i47/n63 ));
 AND2x4_ASAP7_75t_SL \i47/i385  (.A(\i47/n541 ),
    .B(\i47/n14 ),
    .Y(\i47/n61 ));
 AND2x4_ASAP7_75t_SL \i47/i386  (.A(\i47/n542 ),
    .B(\i47/n31 ),
    .Y(\i47/n59 ));
 AND2x4_ASAP7_75t_SL \i47/i387  (.A(\i47/n530 ),
    .B(\i47/n503 ),
    .Y(\i47/n57 ));
 OR2x6_ASAP7_75t_SL \i47/i388  (.A(\i47/n35 ),
    .B(\i47/n429 ),
    .Y(\i47/n56 ));
 INVx3_ASAP7_75t_SL \i47/i389  (.A(\i47/n54 ),
    .Y(\i47/n16 ));
 NAND3xp33_ASAP7_75t_SL \i47/i39  (.A(\i47/n486 ),
    .B(\i47/n351 ),
    .C(\i47/n339 ),
    .Y(\i47/n393 ));
 INVx3_ASAP7_75t_SL \i47/i390  (.A(\i47/n53 ),
    .Y(\i47/n52 ));
 INVx4_ASAP7_75t_SL \i47/i391  (.A(\i47/n51 ),
    .Y(\i47/n50 ));
 INVx2_ASAP7_75t_SL \i47/i392  (.A(\i47/n49 ),
    .Y(\i47/n48 ));
 INVx4_ASAP7_75t_SL \i47/i393  (.A(\i47/n47 ),
    .Y(\i47/n46 ));
 INVx4_ASAP7_75t_SL \i47/i394  (.A(\i47/n45 ),
    .Y(\i47/n15 ));
 INVx4_ASAP7_75t_SL \i47/i395  (.A(\i47/n44 ),
    .Y(\i47/n43 ));
 INVx3_ASAP7_75t_SL \i47/i396  (.A(\i47/n41 ),
    .Y(\i47/n40 ));
 INVx3_ASAP7_75t_SL \i47/i397  (.A(\i47/n39 ),
    .Y(\i47/n38 ));
 AND2x4_ASAP7_75t_SL \i47/i398  (.A(\i47/n34 ),
    .B(\i47/n36 ),
    .Y(\i47/n54 ));
 AND2x4_ASAP7_75t_SL \i47/i399  (.A(\i47/n6 ),
    .B(\i47/n503 ),
    .Y(\i47/n53 ));
 INVx2_ASAP7_75t_SL \i47/i4  (.A(\i47/n10 ),
    .Y(\i47/n4 ));
 NAND2xp5_ASAP7_75t_L \i47/i40  (.A(\i47/n571 ),
    .B(\i47/n383 ),
    .Y(\i47/n392 ));
 NAND2x1p5_ASAP7_75t_SL \i47/i400  (.A(\i47/n541 ),
    .B(\i47/n37 ),
    .Y(\i47/n51 ));
 NAND2x1p5_ASAP7_75t_SL \i47/i401  (.A(\i47/n5 ),
    .B(\i47/n32 ),
    .Y(\i47/n10 ));
 AND2x4_ASAP7_75t_SL \i47/i402  (.A(\i47/n32 ),
    .B(\i47/n14 ),
    .Y(\i47/n49 ));
 OR2x4_ASAP7_75t_SL \i47/i403  (.A(\i47/n29 ),
    .B(\i47/n30 ),
    .Y(\i47/n47 ));
 AND2x4_ASAP7_75t_SL \i47/i404  (.A(\i47/n31 ),
    .B(\i47/n14 ),
    .Y(\i47/n45 ));
 AND2x4_ASAP7_75t_SL \i47/i405  (.A(\i47/n6 ),
    .B(\i47/n531 ),
    .Y(\i47/n44 ));
 NAND2x1_ASAP7_75t_SL \i47/i406  (.A(\i47/n5 ),
    .B(\i47/n438 ),
    .Y(\i47/n42 ));
 AND2x4_ASAP7_75t_SL \i47/i407  (.A(\i47/n36 ),
    .B(\i47/n503 ),
    .Y(\i47/n41 ));
 OR2x6_ASAP7_75t_SL \i47/i408  (.A(\i47/n28 ),
    .B(\i47/n33 ),
    .Y(\i47/n39 ));
 INVx2_ASAP7_75t_SL \i47/i409  (.A(\i47/n468 ),
    .Y(\i47/n36 ));
 NAND2xp33_ASAP7_75t_SL \i47/i41  (.A(\i47/n574 ),
    .B(\i47/n366 ),
    .Y(\i47/n391 ));
 NAND2xp5_ASAP7_75t_SL \i47/i410  (.A(\i47/n11 ),
    .B(\i47/n2 ),
    .Y(\i47/n33 ));
 AND2x2_ASAP7_75t_SL \i47/i411  (.A(\i47/n11 ),
    .B(\i47/n2 ),
    .Y(\i47/n37 ));
 NAND2x1p5_ASAP7_75t_SL \i47/i412  (.A(n27[5]),
    .B(n27[4]),
    .Y(\i47/n35 ));
 AND2x2_ASAP7_75t_SL \i47/i413  (.A(\i47/n0 ),
    .B(\i47/n13 ),
    .Y(\i47/n34 ));
 INVx2_ASAP7_75t_SL \i47/i414  (.A(\i47/n30 ),
    .Y(\i47/n31 ));
 NAND2xp5_ASAP7_75t_SL \i47/i415  (.A(\i47/n27 ),
    .B(\i47/n3 ),
    .Y(\i47/n28 ));
 AND2x4_ASAP7_75t_SL \i47/i416  (.A(n27[0]),
    .B(\i47/n27 ),
    .Y(\i47/n32 ));
 NAND2xp5_ASAP7_75t_SL \i47/i417  (.A(\i47/n3 ),
    .B(n27[1]),
    .Y(\i47/n30 ));
 OR2x2_ASAP7_75t_SL \i47/i418  (.A(\i47/n2 ),
    .B(n27[3]),
    .Y(\i47/n29 ));
 INVx1_ASAP7_75t_SL \i47/i419  (.A(n27[1]),
    .Y(\i47/n27 ));
 NOR2x1_ASAP7_75t_SL \i47/i42  (.A(\i47/n422 ),
    .B(\i47/n374 ),
    .Y(\i47/n397 ));
 INVx4_ASAP7_75t_SL \i47/i420  (.A(n27[5]),
    .Y(\i47/n26 ));
 INVx2_ASAP7_75t_SL \i47/i421  (.A(\i47/n448 ),
    .Y(\i47/n14 ));
 INVx2_ASAP7_75t_SL \i47/i422  (.A(n27[6]),
    .Y(\i47/n13 ));
 INVx2_ASAP7_75t_SL \i47/i423  (.A(n27[3]),
    .Y(\i47/n11 ));
 INVxp67_ASAP7_75t_SL \i47/i424  (.A(\i47/n351 ),
    .Y(\i47/n9 ));
 OR2x2_ASAP7_75t_SL \i47/i425  (.A(\i47/n441 ),
    .B(\i47/n528 ),
    .Y(\i47/n8 ));
 OAI221xp5_ASAP7_75t_SL \i47/i426  (.A1(\i47/n492 ),
    .A2(\i47/n42 ),
    .B1(\i47/n47 ),
    .B2(\i47/n40 ),
    .C(\i47/n101 ),
    .Y(\i47/n418 ));
 NAND4xp25_ASAP7_75t_SL \i47/i427  (.A(\i47/n325 ),
    .B(\i47/n419 ),
    .C(\i47/n319 ),
    .D(\i47/n350 ),
    .Y(\i47/n420 ));
 NOR2x1_ASAP7_75t_SL \i47/i428  (.A(\i47/n520 ),
    .B(\i47/n418 ),
    .Y(\i47/n419 ));
 NAND3xp33_ASAP7_75t_L \i47/i429  (.A(\i47/n303 ),
    .B(\i47/n419 ),
    .C(\i47/n368 ),
    .Y(\i47/n421 ));
 NAND2xp33_ASAP7_75t_L \i47/i43  (.A(\i47/n354 ),
    .B(\i47/n327 ),
    .Y(\i47/n388 ));
 NAND4xp25_ASAP7_75t_SL \i47/i430  (.A(\i47/n312 ),
    .B(\i47/n419 ),
    .C(\i47/n324 ),
    .D(\i47/n308 ),
    .Y(\i47/n422 ));
 AOI211xp5_ASAP7_75t_SL \i47/i431  (.A1(\i47/n112 ),
    .A2(\i47/n432 ),
    .B(\i47/n424 ),
    .C(\i47/n81 ),
    .Y(\i47/n423 ));
 NOR3xp33_ASAP7_75t_SL \i47/i432  (.A(\i47/n239 ),
    .B(\i47/n424 ),
    .C(\i47/n74 ),
    .Y(\i47/n425 ));
 OAI22xp5_ASAP7_75t_SL \i47/i433  (.A1(\i47/n39 ),
    .A2(\i47/n470 ),
    .B1(\i47/n560 ),
    .B2(\i47/n546 ),
    .Y(\i47/n426 ));
 OAI221xp5_ASAP7_75t_SL \i47/i434  (.A1(\i47/n460 ),
    .A2(\i47/n64 ),
    .B1(\i47/n58 ),
    .B2(\i47/n481 ),
    .C(\i47/n173 ),
    .Y(\i47/n427 ));
 INVx1_ASAP7_75t_SL \i47/i435  (.A(\i47/n428 ),
    .Y(\i47/n429 ));
 AND2x4_ASAP7_75t_SL \i47/i436  (.A(n27[7]),
    .B(n27[6]),
    .Y(\i47/n428 ));
 AND2x4_ASAP7_75t_SL \i47/i437  (.A(\i47/n428 ),
    .B(\i47/n36 ),
    .Y(\i47/n430 ));
 AOI211xp5_ASAP7_75t_SL \i47/i438  (.A1(\i47/n451 ),
    .A2(\i47/n428 ),
    .B(\i47/n98 ),
    .C(\i47/n103 ),
    .Y(\i47/n431 ));
 AND2x4_ASAP7_75t_SL \i47/i439  (.A(\i47/n428 ),
    .B(\i47/n530 ),
    .Y(\i47/n432 ));
 NAND2xp33_ASAP7_75t_L \i47/i44  (.A(\i47/n571 ),
    .B(\i47/n333 ),
    .Y(\i47/n387 ));
 AND2x4_ASAP7_75t_SL \i47/i440  (.A(\i47/n428 ),
    .B(\i47/n502 ),
    .Y(\i47/n433 ));
 AND2x4_ASAP7_75t_SL \i47/i441  (.A(\i47/n541 ),
    .B(\i47/n5 ),
    .Y(\i47/n434 ));
 OAI21xp33_ASAP7_75t_SL \i47/i442  (.A1(\i47/n43 ),
    .A2(\i47/n435 ),
    .B(\i47/n159 ),
    .Y(\i47/n436 ));
 NOR2xp33_ASAP7_75t_SL \i47/i443  (.A(\i47/n434 ),
    .B(\i47/n518 ),
    .Y(\i47/n435 ));
 OA21x2_ASAP7_75t_SL \i47/i444  (.A1(\i47/n40 ),
    .A2(\i47/n435 ),
    .B(\i47/n445 ),
    .Y(\i47/n437 ));
 INVx2_ASAP7_75t_SL \i47/i445  (.A(\i47/n449 ),
    .Y(\i47/n438 ));
 AOI221xp5_ASAP7_75t_SL \i47/i446  (.A1(\i47/n54 ),
    .A2(\i47/n38 ),
    .B1(\i47/n439 ),
    .B2(\i47/n55 ),
    .C(\i47/n170 ),
    .Y(\i47/n440 ));
 AND2x4_ASAP7_75t_SL \i47/i447  (.A(\i47/n5 ),
    .B(\i47/n438 ),
    .Y(\i47/n439 ));
 AND2x2_ASAP7_75t_SL \i47/i448  (.A(\i47/n7 ),
    .B(\i47/n439 ),
    .Y(\i47/n441 ));
 NAND2xp5_ASAP7_75t_SL \i47/i449  (.A(\i47/n41 ),
    .B(\i47/n439 ),
    .Y(\i47/n442 ));
 NOR2xp33_ASAP7_75t_SL \i47/i45  (.A(\i47/n332 ),
    .B(\i47/n356 ),
    .Y(\i47/n386 ));
 NAND2xp5_ASAP7_75t_SL \i47/i450  (.A(\i47/n70 ),
    .B(\i47/n439 ),
    .Y(\i47/n443 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i47/i451  (.A1(\i47/n434 ),
    .A2(\i47/n439 ),
    .B(\i47/n57 ),
    .C(\i47/n115 ),
    .Y(\i47/n444 ));
 NAND2xp5_ASAP7_75t_SL \i47/i452  (.A(\i47/n432 ),
    .B(\i47/n439 ),
    .Y(\i47/n445 ));
 OAI21xp5_ASAP7_75t_SL \i47/i453  (.A1(\i47/n61 ),
    .A2(\i47/n439 ),
    .B(\i47/n430 ),
    .Y(\i47/n446 ));
 AOI22xp33_ASAP7_75t_SL \i47/i454  (.A1(\i47/n70 ),
    .A2(\i47/n46 ),
    .B1(\i47/n532 ),
    .B2(\i47/n4 ),
    .Y(\i47/n447 ));
 NAND2x1_ASAP7_75t_SL \i47/i455  (.A(n27[3]),
    .B(\i47/n2 ),
    .Y(\i47/n448 ));
 OR2x2_ASAP7_75t_SL \i47/i456  (.A(n27[0]),
    .B(n27[1]),
    .Y(\i47/n449 ));
 OR2x4_ASAP7_75t_SL \i47/i457  (.A(\i47/n448 ),
    .B(\i47/n449 ),
    .Y(\i47/n450 ));
 INVx3_ASAP7_75t_SL \i47/i458  (.A(\i47/n450 ),
    .Y(\i47/n451 ));
 OAI221xp5_ASAP7_75t_SL \i47/i459  (.A1(\i47/n450 ),
    .A2(\i47/n67 ),
    .B1(\i47/n58 ),
    .B2(\i47/n470 ),
    .C(\i47/n91 ),
    .Y(\i47/n452 ));
 NAND3xp33_ASAP7_75t_SL \i47/i46  (.A(\i47/n322 ),
    .B(\i47/n330 ),
    .C(\i47/n299 ),
    .Y(\i47/n385 ));
 OAI221xp5_ASAP7_75t_SL \i47/i460  (.A1(\i47/n20 ),
    .A2(\i47/n450 ),
    .B1(\i47/n51 ),
    .B2(\i47/n481 ),
    .C(\i47/n139 ),
    .Y(\i47/n453 ));
 OAI22xp5_ASAP7_75t_SL \i47/i461  (.A1(\i47/n71 ),
    .A2(\i47/n450 ),
    .B1(\i47/n40 ),
    .B2(\i47/n10 ),
    .Y(\i47/n454 ));
 OAI22xp5_ASAP7_75t_SL \i47/i462  (.A1(\i47/n492 ),
    .A2(\i47/n450 ),
    .B1(\i47/n56 ),
    .B2(\i47/n68 ),
    .Y(\i47/n455 ));
 OAI22xp5_ASAP7_75t_SL \i47/i463  (.A1(\i47/n450 ),
    .A2(\i47/n43 ),
    .B1(\i47/n507 ),
    .B2(\i47/n15 ),
    .Y(\i47/n456 ));
 OAI22x1_ASAP7_75t_SL \i47/i464  (.A1(\i47/n16 ),
    .A2(\i47/n450 ),
    .B1(\i47/n507 ),
    .B2(\i47/n60 ),
    .Y(\i47/n457 ));
 NOR2xp67_ASAP7_75t_SL \i47/i465  (.A(\i47/n43 ),
    .B(\i47/n460 ),
    .Y(\i47/n461 ));
 OR2x6_ASAP7_75t_SL \i47/i466  (.A(\i47/n458 ),
    .B(\i47/n459 ),
    .Y(\i47/n460 ));
 INVx1_ASAP7_75t_SL \i47/i467  (.A(\i47/n32 ),
    .Y(\i47/n458 ));
 INVx2_ASAP7_75t_SL \i47/i468  (.A(\i47/n37 ),
    .Y(\i47/n459 ));
 OAI22xp5_ASAP7_75t_SL \i47/i469  (.A1(\i47/n69 ),
    .A2(\i47/n10 ),
    .B1(\i47/n470 ),
    .B2(\i47/n460 ),
    .Y(\i47/n462 ));
 NOR2x1_ASAP7_75t_SL \i47/i47  (.A(\i47/n285 ),
    .B(\i47/n341 ),
    .Y(\i47/n384 ));
 OAI221xp5_ASAP7_75t_SL \i47/i470  (.A1(\i47/n460 ),
    .A2(\i47/n65 ),
    .B1(\i47/n17 ),
    .B2(\i47/n16 ),
    .C(\i47/n203 ),
    .Y(\i47/n463 ));
 OAI222xp33_ASAP7_75t_SL \i47/i471  (.A1(\i47/n460 ),
    .A2(\i47/n40 ),
    .B1(\i47/n42 ),
    .B2(\i47/n16 ),
    .C1(\i47/n546 ),
    .C2(\i47/n56 ),
    .Y(\i47/n464 ));
 AOI21xp5_ASAP7_75t_L \i47/i472  (.A1(\i47/n52 ),
    .A2(\i47/n514 ),
    .B(\i47/n460 ),
    .Y(\i47/n465 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i47/i473  (.A1(\i47/n460 ),
    .A2(\i47/n42 ),
    .B(\i47/n481 ),
    .C(\i47/n517 ),
    .Y(\i47/n466 ));
 INVx3_ASAP7_75t_SL \i47/i474  (.A(\i47/n460 ),
    .Y(\i47/n467 ));
 NAND2xp5_ASAP7_75t_SL \i47/i475  (.A(\i47/n1 ),
    .B(n27[5]),
    .Y(\i47/n468 ));
 OAI221xp5_ASAP7_75t_SL \i47/i476  (.A1(\i47/n95 ),
    .A2(\i47/n69 ),
    .B1(\i47/n95 ),
    .B2(\i47/n470 ),
    .C(\i47/n539 ),
    .Y(\i47/n471 ));
 OR2x2_ASAP7_75t_SL \i47/i477  (.A(\i47/n469 ),
    .B(\i47/n468 ),
    .Y(\i47/n470 ));
 NAND2xp5_ASAP7_75t_SL \i47/i478  (.A(\i47/n0 ),
    .B(n27[6]),
    .Y(\i47/n469 ));
 NAND2xp5_ASAP7_75t_SL \i47/i479  (.A(\i47/n56 ),
    .B(\i47/n470 ),
    .Y(\i47/n472 ));
 NOR2xp33_ASAP7_75t_SL \i47/i48  (.A(\i47/n347 ),
    .B(\i47/n265 ),
    .Y(\i47/n383 ));
 OAI21xp5_ASAP7_75t_SL \i47/i480  (.A1(\i47/n470 ),
    .A2(\i47/n10 ),
    .B(\i47/n442 ),
    .Y(\i47/n473 ));
 AOI21xp5_ASAP7_75t_SL \i47/i481  (.A1(\i47/n476 ),
    .A2(\i47/n43 ),
    .B(\i47/n68 ),
    .Y(\i47/n474 ));
 OAI221xp5_ASAP7_75t_SL \i47/i482  (.A1(\i47/n48 ),
    .A2(\i47/n476 ),
    .B1(\i47/n43 ),
    .B2(\i47/n47 ),
    .C(\i47/n496 ),
    .Y(\i47/n475 ));
 OA21x2_ASAP7_75t_SL \i47/i483  (.A1(\i47/n476 ),
    .A2(\i47/n15 ),
    .B(\i47/n147 ),
    .Y(\i47/n477 ));
 AOI21xp33_ASAP7_75t_SL \i47/i484  (.A1(\i47/n56 ),
    .A2(\i47/n476 ),
    .B(\i47/n39 ),
    .Y(\i47/n478 ));
 NOR2xp67_ASAP7_75t_SL \i47/i485  (.A(\i47/n476 ),
    .B(\i47/n58 ),
    .Y(\i47/n479 ));
 NOR2xp33_ASAP7_75t_SL \i47/i486  (.A(\i47/n47 ),
    .B(\i47/n476 ),
    .Y(\i47/n480 ));
 INVx3_ASAP7_75t_SL \i47/i487  (.A(\i47/n57 ),
    .Y(\i47/n481 ));
 NAND2xp5_ASAP7_75t_SL \i47/i488  (.A(\i47/n433 ),
    .B(\i47/n66 ),
    .Y(\i47/n482 ));
 NAND2xp5_ASAP7_75t_SL \i47/i489  (.A(\i47/n72 ),
    .B(\i47/n4 ),
    .Y(\i47/n483 ));
 NAND2xp5_ASAP7_75t_SL \i47/i49  (.A(\i47/n354 ),
    .B(\i47/n349 ),
    .Y(\i47/n382 ));
 NOR2xp33_ASAP7_75t_SL \i47/i490  (.A(\i47/n418 ),
    .B(\i47/n485 ),
    .Y(\i47/n486 ));
 OAI211xp5_ASAP7_75t_SL \i47/i491  (.A1(\i47/n481 ),
    .A2(\i47/n484 ),
    .B(\i47/n482 ),
    .C(\i47/n483 ),
    .Y(\i47/n485 ));
 NOR2xp33_ASAP7_75t_SL \i47/i492  (.A(\i47/n434 ),
    .B(\i47/n4 ),
    .Y(\i47/n484 ));
 NOR5xp2_ASAP7_75t_SL \i47/i493  (.A(\i47/n485 ),
    .B(\i47/n475 ),
    .C(\i47/n452 ),
    .D(\i47/n24 ),
    .E(\i47/n427 ),
    .Y(\i47/n487 ));
 OR3x1_ASAP7_75t_SL \i47/i494  (.A(\i47/n488 ),
    .B(\i47/n452 ),
    .C(\i47/n24 ),
    .Y(\i47/n489 ));
 OAI211xp5_ASAP7_75t_SL \i47/i495  (.A1(\i47/n481 ),
    .A2(\i47/n484 ),
    .B(\i47/n482 ),
    .C(\i47/n483 ),
    .Y(\i47/n488 ));
 OAI21xp33_ASAP7_75t_SL \i47/i496  (.A1(\i47/n46 ),
    .A2(\i47/n439 ),
    .B(\i47/n490 ),
    .Y(\i47/n491 ));
 AND2x4_ASAP7_75t_SL \i47/i497  (.A(\i47/n502 ),
    .B(\i47/n531 ),
    .Y(\i47/n490 ));
 INVx4_ASAP7_75t_SL \i47/i498  (.A(\i47/n490 ),
    .Y(\i47/n492 ));
 OAI21xp5_ASAP7_75t_SL \i47/i499  (.A1(\i47/n490 ),
    .A2(\i47/n57 ),
    .B(\i47/n59 ),
    .Y(\i47/n493 ));
 INVx1_ASAP7_75t_SL \i47/i5  (.A(\i47/n29 ),
    .Y(\i47/n5 ));
 NOR2x1_ASAP7_75t_SL \i47/i50  (.A(\i47/n525 ),
    .B(\i47/n356 ),
    .Y(\i47/n381 ));
 OAI21xp5_ASAP7_75t_SL \i47/i500  (.A1(\i47/n432 ),
    .A2(\i47/n490 ),
    .B(\i47/n46 ),
    .Y(\i47/n494 ));
 AOI22xp5_ASAP7_75t_R \i47/i501  (.A1(\i47/n490 ),
    .A2(\i47/n66 ),
    .B1(\i47/n41 ),
    .B2(\i47/n50 ),
    .Y(\i47/n495 ));
 NAND2xp5_ASAP7_75t_SL \i47/i502  (.A(\i47/n490 ),
    .B(\i47/n61 ),
    .Y(\i47/n496 ));
 NAND2xp5_ASAP7_75t_SL \i47/i503  (.A(\i47/n490 ),
    .B(\i47/n63 ),
    .Y(\i47/n497 ));
 NAND2xp5_ASAP7_75t_SL \i47/i504  (.A(\i47/n4 ),
    .B(\i47/n490 ),
    .Y(\i47/n498 ));
 NAND2xp5_ASAP7_75t_SL \i47/i505  (.A(\i47/n490 ),
    .B(\i47/n45 ),
    .Y(\i47/n499 ));
 NAND2xp5_ASAP7_75t_SL \i47/i506  (.A(\i47/n490 ),
    .B(\i47/n518 ),
    .Y(\i47/n500 ));
 NAND2xp5_ASAP7_75t_SL \i47/i507  (.A(\i47/n490 ),
    .B(\i47/n467 ),
    .Y(\i47/n501 ));
 AND2x2_ASAP7_75t_SL \i47/i508  (.A(n27[4]),
    .B(\i47/n26 ),
    .Y(\i47/n502 ));
 AND2x2_ASAP7_75t_SL \i47/i509  (.A(n27[7]),
    .B(\i47/n13 ),
    .Y(\i47/n503 ));
 NOR2x1_ASAP7_75t_SL \i47/i51  (.A(\i47/n331 ),
    .B(\i47/n342 ),
    .Y(\i47/n380 ));
 AND2x4_ASAP7_75t_SL \i47/i510  (.A(\i47/n502 ),
    .B(\i47/n503 ),
    .Y(\i47/n504 ));
 OAI21xp5_ASAP7_75t_SL \i47/i511  (.A1(\i47/n38 ),
    .A2(\i47/n439 ),
    .B(\i47/n504 ),
    .Y(\i47/n505 ));
 AOI22xp5_ASAP7_75t_SL \i47/i512  (.A1(\i47/n504 ),
    .A2(\i47/n439 ),
    .B1(\i47/n50 ),
    .B2(\i47/n54 ),
    .Y(\i47/n506 ));
 INVx3_ASAP7_75t_SL \i47/i513  (.A(\i47/n504 ),
    .Y(\i47/n507 ));
 OAI31xp33_ASAP7_75t_SL \i47/i514  (.A1(\i47/n41 ),
    .A2(\i47/n504 ),
    .A3(\i47/n57 ),
    .B(\i47/n451 ),
    .Y(\i47/n508 ));
 OAI21xp5_ASAP7_75t_SL \i47/i515  (.A1(\i47/n59 ),
    .A2(\i47/n49 ),
    .B(\i47/n504 ),
    .Y(\i47/n509 ));
 OAI21xp5_ASAP7_75t_SL \i47/i516  (.A1(\i47/n434 ),
    .A2(\i47/n61 ),
    .B(\i47/n504 ),
    .Y(\i47/n510 ));
 AOI22xp5_ASAP7_75t_SL \i47/i517  (.A1(\i47/n432 ),
    .A2(\i47/n50 ),
    .B1(\i47/n504 ),
    .B2(\i47/n4 ),
    .Y(\i47/n511 ));
 AOI22xp5_ASAP7_75t_SL \i47/i518  (.A1(\i47/n504 ),
    .A2(\i47/n50 ),
    .B1(\i47/n41 ),
    .B2(\i47/n434 ),
    .Y(\i47/n512 ));
 AOI22xp5_ASAP7_75t_SL \i47/i519  (.A1(\i47/n38 ),
    .A2(\i47/n504 ),
    .B1(\i47/n57 ),
    .B2(\i47/n66 ),
    .Y(\i47/n513 ));
 NAND2xp5_ASAP7_75t_SL \i47/i52  (.A(\i47/n298 ),
    .B(\i47/n336 ),
    .Y(\i47/n379 ));
 NOR2xp33_ASAP7_75t_L \i47/i520  (.A(\i47/n70 ),
    .B(\i47/n504 ),
    .Y(\i47/n514 ));
 NAND2xp5_ASAP7_75t_SL \i47/i521  (.A(\i47/n504 ),
    .B(\i47/n63 ),
    .Y(\i47/n515 ));
 NAND2xp5_ASAP7_75t_SL \i47/i522  (.A(\i47/n504 ),
    .B(\i47/n518 ),
    .Y(\i47/n516 ));
 NAND2xp5_ASAP7_75t_SL \i47/i523  (.A(\i47/n504 ),
    .B(\i47/n66 ),
    .Y(\i47/n517 ));
 AND2x4_ASAP7_75t_SL \i47/i524  (.A(\i47/n37 ),
    .B(\i47/n31 ),
    .Y(\i47/n518 ));
 OAI22xp5_ASAP7_75t_SL \i47/i525  (.A1(\i47/n476 ),
    .A2(\i47/n519 ),
    .B1(\i47/n481 ),
    .B2(\i47/n460 ),
    .Y(\i47/n520 ));
 INVx4_ASAP7_75t_SL \i47/i526  (.A(\i47/n518 ),
    .Y(\i47/n519 ));
 OAI222xp33_ASAP7_75t_SL \i47/i527  (.A1(\i47/n519 ),
    .A2(\i47/n65 ),
    .B1(\i47/n450 ),
    .B2(\i47/n64 ),
    .C1(\i47/n17 ),
    .C2(\i47/n52 ),
    .Y(\i47/n521 ));
 OAI22xp5_ASAP7_75t_SL \i47/i528  (.A1(\i47/n69 ),
    .A2(\i47/n48 ),
    .B1(\i47/n519 ),
    .B2(\i47/n492 ),
    .Y(\i47/n522 ));
 OAI22xp5_ASAP7_75t_L \i47/i529  (.A1(\i47/n65 ),
    .A2(\i47/n39 ),
    .B1(\i47/n40 ),
    .B2(\i47/n519 ),
    .Y(\i47/n523 ));
 NOR2x1_ASAP7_75t_SL \i47/i53  (.A(\i47/n343 ),
    .B(\i47/n9 ),
    .Y(\i47/n378 ));
 OAI22xp5_ASAP7_75t_SL \i47/i530  (.A1(\i47/n519 ),
    .A2(\i47/n137 ),
    .B1(\i47/n56 ),
    .B2(\i47/n80 ),
    .Y(\i47/n524 ));
 OAI211xp5_ASAP7_75t_SL \i47/i531  (.A1(\i47/n69 ),
    .A2(\i47/n519 ),
    .B(\i47/n155 ),
    .C(\i47/n109 ),
    .Y(\i47/n525 ));
 OAI22xp5_ASAP7_75t_SL \i47/i532  (.A1(\i47/n481 ),
    .A2(\i47/n519 ),
    .B1(\i47/n58 ),
    .B2(\i47/n507 ),
    .Y(\i47/n526 ));
 AOI21xp33_ASAP7_75t_SL \i47/i533  (.A1(\i47/n58 ),
    .A2(\i47/n519 ),
    .B(\i47/n65 ),
    .Y(\i47/n527 ));
 OAI22xp5_ASAP7_75t_SL \i47/i534  (.A1(\i47/n43 ),
    .A2(\i47/n519 ),
    .B1(\i47/n56 ),
    .B2(\i47/n47 ),
    .Y(\i47/n528 ));
 OAI22xp5_ASAP7_75t_SL \i47/i535  (.A1(\i47/n52 ),
    .A2(\i47/n42 ),
    .B1(\i47/n56 ),
    .B2(\i47/n519 ),
    .Y(\i47/n529 ));
 AND2x4_ASAP7_75t_SL \i47/i536  (.A(\i47/n26 ),
    .B(\i47/n1 ),
    .Y(\i47/n530 ));
 AND2x2_ASAP7_75t_L \i47/i537  (.A(\i47/n0 ),
    .B(n27[6]),
    .Y(\i47/n531 ));
 OR2x2_ASAP7_75t_SL \i47/i538  (.A(\i47/n504 ),
    .B(\i47/n532 ),
    .Y(\i47/n533 ));
 AND2x4_ASAP7_75t_SL \i47/i539  (.A(\i47/n530 ),
    .B(\i47/n531 ),
    .Y(\i47/n532 ));
 NAND2xp5_ASAP7_75t_SL \i47/i54  (.A(\i47/n340 ),
    .B(\i47/n320 ),
    .Y(\i47/n390 ));
 INVx3_ASAP7_75t_SL \i47/i540  (.A(\i47/n532 ),
    .Y(\i47/n476 ));
 NAND2xp5_ASAP7_75t_SL \i47/i541  (.A(\i47/n63 ),
    .B(\i47/n532 ),
    .Y(\i47/n534 ));
 NAND2xp5_ASAP7_75t_SL \i47/i542  (.A(\i47/n532 ),
    .B(\i47/n4 ),
    .Y(\i47/n535 ));
 AOI22xp33_ASAP7_75t_SL \i47/i543  (.A1(\i47/n532 ),
    .A2(\i47/n61 ),
    .B1(\i47/n7 ),
    .B2(\i47/n46 ),
    .Y(\i47/n536 ));
 AOI22xp5_ASAP7_75t_SL \i47/i544  (.A1(\i47/n532 ),
    .A2(\i47/n50 ),
    .B1(\i47/n72 ),
    .B2(\i47/n49 ),
    .Y(\i47/n537 ));
 AOI22xp5_ASAP7_75t_SL \i47/i545  (.A1(\i47/n532 ),
    .A2(\i47/n451 ),
    .B1(\i47/n7 ),
    .B2(\i47/n66 ),
    .Y(\i47/n538 ));
 AOI211x1_ASAP7_75t_SL \i47/i546  (.A1(\i47/n85 ),
    .A2(\i47/n532 ),
    .B(\i47/n156 ),
    .C(\i47/n158 ),
    .Y(\i47/n539 ));
 NAND2xp5_ASAP7_75t_SL \i47/i547  (.A(\i47/n532 ),
    .B(\i47/n439 ),
    .Y(\i47/n540 ));
 AND2x2_ASAP7_75t_SL \i47/i548  (.A(n27[0]),
    .B(n27[1]),
    .Y(\i47/n541 ));
 AND2x4_ASAP7_75t_SL \i47/i549  (.A(n27[2]),
    .B(n27[3]),
    .Y(\i47/n542 ));
 NOR2x1_ASAP7_75t_SL \i47/i55  (.A(\i47/n357 ),
    .B(\i47/n342 ),
    .Y(\i47/n377 ));
 OAI31xp33_ASAP7_75t_SL \i47/i550  (.A1(\i47/n543 ),
    .A2(\i47/n4 ),
    .A3(\i47/n45 ),
    .B(\i47/n504 ),
    .Y(\i47/n544 ));
 AND2x4_ASAP7_75t_SL \i47/i551  (.A(\i47/n541 ),
    .B(\i47/n542 ),
    .Y(\i47/n543 ));
 AOI22xp5_ASAP7_75t_SL \i47/i552  (.A1(\i47/n72 ),
    .A2(\i47/n439 ),
    .B1(\i47/n53 ),
    .B2(\i47/n543 ),
    .Y(\i47/n545 ));
 INVx2_ASAP7_75t_SL \i47/i553  (.A(\i47/n543 ),
    .Y(\i47/n546 ));
 AOI211xp5_ASAP7_75t_SL \i47/i554  (.A1(\i47/n138 ),
    .A2(\i47/n543 ),
    .B(\i47/n564 ),
    .C(\i47/n154 ),
    .Y(\i47/n547 ));
 OAI31xp33_ASAP7_75t_R \i47/i555  (.A1(\i47/n543 ),
    .A2(\i47/n61 ),
    .A3(\i47/n63 ),
    .B(\i47/n57 ),
    .Y(\i47/n548 ));
 OAI21xp5_ASAP7_75t_SL \i47/i556  (.A1(\i47/n559 ),
    .A2(\i47/n136 ),
    .B(\i47/n543 ),
    .Y(\i47/n549 ));
 AOI22xp5_ASAP7_75t_SL \i47/i557  (.A1(\i47/n70 ),
    .A2(\i47/n84 ),
    .B1(\i47/n41 ),
    .B2(\i47/n543 ),
    .Y(\i47/n550 ));
 AOI222xp33_ASAP7_75t_SL \i47/i558  (.A1(\i47/n63 ),
    .A2(\i47/n54 ),
    .B1(\i47/n7 ),
    .B2(\i47/n38 ),
    .C1(\i47/n543 ),
    .C2(\i47/n559 ),
    .Y(\i47/n551 ));
 AOI22xp5_ASAP7_75t_SL \i47/i559  (.A1(\i47/n430 ),
    .A2(\i47/n49 ),
    .B1(\i47/n433 ),
    .B2(\i47/n543 ),
    .Y(\i47/n552 ));
 NOR2x1_ASAP7_75t_SL \i47/i56  (.A(\i47/n284 ),
    .B(\i47/n341 ),
    .Y(\i47/n389 ));
 AOI22xp5_ASAP7_75t_SL \i47/i560  (.A1(\i47/n434 ),
    .A2(\i47/n72 ),
    .B1(\i47/n432 ),
    .B2(\i47/n543 ),
    .Y(\i47/n553 ));
 NAND2xp5_ASAP7_75t_SL \i47/i561  (.A(\i47/n543 ),
    .B(\i47/n57 ),
    .Y(\i47/n554 ));
 NAND2xp5_ASAP7_75t_SL \i47/i562  (.A(\i47/n54 ),
    .B(\i47/n543 ),
    .Y(\i47/n555 ));
 AND2x2_ASAP7_75t_SL \i47/i563  (.A(\i47/n72 ),
    .B(\i47/n543 ),
    .Y(\i47/n556 ));
 NAND2xp5_ASAP7_75t_SL \i47/i564  (.A(\i47/n543 ),
    .B(\i47/n7 ),
    .Y(\i47/n557 ));
 NAND2xp5_ASAP7_75t_SL \i47/i565  (.A(\i47/n70 ),
    .B(\i47/n543 ),
    .Y(\i47/n558 ));
 AND2x4_ASAP7_75t_SL \i47/i566  (.A(\i47/n502 ),
    .B(\i47/n34 ),
    .Y(\i47/n559 ));
 NOR2xp33_ASAP7_75t_SL \i47/i567  (.A(\i47/n560 ),
    .B(\i47/n519 ),
    .Y(\i47/n424 ));
 INVx3_ASAP7_75t_SL \i47/i568  (.A(\i47/n559 ),
    .Y(\i47/n560 ));
 OAI22xp5_ASAP7_75t_SL \i47/i569  (.A1(\i47/n17 ),
    .A2(\i47/n560 ),
    .B1(\i47/n519 ),
    .B2(\i47/n67 ),
    .Y(\i47/n561 ));
 INVxp67_ASAP7_75t_SL \i47/i57  (.A(\i47/n375 ),
    .Y(\i47/n376 ));
 OAI22x1_ASAP7_75t_SL \i47/i570  (.A1(\i47/n62 ),
    .A2(\i47/n560 ),
    .B1(\i47/n546 ),
    .B2(\i47/n476 ),
    .Y(\i47/n562 ));
 OAI22xp33_ASAP7_75t_SL \i47/i571  (.A1(\i47/n560 ),
    .A2(\i47/n39 ),
    .B1(\i47/n460 ),
    .B2(\i47/n52 ),
    .Y(\i47/n563 ));
 OAI22xp5_ASAP7_75t_SL \i47/i572  (.A1(\i47/n560 ),
    .A2(\i47/n460 ),
    .B1(\i47/n71 ),
    .B2(\i47/n15 ),
    .Y(\i47/n564 ));
 OAI22xp33_ASAP7_75t_SL \i47/i573  (.A1(\i47/n507 ),
    .A2(\i47/n450 ),
    .B1(\i47/n47 ),
    .B2(\i47/n560 ),
    .Y(\i47/n565 ));
 OAI22xp5_ASAP7_75t_SL \i47/i574  (.A1(\i47/n560 ),
    .A2(\i47/n450 ),
    .B1(\i47/n56 ),
    .B2(\i47/n15 ),
    .Y(\i47/n566 ));
 NOR2xp33_ASAP7_75t_SL \i47/i575  (.A(\i47/n560 ),
    .B(\i47/n68 ),
    .Y(\i47/n567 ));
 OAI22xp33_ASAP7_75t_SL \i47/i576  (.A1(\i47/n42 ),
    .A2(\i47/n560 ),
    .B1(\i47/n15 ),
    .B2(\i47/n43 ),
    .Y(\i47/n568 ));
 OAI21xp33_ASAP7_75t_SL \i47/i577  (.A1(\i47/n60 ),
    .A2(\i47/n560 ),
    .B(\i47/n150 ),
    .Y(\i47/n569 ));
 AND4x1_ASAP7_75t_SL \i47/i578  (.A(\i47/n551 ),
    .B(\i47/n267 ),
    .C(\i47/n575 ),
    .D(\i47/n477 ),
    .Y(\i47/n570 ));
 AND4x1_ASAP7_75t_SL \i47/i579  (.A(\i47/n229 ),
    .B(\i47/n269 ),
    .C(\i47/n245 ),
    .D(\i47/n551 ),
    .Y(\i47/n571 ));
 INVxp67_ASAP7_75t_SL \i47/i58  (.A(\i47/n371 ),
    .Y(\i47/n372 ));
 OR4x1_ASAP7_75t_SL \i47/i580  (.A(\i47/n474 ),
    .B(\i47/n211 ),
    .C(\i47/n210 ),
    .D(\i47/n206 ),
    .Y(\i47/n572 ));
 OAI21xp5_ASAP7_75t_SL \i47/i581  (.A1(\i47/n4 ),
    .A2(\i47/n61 ),
    .B(\i47/n41 ),
    .Y(\i47/n573 ));
 AND3x1_ASAP7_75t_SL \i47/i582  (.A(\i47/n573 ),
    .B(\i47/n237 ),
    .C(\i47/n302 ),
    .Y(\i47/n574 ));
 AOI21xp5_ASAP7_75t_SL \i47/i583  (.A1(\i47/n44 ),
    .A2(\i47/n543 ),
    .B(\i47/n170 ),
    .Y(\i47/n575 ));
 NOR3xp33_ASAP7_75t_SL \i47/i584  (.A(\i47/n576 ),
    .B(\i47/n257 ),
    .C(\i47/n121 ),
    .Y(\i47/n577 ));
 OAI21xp5_ASAP7_75t_SL \i47/i585  (.A1(\i47/n481 ),
    .A2(\i47/n519 ),
    .B(\i47/n558 ),
    .Y(\i47/n576 ));
 NOR3xp33_ASAP7_75t_SL \i47/i586  (.A(\i47/n578 ),
    .B(\i47/n436 ),
    .C(\i47/n562 ),
    .Y(\i47/n579 ));
 OAI21xp5_ASAP7_75t_SL \i47/i587  (.A1(\i47/n56 ),
    .A2(\i47/n17 ),
    .B(\i47/n498 ),
    .Y(\i47/n578 ));
 AND5x1_ASAP7_75t_SL \i47/i59  (.A(\i47/n295 ),
    .B(\i47/n575 ),
    .C(\i47/n289 ),
    .D(\i47/n228 ),
    .E(\i47/n446 ),
    .Y(\i47/n370 ));
 INVx2_ASAP7_75t_SL \i47/i6  (.A(\i47/n35 ),
    .Y(\i47/n6 ));
 NOR3xp33_ASAP7_75t_SL \i47/i60  (.A(\i47/n304 ),
    .B(\i47/n288 ),
    .C(\i47/n270 ),
    .Y(\i47/n369 ));
 NOR3xp33_ASAP7_75t_SL \i47/i61  (.A(\i47/n328 ),
    .B(\i47/n271 ),
    .C(\i47/n236 ),
    .Y(\i47/n368 ));
 AND5x1_ASAP7_75t_SL \i47/i62  (.A(\i47/n261 ),
    .B(\i47/n274 ),
    .C(\i47/n431 ),
    .D(\i47/n264 ),
    .E(\i47/n212 ),
    .Y(\i47/n367 ));
 NOR2xp33_ASAP7_75t_SL \i47/i63  (.A(\i47/n329 ),
    .B(\i47/n334 ),
    .Y(\i47/n366 ));
 NAND5xp2_ASAP7_75t_SL \i47/i64  (.A(\i47/n547 ),
    .B(\i47/n182 ),
    .C(\i47/n256 ),
    .D(\i47/n172 ),
    .E(\i47/n12 ),
    .Y(\i47/n365 ));
 NOR4xp25_ASAP7_75t_SL \i47/i65  (.A(\i47/n286 ),
    .B(\i47/n475 ),
    .C(\i47/n246 ),
    .D(\i47/n230 ),
    .Y(\i47/n364 ));
 NAND4xp25_ASAP7_75t_SL \i47/i66  (.A(\i47/n302 ),
    .B(\i47/n314 ),
    .C(\i47/n317 ),
    .D(\i47/n319 ),
    .Y(\i47/n363 ));
 NAND4xp25_ASAP7_75t_SL \i47/i67  (.A(\i47/n326 ),
    .B(\i47/n324 ),
    .C(\i47/n164 ),
    .D(\i47/n208 ),
    .Y(\i47/n362 ));
 NOR2x1_ASAP7_75t_SL \i47/i68  (.A(\i47/n168 ),
    .B(\i47/n353 ),
    .Y(\i47/n361 ));
 NAND3xp33_ASAP7_75t_SL \i47/i69  (.A(\i47/n319 ),
    .B(\i47/n294 ),
    .C(\i47/n516 ),
    .Y(\i47/n375 ));
 INVx2_ASAP7_75t_SL \i47/i7  (.A(\i47/n470 ),
    .Y(\i47/n7 ));
 NAND4xp75_ASAP7_75t_SL \i47/i70  (.A(\i47/n539 ),
    .B(\i47/n220 ),
    .C(\i47/n283 ),
    .D(\i47/n557 ),
    .Y(\i47/n374 ));
 NAND2xp33_ASAP7_75t_L \i47/i71  (.A(\i47/n301 ),
    .B(\i47/n358 ),
    .Y(\i47/n360 ));
 AND2x2_ASAP7_75t_SL \i47/i72  (.A(\i47/n303 ),
    .B(\i47/n348 ),
    .Y(\i47/n373 ));
 NAND2x1p5_ASAP7_75t_SL \i47/i73  (.A(\i47/n355 ),
    .B(\i47/n313 ),
    .Y(\i47/n371 ));
 INVx1_ASAP7_75t_L \i47/i74  (.A(\i47/n358 ),
    .Y(\i47/n359 ));
 INVxp67_ASAP7_75t_SL \i47/i75  (.A(\i47/n352 ),
    .Y(\i47/n353 ));
 NOR5xp2_ASAP7_75t_SL \i47/i76  (.A(\i47/n465 ),
    .B(\i47/n235 ),
    .C(\i47/n457 ),
    .D(\i47/n556 ),
    .E(\i47/n76 ),
    .Y(\i47/n350 ));
 NOR3xp33_ASAP7_75t_SL \i47/i77  (.A(\i47/n323 ),
    .B(\i47/n249 ),
    .C(\i47/n521 ),
    .Y(\i47/n349 ));
 NOR2xp33_ASAP7_75t_SL \i47/i78  (.A(\i47/n321 ),
    .B(\i47/n276 ),
    .Y(\i47/n348 ));
 NOR2x1_ASAP7_75t_SL \i47/i79  (.A(\i47/n290 ),
    .B(\i47/n262 ),
    .Y(\i47/n358 ));
 NOR2x2_ASAP7_75t_SL \i47/i8  (.A(\i47/n413 ),
    .B(\i47/n412 ),
    .Y(n26[4]));
 NAND3xp33_ASAP7_75t_SL \i47/i80  (.A(\i47/n550 ),
    .B(\i47/n544 ),
    .C(\i47/n553 ),
    .Y(\i47/n347 ));
 NAND2xp5_ASAP7_75t_L \i47/i81  (.A(\i47/n320 ),
    .B(\i47/n293 ),
    .Y(\i47/n346 ));
 NAND2xp5_ASAP7_75t_SL \i47/i82  (.A(\i47/n311 ),
    .B(\i47/n275 ),
    .Y(\i47/n345 ));
 NAND3xp33_ASAP7_75t_SL \i47/i83  (.A(\i47/n575 ),
    .B(\i47/n232 ),
    .C(\i47/n477 ),
    .Y(\i47/n357 ));
 NOR3xp33_ASAP7_75t_SL \i47/i84  (.A(\i47/n471 ),
    .B(\i47/n8 ),
    .C(\i47/n463 ),
    .Y(\i47/n344 ));
 NAND2xp5_ASAP7_75t_SL \i47/i85  (.A(\i47/n21 ),
    .B(\i47/n302 ),
    .Y(\i47/n356 ));
 NOR2x1_ASAP7_75t_SL \i47/i86  (.A(\i47/n521 ),
    .B(\i47/n323 ),
    .Y(\i47/n355 ));
 NOR2xp33_ASAP7_75t_SL \i47/i87  (.A(\i47/n287 ),
    .B(\i47/n273 ),
    .Y(\i47/n354 ));
 NOR2xp33_ASAP7_75t_SL \i47/i88  (.A(\i47/n453 ),
    .B(\i47/n310 ),
    .Y(\i47/n352 ));
 NOR3x1_ASAP7_75t_SL \i47/i89  (.A(\i47/n242 ),
    .B(\i47/n167 ),
    .C(\i47/n280 ),
    .Y(\i47/n351 ));
 NOR2x2_ASAP7_75t_SL \i47/i9  (.A(\i47/n408 ),
    .B(\i47/n414 ),
    .Y(n26[3]));
 NOR3xp33_ASAP7_75t_SL \i47/i90  (.A(\i47/n247 ),
    .B(\i47/n181 ),
    .C(\i47/n239 ),
    .Y(\i47/n340 ));
 NOR2xp33_ASAP7_75t_SL \i47/i91  (.A(\i47/n297 ),
    .B(\i47/n572 ),
    .Y(\i47/n339 ));
 NAND3xp33_ASAP7_75t_SL \i47/i92  (.A(\i47/n551 ),
    .B(\i47/n425 ),
    .C(\i47/n245 ),
    .Y(\i47/n338 ));
 NAND4xp25_ASAP7_75t_SL \i47/i93  (.A(\i47/n437 ),
    .B(\i47/n444 ),
    .C(\i47/n548 ),
    .D(\i47/n231 ),
    .Y(\i47/n337 ));
 NAND2xp5_ASAP7_75t_SL \i47/i94  (.A(\i47/n309 ),
    .B(\i47/n322 ),
    .Y(\i47/n343 ));
 NOR5xp2_ASAP7_75t_SL \i47/i95  (.A(\i47/n318 ),
    .B(\i47/n466 ),
    .C(\i47/n107 ),
    .D(\i47/n478 ),
    .E(\i47/n140 ),
    .Y(\i47/n336 ));
 NAND3xp33_ASAP7_75t_SL \i47/i96  (.A(\i47/n279 ),
    .B(\i47/n577 ),
    .C(\i47/n184 ),
    .Y(\i47/n335 ));
 NAND2xp33_ASAP7_75t_SL \i47/i97  (.A(\i47/n233 ),
    .B(\i47/n315 ),
    .Y(\i47/n334 ));
 NOR5xp2_ASAP7_75t_SL \i47/i98  (.A(\i47/n263 ),
    .B(\i47/n453 ),
    .C(\i47/n253 ),
    .D(\i47/n213 ),
    .E(\i47/n175 ),
    .Y(\i47/n333 ));
 NAND5xp2_ASAP7_75t_SL \i47/i99  (.A(\i47/n440 ),
    .B(\i47/n277 ),
    .C(\i47/n545 ),
    .D(\i47/n251 ),
    .E(\i47/n537 ),
    .Y(\i47/n332 ));
 XOR2xp5_ASAP7_75t_SL i470 (.A(n812),
    .B(n587),
    .Y(n1002));
 OAI22xp5_ASAP7_75t_SL i471 (.A1(n825),
    .A2(n1167),
    .B1(n795),
    .B2(n824),
    .Y(n1001));
 XNOR2xp5_ASAP7_75t_SL i472 (.A(n586),
    .B(n804),
    .Y(n1000));
 XOR2xp5_ASAP7_75t_SL i473 (.A(n585),
    .B(n584),
    .Y(n999));
 AOI22xp5_ASAP7_75t_SL i474 (.A1(n1175),
    .A2(n820),
    .B1(n792),
    .B2(n821),
    .Y(n998));
 OAI22xp5_ASAP7_75t_SL i475 (.A1(n1174),
    .A2(n809),
    .B1(n810),
    .B2(n822),
    .Y(n997));
 XNOR2xp5_ASAP7_75t_SL i476 (.A(n605),
    .B(n811),
    .Y(n996));
 OAI22xp5_ASAP7_75t_SL i477 (.A1(n832),
    .A2(n810),
    .B1(n833),
    .B2(n809),
    .Y(n995));
 AOI22xp5_ASAP7_75t_SL i478 (.A1(n836),
    .A2(n1155),
    .B1(n224),
    .B2(n226),
    .Y(n994));
 XNOR2xp5_ASAP7_75t_SL i479 (.A(n330),
    .B(n595),
    .Y(n993));
 INVx2_ASAP7_75t_SL \i48/i0  (.A(n25[5]),
    .Y(\i48/n0 ));
 INVxp67_ASAP7_75t_SL \i48/i1  (.A(n25[4]),
    .Y(\i48/n1 ));
 NOR2x1p5_ASAP7_75t_SL \i48/i10  (.A(\i48/n447 ),
    .B(\i48/n438 ),
    .Y(n24[5]));
 NAND5xp2_ASAP7_75t_SL \i48/i100  (.A(\i48/n236 ),
    .B(\i48/n474 ),
    .C(\i48/n495 ),
    .D(\i48/n272 ),
    .E(\i48/n523 ),
    .Y(\i48/n360 ));
 NAND3xp33_ASAP7_75t_SL \i48/i101  (.A(\i48/n232 ),
    .B(\i48/n258 ),
    .C(\i48/n327 ),
    .Y(\i48/n359 ));
 NOR5xp2_ASAP7_75t_SL \i48/i102  (.A(\i48/n230 ),
    .B(\i48/n240 ),
    .C(\i48/n225 ),
    .D(\i48/n91 ),
    .E(\i48/n460 ),
    .Y(\i48/n358 ));
 NAND5xp2_ASAP7_75t_SL \i48/i103  (.A(\i48/n21 ),
    .B(\i48/n513 ),
    .C(\i48/n495 ),
    .D(\i48/n542 ),
    .E(\i48/n159 ),
    .Y(\i48/n357 ));
 NOR5xp2_ASAP7_75t_SL \i48/i104  (.A(\i48/n195 ),
    .B(\i48/n514 ),
    .C(\i48/n183 ),
    .D(\i48/n154 ),
    .E(\i48/n152 ),
    .Y(\i48/n356 ));
 NOR2xp33_ASAP7_75t_SL \i48/i105  (.A(\i48/n317 ),
    .B(\i48/n350 ),
    .Y(\i48/n355 ));
 NOR2xp33_ASAP7_75t_SL \i48/i106  (.A(\i48/n305 ),
    .B(\i48/n336 ),
    .Y(\i48/n354 ));
 NAND3x1_ASAP7_75t_SL \i48/i107  (.A(\i48/n499 ),
    .B(\i48/n334 ),
    .C(\i48/n474 ),
    .Y(\i48/n370 ));
 NAND3x1_ASAP7_75t_SL \i48/i108  (.A(\i48/n296 ),
    .B(\i48/n278 ),
    .C(\i48/n248 ),
    .Y(\i48/n369 ));
 AOI21xp5_ASAP7_75t_L \i48/i109  (.A1(\i48/n56 ),
    .A2(\i48/n198 ),
    .B(\i48/n136 ),
    .Y(\i48/n347 ));
 AND2x4_ASAP7_75t_SL \i48/i11  (.A(\i48/n448 ),
    .B(\i48/n431 ),
    .Y(n24[0]));
 NOR2xp33_ASAP7_75t_SL \i48/i110  (.A(\i48/n509 ),
    .B(\i48/n287 ),
    .Y(\i48/n346 ));
 NAND2xp5_ASAP7_75t_SL \i48/i111  (.A(\i48/n276 ),
    .B(\i48/n304 ),
    .Y(\i48/n345 ));
 NOR2xp33_ASAP7_75t_SL \i48/i112  (.A(\i48/n303 ),
    .B(\i48/n22 ),
    .Y(\i48/n344 ));
 NOR2xp33_ASAP7_75t_SL \i48/i113  (.A(\i48/n282 ),
    .B(\i48/n292 ),
    .Y(\i48/n343 ));
 NOR2xp67_ASAP7_75t_SL \i48/i114  (.A(\i48/n144 ),
    .B(\i48/n289 ),
    .Y(\i48/n342 ));
 NOR2xp33_ASAP7_75t_SL \i48/i115  (.A(\i48/n18 ),
    .B(\i48/n287 ),
    .Y(\i48/n341 ));
 NOR4xp25_ASAP7_75t_SL \i48/i116  (.A(\i48/n261 ),
    .B(\i48/n18 ),
    .C(\i48/n477 ),
    .D(\i48/n519 ),
    .Y(\i48/n340 ));
 NAND2xp5_ASAP7_75t_SL \i48/i117  (.A(\i48/n222 ),
    .B(\i48/n269 ),
    .Y(\i48/n339 ));
 NOR4xp25_ASAP7_75t_SL \i48/i118  (.A(\i48/n89 ),
    .B(\i48/n215 ),
    .C(\i48/n186 ),
    .D(\i48/n199 ),
    .Y(\i48/n338 ));
 NOR3xp33_ASAP7_75t_SL \i48/i119  (.A(\i48/n219 ),
    .B(\i48/n458 ),
    .C(\i48/n218 ),
    .Y(\i48/n337 ));
 NOR3xp33_ASAP7_75t_SL \i48/i12  (.A(\i48/n422 ),
    .B(\i48/n418 ),
    .C(\i48/n451 ),
    .Y(\i48/n448 ));
 NAND2xp33_ASAP7_75t_SL \i48/i120  (.A(\i48/n525 ),
    .B(\i48/n19 ),
    .Y(\i48/n336 ));
 NOR2xp33_ASAP7_75t_SL \i48/i121  (.A(\i48/n509 ),
    .B(\i48/n254 ),
    .Y(\i48/n335 ));
 NOR2x1p5_ASAP7_75t_SL \i48/i122  (.A(\i48/n237 ),
    .B(\i48/n570 ),
    .Y(\i48/n334 ));
 NAND2xp33_ASAP7_75t_SL \i48/i123  (.A(\i48/n301 ),
    .B(\i48/n285 ),
    .Y(\i48/n333 ));
 NAND3xp33_ASAP7_75t_SL \i48/i124  (.A(\i48/n20 ),
    .B(\i48/n539 ),
    .C(\i48/n566 ),
    .Y(\i48/n332 ));
 NOR3xp33_ASAP7_75t_SL \i48/i125  (.A(\i48/n179 ),
    .B(\i48/n192 ),
    .C(\i48/n167 ),
    .Y(\i48/n353 ));
 NAND2xp5_ASAP7_75t_SL \i48/i126  (.A(\i48/n12 ),
    .B(\i48/n178 ),
    .Y(\i48/n352 ));
 NOR2x1_ASAP7_75t_SL \i48/i127  (.A(\i48/n235 ),
    .B(\i48/n256 ),
    .Y(\i48/n351 ));
 NAND2xp5_ASAP7_75t_SL \i48/i128  (.A(\i48/n495 ),
    .B(\i48/n262 ),
    .Y(\i48/n350 ));
 NOR2x1_ASAP7_75t_SL \i48/i129  (.A(\i48/n577 ),
    .B(\i48/n290 ),
    .Y(\i48/n349 ));
 NOR2x2_ASAP7_75t_SL \i48/i13  (.A(\i48/n440 ),
    .B(\i48/n441 ),
    .Y(n24[2]));
 NOR3x1_ASAP7_75t_SL \i48/i130  (.A(\i48/n183 ),
    .B(\i48/n554 ),
    .C(\i48/n151 ),
    .Y(\i48/n348 ));
 INVx1_ASAP7_75t_SL \i48/i131  (.A(\i48/n329 ),
    .Y(\i48/n330 ));
 INVx1_ASAP7_75t_SL \i48/i132  (.A(\i48/n23 ),
    .Y(\i48/n328 ));
 NOR4xp25_ASAP7_75t_SL \i48/i133  (.A(\i48/n463 ),
    .B(\i48/n202 ),
    .C(\i48/n190 ),
    .D(\i48/n165 ),
    .Y(\i48/n327 ));
 AOI211xp5_ASAP7_75t_SL \i48/i134  (.A1(\i48/n55 ),
    .A2(\i48/n50 ),
    .B(\i48/n570 ),
    .C(\i48/n148 ),
    .Y(\i48/n326 ));
 AOI211xp5_ASAP7_75t_SL \i48/i135  (.A1(\i48/n93 ),
    .A2(\i48/n43 ),
    .B(\i48/n273 ),
    .C(\i48/n217 ),
    .Y(\i48/n325 ));
 NAND2xp33_ASAP7_75t_SL \i48/i136  (.A(\i48/n249 ),
    .B(\i48/n271 ),
    .Y(\i48/n324 ));
 NAND5xp2_ASAP7_75t_SL \i48/i137  (.A(\i48/n200 ),
    .B(\i48/n213 ),
    .C(\i48/n224 ),
    .D(\i48/n488 ),
    .E(\i48/n505 ),
    .Y(\i48/n323 ));
 NOR4xp25_ASAP7_75t_SL \i48/i138  (.A(\i48/n280 ),
    .B(\i48/n118 ),
    .C(\i48/n120 ),
    .D(\i48/n141 ),
    .Y(\i48/n322 ));
 NOR2xp33_ASAP7_75t_SL \i48/i139  (.A(\i48/n241 ),
    .B(\i48/n244 ),
    .Y(\i48/n321 ));
 NAND4xp75_ASAP7_75t_SL \i48/i14  (.A(\i48/n408 ),
    .B(\i48/n426 ),
    .C(\i48/n406 ),
    .D(\i48/n575 ),
    .Y(\i48/n447 ));
 AOI211xp5_ASAP7_75t_SL \i48/i140  (.A1(\i48/n139 ),
    .A2(\i48/n57 ),
    .B(\i48/n465 ),
    .C(\i48/n156 ),
    .Y(\i48/n320 ));
 OA21x2_ASAP7_75t_SL \i48/i141  (.A1(\i48/n535 ),
    .A2(\i48/n56 ),
    .B(\i48/n513 ),
    .Y(\i48/n319 ));
 NOR4xp25_ASAP7_75t_SL \i48/i142  (.A(\i48/n226 ),
    .B(\i48/n147 ),
    .C(\i48/n174 ),
    .D(\i48/n151 ),
    .Y(\i48/n318 ));
 NAND5xp2_ASAP7_75t_SL \i48/i143  (.A(\i48/n119 ),
    .B(\i48/n80 ),
    .C(\i48/n129 ),
    .D(\i48/n121 ),
    .E(\i48/n74 ),
    .Y(\i48/n317 ));
 NOR3xp33_ASAP7_75t_SL \i48/i144  (.A(\i48/n257 ),
    .B(\i48/n149 ),
    .C(\i48/n73 ),
    .Y(\i48/n316 ));
 NAND2xp5_ASAP7_75t_SL \i48/i145  (.A(\i48/n239 ),
    .B(\i48/n21 ),
    .Y(\i48/n315 ));
 NAND5xp2_ASAP7_75t_SL \i48/i146  (.A(\i48/n176 ),
    .B(\i48/n85 ),
    .C(\i48/n538 ),
    .D(\i48/n164 ),
    .E(\i48/n163 ),
    .Y(\i48/n314 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i48/i147  (.A1(\i48/n61 ),
    .A2(\i48/n75 ),
    .B(\i48/n549 ),
    .C(\i48/n233 ),
    .Y(\i48/n313 ));
 NAND4xp25_ASAP7_75t_SL \i48/i148  (.A(\i48/n268 ),
    .B(\i48/n214 ),
    .C(\i48/n90 ),
    .D(\i48/n528 ),
    .Y(\i48/n312 ));
 NAND5xp2_ASAP7_75t_SL \i48/i149  (.A(\i48/n140 ),
    .B(\i48/n527 ),
    .C(\i48/n206 ),
    .D(\i48/n87 ),
    .E(\i48/n83 ),
    .Y(\i48/n311 ));
 NOR3xp33_ASAP7_75t_SL \i48/i15  (.A(\i48/n450 ),
    .B(\i48/n392 ),
    .C(\i48/n434 ),
    .Y(\i48/n446 ));
 NAND2xp5_ASAP7_75t_SL \i48/i150  (.A(\i48/n238 ),
    .B(\i48/n260 ),
    .Y(\i48/n310 ));
 NAND3xp33_ASAP7_75t_SL \i48/i151  (.A(\i48/n255 ),
    .B(\i48/n461 ),
    .C(\i48/n77 ),
    .Y(\i48/n309 ));
 NAND2xp5_ASAP7_75t_SL \i48/i152  (.A(\i48/n499 ),
    .B(\i48/n474 ),
    .Y(\i48/n308 ));
 NOR2xp33_ASAP7_75t_L \i48/i153  (.A(\i48/n281 ),
    .B(\i48/n292 ),
    .Y(\i48/n331 ));
 NAND2xp5_ASAP7_75t_SL \i48/i154  (.A(\i48/n496 ),
    .B(\i48/n301 ),
    .Y(\i48/n307 ));
 NOR2x1p5_ASAP7_75t_SL \i48/i155  (.A(\i48/n481 ),
    .B(\i48/n284 ),
    .Y(\i48/n329 ));
 NAND3x1_ASAP7_75t_SL \i48/i156  (.A(\i48/n228 ),
    .B(\i48/n501 ),
    .C(\i48/n124 ),
    .Y(\i48/n23 ));
 INVxp67_ASAP7_75t_SL \i48/i157  (.A(\i48/n305 ),
    .Y(\i48/n306 ));
 INVxp67_ASAP7_75t_SL \i48/i158  (.A(\i48/n7 ),
    .Y(\i48/n304 ));
 INVxp67_ASAP7_75t_SL \i48/i159  (.A(\i48/n299 ),
    .Y(\i48/n300 ));
 NAND4xp75_ASAP7_75t_SL \i48/i16  (.A(\i48/n407 ),
    .B(\i48/n436 ),
    .C(\i48/n412 ),
    .D(\i48/n402 ),
    .Y(\i48/n445 ));
 INVxp67_ASAP7_75t_SL \i48/i160  (.A(\i48/n297 ),
    .Y(\i48/n298 ));
 INVx2_ASAP7_75t_SL \i48/i161  (.A(\i48/n295 ),
    .Y(\i48/n296 ));
 INVxp67_ASAP7_75t_SL \i48/i162  (.A(\i48/n486 ),
    .Y(\i48/n294 ));
 INVxp67_ASAP7_75t_SL \i48/i163  (.A(\i48/n290 ),
    .Y(\i48/n291 ));
 INVxp67_ASAP7_75t_SL \i48/i164  (.A(\i48/n512 ),
    .Y(\i48/n288 ));
 INVx1_ASAP7_75t_SL \i48/i165  (.A(\i48/n285 ),
    .Y(\i48/n286 ));
 NAND2x1_ASAP7_75t_SL \i48/i166  (.A(\i48/n189 ),
    .B(\i48/n188 ),
    .Y(\i48/n284 ));
 NOR2xp33_ASAP7_75t_SL \i48/i167  (.A(\i48/n558 ),
    .B(\i48/n219 ),
    .Y(\i48/n283 ));
 NAND2xp33_ASAP7_75t_SL \i48/i168  (.A(\i48/n539 ),
    .B(\i48/n495 ),
    .Y(\i48/n282 ));
 NAND2xp5_ASAP7_75t_SL \i48/i169  (.A(\i48/n150 ),
    .B(\i48/n539 ),
    .Y(\i48/n281 ));
 AND3x4_ASAP7_75t_SL \i48/i17  (.A(\i48/n427 ),
    .B(\i48/n442 ),
    .C(\i48/n432 ),
    .Y(n24[7]));
 AOI31xp33_ASAP7_75t_SL \i48/i170  (.A1(\i48/n42 ),
    .A2(\i48/n15 ),
    .A3(\i48/n484 ),
    .B(\i48/n35 ),
    .Y(\i48/n280 ));
 NOR3xp33_ASAP7_75t_SL \i48/i171  (.A(\i48/n458 ),
    .B(\i48/n112 ),
    .C(\i48/n97 ),
    .Y(\i48/n279 ));
 NOR3xp33_ASAP7_75t_SL \i48/i172  (.A(\i48/n504 ),
    .B(\i48/n105 ),
    .C(\i48/n558 ),
    .Y(\i48/n278 ));
 OAI31xp33_ASAP7_75t_SL \i48/i173  (.A1(\i48/n37 ),
    .A2(\i48/n39 ),
    .A3(\i48/n53 ),
    .B(\i48/n68 ),
    .Y(\i48/n277 ));
 AOI221xp5_ASAP7_75t_SL \i48/i174  (.A1(\i48/n61 ),
    .A2(\i48/n71 ),
    .B1(\i48/n511 ),
    .B2(\i48/n49 ),
    .C(\i48/n166 ),
    .Y(\i48/n276 ));
 OAI31xp33_ASAP7_75t_SL \i48/i175  (.A1(\i48/n57 ),
    .A2(\i48/n59 ),
    .A3(\i48/n61 ),
    .B(\i48/n53 ),
    .Y(\i48/n275 ));
 AOI21xp5_ASAP7_75t_SL \i48/i176  (.A1(\i48/n136 ),
    .A2(\i48/n484 ),
    .B(\i48/n67 ),
    .Y(\i48/n305 ));
 OAI221xp5_ASAP7_75t_SL \i48/i177  (.A1(\i48/n16 ),
    .A2(\i48/n70 ),
    .B1(\i48/n38 ),
    .B2(\i48/n45 ),
    .C(\i48/n185 ),
    .Y(\i48/n274 ));
 AOI21xp33_ASAP7_75t_SL \i48/i178  (.A1(\i48/n145 ),
    .A2(\i48/n36 ),
    .B(\i48/n60 ),
    .Y(\i48/n273 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i48/i179  (.A1(\i48/n546 ),
    .A2(\i48/n5 ),
    .B(\i48/n559 ),
    .C(\i48/n557 ),
    .Y(\i48/n272 ));
 NAND4xp75_ASAP7_75t_SL \i48/i18  (.A(\i48/n391 ),
    .B(\i48/n411 ),
    .C(\i48/n420 ),
    .D(\i48/n435 ),
    .Y(\i48/n444 ));
 NOR3xp33_ASAP7_75t_SL \i48/i180  (.A(\i48/n196 ),
    .B(\i48/n504 ),
    .C(\i48/n117 ),
    .Y(\i48/n271 ));
 NAND3xp33_ASAP7_75t_SL \i48/i181  (.A(\i48/n17 ),
    .B(\i48/n490 ),
    .C(\i48/n471 ),
    .Y(\i48/n270 ));
 AOI22xp5_ASAP7_75t_SL \i48/i182  (.A1(\i48/n457 ),
    .A2(\i48/n131 ),
    .B1(\i48/n49 ),
    .B2(\i48/n470 ),
    .Y(\i48/n269 ));
 OAI21xp5_ASAP7_75t_SL \i48/i183  (.A1(\i48/n48 ),
    .A2(\i48/n137 ),
    .B(\i48/n57 ),
    .Y(\i48/n268 ));
 NAND4xp25_ASAP7_75t_SL \i48/i184  (.A(\i48/n153 ),
    .B(\i48/n528 ),
    .C(\i48/n122 ),
    .D(\i48/n125 ),
    .Y(\i48/n267 ));
 NAND2xp33_ASAP7_75t_SL \i48/i185  (.A(\i48/n472 ),
    .B(\i48/n116 ),
    .Y(\i48/n266 ));
 OAI211xp5_ASAP7_75t_SL \i48/i186  (.A1(\i48/n60 ),
    .A2(\i48/n51 ),
    .B(\i48/n127 ),
    .C(\i48/n130 ),
    .Y(\i48/n303 ));
 NOR2x1_ASAP7_75t_SL \i48/i187  (.A(\i48/n135 ),
    .B(\i48/n518 ),
    .Y(\i48/n302 ));
 NOR2xp67_ASAP7_75t_SL \i48/i188  (.A(\i48/n515 ),
    .B(\i48/n225 ),
    .Y(\i48/n301 ));
 NAND2xp5_ASAP7_75t_SL \i48/i189  (.A(\i48/n210 ),
    .B(\i48/n497 ),
    .Y(\i48/n22 ));
 NAND2x1_ASAP7_75t_SL \i48/i19  (.A(\i48/n399 ),
    .B(\i48/n428 ),
    .Y(\i48/n443 ));
 NOR2xp33_ASAP7_75t_SL \i48/i190  (.A(\i48/n211 ),
    .B(\i48/n226 ),
    .Y(\i48/n299 ));
 OAI211xp5_ASAP7_75t_SL \i48/i191  (.A1(\i48/n484 ),
    .A2(\i48/n60 ),
    .B(\i48/n161 ),
    .C(\i48/n162 ),
    .Y(\i48/n297 ));
 OR2x2_ASAP7_75t_SL \i48/i192  (.A(\i48/n464 ),
    .B(\i48/n517 ),
    .Y(\i48/n295 ));
 OAI211xp5_ASAP7_75t_SL \i48/i193  (.A1(\i48/n70 ),
    .A2(\i48/n63 ),
    .B(\i48/n157 ),
    .C(\i48/n107 ),
    .Y(\i48/n293 ));
 NAND2xp5_ASAP7_75t_SL \i48/i194  (.A(\i48/n523 ),
    .B(\i48/n526 ),
    .Y(\i48/n292 ));
 NAND2xp5_ASAP7_75t_SL \i48/i195  (.A(\i48/n20 ),
    .B(\i48/n168 ),
    .Y(\i48/n290 ));
 NAND2xp5_ASAP7_75t_SL \i48/i196  (.A(\i48/n208 ),
    .B(\i48/n568 ),
    .Y(\i48/n289 ));
 NAND2xp5_ASAP7_75t_SL \i48/i197  (.A(\i48/n155 ),
    .B(\i48/n573 ),
    .Y(\i48/n287 ));
 NOR2x1_ASAP7_75t_SL \i48/i198  (.A(\i48/n209 ),
    .B(\i48/n184 ),
    .Y(\i48/n285 ));
 INVxp67_ASAP7_75t_SL \i48/i199  (.A(\i48/n261 ),
    .Y(\i48/n262 ));
 INVx2_ASAP7_75t_SL \i48/i2  (.A(n25[2]),
    .Y(\i48/n2 ));
 NOR2xp67_ASAP7_75t_SL \i48/i20  (.A(\i48/n393 ),
    .B(\i48/n429 ),
    .Y(\i48/n442 ));
 INVx1_ASAP7_75t_SL \i48/i200  (.A(\i48/n258 ),
    .Y(\i48/n259 ));
 INVx1_ASAP7_75t_SL \i48/i201  (.A(\i48/n255 ),
    .Y(\i48/n256 ));
 NAND4xp25_ASAP7_75t_SL \i48/i202  (.A(\i48/n534 ),
    .B(\i48/n108 ),
    .C(\i48/n94 ),
    .D(\i48/n565 ),
    .Y(\i48/n252 ));
 AOI31xp33_ASAP7_75t_SL \i48/i203  (.A1(\i48/n109 ),
    .A2(\i48/n56 ),
    .A3(\i48/n35 ),
    .B(\i48/n36 ),
    .Y(\i48/n251 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i48/i204  (.A1(\i48/n559 ),
    .A2(\i48/n41 ),
    .B(\i48/n53 ),
    .C(\i48/n113 ),
    .Y(\i48/n250 ));
 NOR4xp25_ASAP7_75t_SL \i48/i205  (.A(\i48/n89 ),
    .B(\i48/n462 ),
    .C(\i48/n160 ),
    .D(\i48/n72 ),
    .Y(\i48/n249 ));
 AOI211xp5_ASAP7_75t_SL \i48/i206  (.A1(\i48/n110 ),
    .A2(\i48/n548 ),
    .B(\i48/n149 ),
    .C(\i48/n78 ),
    .Y(\i48/n248 ));
 AOI21xp5_ASAP7_75t_R \i48/i207  (.A1(\i48/n530 ),
    .A2(\i48/n559 ),
    .B(\i48/n201 ),
    .Y(\i48/n247 ));
 NOR2xp33_ASAP7_75t_L \i48/i208  (.A(\i48/n510 ),
    .B(\i48/n220 ),
    .Y(\i48/n246 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i48/i209  (.A1(\i48/n60 ),
    .A2(\i48/n40 ),
    .B(\i48/n66 ),
    .C(\i48/n197 ),
    .Y(\i48/n245 ));
 NAND4xp75_ASAP7_75t_SL \i48/i21  (.A(\i48/n403 ),
    .B(\i48/n415 ),
    .C(\i48/n397 ),
    .D(\i48/n400 ),
    .Y(\i48/n441 ));
 OAI22xp5_ASAP7_75t_SL \i48/i210  (.A1(\i48/n63 ),
    .A2(\i48/n138 ),
    .B1(\i48/n51 ),
    .B2(\i48/n76 ),
    .Y(\i48/n244 ));
 NOR2xp33_ASAP7_75t_SL \i48/i211  (.A(\i48/n181 ),
    .B(\i48/n169 ),
    .Y(\i48/n243 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i48/i212  (.A1(\i48/n457 ),
    .A2(\i48/n46 ),
    .B(\i48/n5 ),
    .C(\i48/n146 ),
    .Y(\i48/n242 ));
 NAND2xp33_ASAP7_75t_L \i48/i213  (.A(\i48/n543 ),
    .B(\i48/n536 ),
    .Y(\i48/n241 ));
 NAND2xp33_ASAP7_75t_SL \i48/i214  (.A(\i48/n473 ),
    .B(\i48/n106 ),
    .Y(\i48/n240 ));
 AOI22xp5_ASAP7_75t_SL \i48/i215  (.A1(\i48/n59 ),
    .A2(\i48/n86 ),
    .B1(\i48/n548 ),
    .B2(\i48/n61 ),
    .Y(\i48/n239 ));
 OAI21xp33_ASAP7_75t_SL \i48/i216  (.A1(\i48/n93 ),
    .A2(\i48/n59 ),
    .B(\i48/n548 ),
    .Y(\i48/n238 ));
 NAND4xp25_ASAP7_75t_SL \i48/i217  (.A(\i48/n103 ),
    .B(\i48/n126 ),
    .C(\i48/n84 ),
    .D(\i48/n82 ),
    .Y(\i48/n237 ));
 AOI221xp5_ASAP7_75t_SL \i48/i218  (.A1(\i48/n49 ),
    .A2(\i48/n34 ),
    .B1(\i48/n41 ),
    .B2(\i48/n50 ),
    .C(\i48/n518 ),
    .Y(\i48/n236 ));
 OAI221xp5_ASAP7_75t_SL \i48/i219  (.A1(\i48/n69 ),
    .A2(\i48/n66 ),
    .B1(\i48/n54 ),
    .B2(\i48/n552 ),
    .C(\i48/n88 ),
    .Y(\i48/n265 ));
 OR3x1_ASAP7_75t_SL \i48/i22  (.A(\i48/n423 ),
    .B(\i48/n421 ),
    .C(\i48/n404 ),
    .Y(\i48/n440 ));
 OAI222xp33_ASAP7_75t_SL \i48/i220  (.A1(\i48/n564 ),
    .A2(\i48/n42 ),
    .B1(\i48/n45 ),
    .B2(\i48/n51 ),
    .C1(\i48/n54 ),
    .C2(\i48/n62 ),
    .Y(\i48/n235 ));
 AND3x1_ASAP7_75t_SL \i48/i221  (.A(\i48/n100 ),
    .B(\i48/n108 ),
    .C(\i48/n203 ),
    .Y(\i48/n234 ));
 AOI22xp5_ASAP7_75t_SL \i48/i222  (.A1(\i48/n478 ),
    .A2(\i48/n133 ),
    .B1(\i48/n48 ),
    .B2(\i48/n559 ),
    .Y(\i48/n264 ));
 NAND2xp33_ASAP7_75t_SL \i48/i223  (.A(\i48/n172 ),
    .B(\i48/n204 ),
    .Y(\i48/n233 ));
 OAI222xp33_ASAP7_75t_SL \i48/i224  (.A1(\i48/n63 ),
    .A2(\i48/n64 ),
    .B1(\i48/n69 ),
    .B2(\i48/n62 ),
    .C1(\i48/n16 ),
    .C2(\i48/n484 ),
    .Y(\i48/n263 ));
 NAND3x1_ASAP7_75t_SL \i48/i225  (.A(\i48/n537 ),
    .B(\i48/n128 ),
    .C(\i48/n123 ),
    .Y(\i48/n261 ));
 AOI22x1_ASAP7_75t_SL \i48/i226  (.A1(\i48/n553 ),
    .A2(\i48/n68 ),
    .B1(\i48/n511 ),
    .B2(\i48/n53 ),
    .Y(\i48/n12 ));
 AOI22xp5_ASAP7_75t_SL \i48/i227  (.A1(\i48/n71 ),
    .A2(\i48/n469 ),
    .B1(\i48/n37 ),
    .B2(\i48/n57 ),
    .Y(\i48/n260 ));
 AOI221xp5_ASAP7_75t_SL \i48/i228  (.A1(\i48/n68 ),
    .A2(\i48/n53 ),
    .B1(\i48/n61 ),
    .B2(\i48/n549 ),
    .C(\i48/n205 ),
    .Y(\i48/n258 ));
 OAI21xp33_ASAP7_75t_SL \i48/i229  (.A1(\i48/n35 ),
    .A2(\i48/n66 ),
    .B(\i48/n212 ),
    .Y(\i48/n257 ));
 OR3x1_ASAP7_75t_SL \i48/i23  (.A(\i48/n424 ),
    .B(\i48/n390 ),
    .C(\i48/n363 ),
    .Y(\i48/n439 ));
 NOR2x1_ASAP7_75t_SL \i48/i230  (.A(\i48/n102 ),
    .B(\i48/n171 ),
    .Y(\i48/n255 ));
 OAI211xp5_ASAP7_75t_SL \i48/i231  (.A1(\i48/n52 ),
    .A2(\i48/n572 ),
    .B(\i48/n90 ),
    .C(\i48/n567 ),
    .Y(\i48/n254 ));
 NOR2xp33_ASAP7_75t_SL \i48/i232  (.A(\i48/n113 ),
    .B(\i48/n175 ),
    .Y(\i48/n21 ));
 NOR2xp33_ASAP7_75t_SL \i48/i233  (.A(\i48/n114 ),
    .B(\i48/n227 ),
    .Y(\i48/n232 ));
 AOI222xp33_ASAP7_75t_SL \i48/i234  (.A1(\i48/n61 ),
    .A2(\i48/n49 ),
    .B1(\i48/n5 ),
    .B2(\i48/n34 ),
    .C1(\i48/n57 ),
    .C2(\i48/n48 ),
    .Y(\i48/n253 ));
 INVx1_ASAP7_75t_R \i48/i235  (.A(\i48/n568 ),
    .Y(\i48/n230 ));
 INVx1_ASAP7_75t_SL \i48/i236  (.A(\i48/n227 ),
    .Y(\i48/n228 ));
 INVxp67_ASAP7_75t_SL \i48/i237  (.A(\i48/n223 ),
    .Y(\i48/n224 ));
 INVx1_ASAP7_75t_SL \i48/i238  (.A(\i48/n220 ),
    .Y(\i48/n221 ));
 OAI21xp33_ASAP7_75t_SL \i48/i239  (.A1(\i48/n58 ),
    .A2(\i48/n47 ),
    .B(\i48/n487 ),
    .Y(\i48/n218 ));
 NAND3xp33_ASAP7_75t_SL \i48/i24  (.A(\i48/n433 ),
    .B(\i48/n420 ),
    .C(\i48/n403 ),
    .Y(\i48/n438 ));
 NAND2xp5_ASAP7_75t_SL \i48/i240  (.A(\i48/n569 ),
    .B(\i48/n107 ),
    .Y(\i48/n217 ));
 NOR2xp33_ASAP7_75t_SL \i48/i241  (.A(\i48/n115 ),
    .B(\i48/n148 ),
    .Y(\i48/n216 ));
 NAND2xp33_ASAP7_75t_L \i48/i242  (.A(\i48/n571 ),
    .B(\i48/n79 ),
    .Y(\i48/n215 ));
 OAI21xp5_ASAP7_75t_SL \i48/i243  (.A1(\i48/n55 ),
    .A2(\i48/n46 ),
    .B(\i48/n39 ),
    .Y(\i48/n214 ));
 NOR2xp33_ASAP7_75t_SL \i48/i244  (.A(\i48/n557 ),
    .B(\i48/n95 ),
    .Y(\i48/n213 ));
 OAI21xp5_ASAP7_75t_SL \i48/i245  (.A1(\i48/n59 ),
    .A2(\i48/n65 ),
    .B(\i48/n49 ),
    .Y(\i48/n212 ));
 OAI21xp5_ASAP7_75t_SL \i48/i246  (.A1(\i48/n535 ),
    .A2(\i48/n67 ),
    .B(\i48/n529 ),
    .Y(\i48/n211 ));
 AOI22xp5_ASAP7_75t_SL \i48/i247  (.A1(\i48/n546 ),
    .A2(\i48/n46 ),
    .B1(\i48/n549 ),
    .B2(\i48/n57 ),
    .Y(\i48/n210 ));
 OAI21xp5_ASAP7_75t_SL \i48/i248  (.A1(\i48/n15 ),
    .A2(\i48/n54 ),
    .B(\i48/n111 ),
    .Y(\i48/n209 ));
 AOI22xp5_ASAP7_75t_SL \i48/i249  (.A1(\i48/n34 ),
    .A2(\i48/n71 ),
    .B1(\i48/n37 ),
    .B2(\i48/n59 ),
    .Y(\i48/n208 ));
 NOR2x1_ASAP7_75t_SL \i48/i25  (.A(\i48/n345 ),
    .B(\i48/n421 ),
    .Y(\i48/n436 ));
 OA21x2_ASAP7_75t_SL \i48/i250  (.A1(\i48/n524 ),
    .A2(\i48/n44 ),
    .B(\i48/n488 ),
    .Y(\i48/n231 ));
 AOI21xp33_ASAP7_75t_SL \i48/i251  (.A1(\i48/n51 ),
    .A2(\i48/n524 ),
    .B(\i48/n35 ),
    .Y(\i48/n207 ));
 OAI21xp5_ASAP7_75t_SL \i48/i252  (.A1(\i48/n549 ),
    .A2(\i48/n71 ),
    .B(\i48/n478 ),
    .Y(\i48/n206 ));
 OA21x2_ASAP7_75t_SL \i48/i253  (.A1(\i48/n5 ),
    .A2(\i48/n71 ),
    .B(\i48/n559 ),
    .Y(\i48/n205 ));
 OAI21xp5_ASAP7_75t_SL \i48/i254  (.A1(\i48/n50 ),
    .A2(\i48/n37 ),
    .B(\i48/n478 ),
    .Y(\i48/n204 ));
 OAI21xp5_ASAP7_75t_SL \i48/i255  (.A1(\i48/n59 ),
    .A2(\i48/n55 ),
    .B(\i48/n71 ),
    .Y(\i48/n203 ));
 AOI21xp33_ASAP7_75t_SL \i48/i256  (.A1(\i48/n484 ),
    .A2(\i48/n66 ),
    .B(\i48/n35 ),
    .Y(\i48/n202 ));
 OAI21xp5_ASAP7_75t_SL \i48/i257  (.A1(\i48/n535 ),
    .A2(\i48/n54 ),
    .B(\i48/n19 ),
    .Y(\i48/n201 ));
 AOI22xp5_ASAP7_75t_SL \i48/i258  (.A1(\i48/n48 ),
    .A2(\i48/n457 ),
    .B1(\i48/n549 ),
    .B2(\i48/n46 ),
    .Y(\i48/n200 ));
 AOI21xp33_ASAP7_75t_SL \i48/i259  (.A1(\i48/n60 ),
    .A2(\i48/n35 ),
    .B(\i48/n52 ),
    .Y(\i48/n199 ));
 NOR2x1_ASAP7_75t_SL \i48/i26  (.A(\i48/n405 ),
    .B(\i48/n401 ),
    .Y(\i48/n435 ));
 OAI21xp5_ASAP7_75t_SL \i48/i260  (.A1(\i48/n559 ),
    .A2(\i48/n59 ),
    .B(\i48/n39 ),
    .Y(\i48/n198 ));
 OAI21xp5_ASAP7_75t_SL \i48/i261  (.A1(\i48/n55 ),
    .A2(\i48/n457 ),
    .B(\i48/n549 ),
    .Y(\i48/n197 ));
 NAND2xp5_ASAP7_75t_SL \i48/i262  (.A(\i48/n478 ),
    .B(\i48/n530 ),
    .Y(\i48/n20 ));
 NAND2xp5_ASAP7_75t_L \i48/i263  (.A(\i48/n161 ),
    .B(\i48/n162 ),
    .Y(\i48/n196 ));
 OAI22xp5_ASAP7_75t_SL \i48/i264  (.A1(\i48/n498 ),
    .A2(\i48/n54 ),
    .B1(\i48/n16 ),
    .B2(\i48/n51 ),
    .Y(\i48/n229 ));
 OAI22xp5_ASAP7_75t_SL \i48/i265  (.A1(\i48/n70 ),
    .A2(\i48/n45 ),
    .B1(\i48/n535 ),
    .B2(\i48/n63 ),
    .Y(\i48/n227 ));
 OAI22xp5_ASAP7_75t_SL \i48/i266  (.A1(\i48/n52 ),
    .A2(\i48/n63 ),
    .B1(\i48/n54 ),
    .B2(\i48/n38 ),
    .Y(\i48/n226 ));
 OAI22xp5_ASAP7_75t_SL \i48/i267  (.A1(\i48/n498 ),
    .A2(\i48/n69 ),
    .B1(\i48/n36 ),
    .B2(\i48/n564 ),
    .Y(\i48/n225 ));
 OAI22xp5_ASAP7_75t_SL \i48/i268  (.A1(\i48/n535 ),
    .A2(\i48/n69 ),
    .B1(\i48/n51 ),
    .B2(\i48/n67 ),
    .Y(\i48/n223 ));
 OAI21xp5_ASAP7_75t_SL \i48/i269  (.A1(\i48/n59 ),
    .A2(\i48/n41 ),
    .B(\i48/n546 ),
    .Y(\i48/n222 ));
 NAND3xp33_ASAP7_75t_SL \i48/i27  (.A(\i48/n385 ),
    .B(\i48/n581 ),
    .C(\i48/n382 ),
    .Y(\i48/n434 ));
 NOR2xp33_ASAP7_75t_L \i48/i270  (.A(\i48/n44 ),
    .B(\i48/n491 ),
    .Y(\i48/n220 ));
 NAND2xp33_ASAP7_75t_L \i48/i271  (.A(\i48/n90 ),
    .B(\i48/n567 ),
    .Y(\i48/n195 ));
 OAI21xp5_ASAP7_75t_SL \i48/i272  (.A1(\i48/n52 ),
    .A2(\i48/n45 ),
    .B(\i48/n505 ),
    .Y(\i48/n219 ));
 INVxp67_ASAP7_75t_SL \i48/i273  (.A(\i48/n193 ),
    .Y(\i48/n194 ));
 INVxp67_ASAP7_75t_SL \i48/i274  (.A(\i48/n191 ),
    .Y(\i48/n192 ));
 INVx1_ASAP7_75t_SL \i48/i275  (.A(\i48/n189 ),
    .Y(\i48/n190 ));
 INVx1_ASAP7_75t_SL \i48/i276  (.A(\i48/n187 ),
    .Y(\i48/n188 ));
 INVxp67_ASAP7_75t_SL \i48/i277  (.A(\i48/n185 ),
    .Y(\i48/n186 ));
 INVxp67_ASAP7_75t_SL \i48/i278  (.A(\i48/n181 ),
    .Y(\i48/n182 ));
 INVxp67_ASAP7_75t_SL \i48/i279  (.A(\i48/n179 ),
    .Y(\i48/n180 ));
 NOR2xp33_ASAP7_75t_L \i48/i28  (.A(\i48/n410 ),
    .B(\i48/n372 ),
    .Y(\i48/n433 ));
 OAI21xp5_ASAP7_75t_SL \i48/i280  (.A1(\i48/n46 ),
    .A2(\i48/n560 ),
    .B(\i48/n549 ),
    .Y(\i48/n176 ));
 OAI22xp5_ASAP7_75t_SL \i48/i281  (.A1(\i48/n69 ),
    .A2(\i48/n42 ),
    .B1(\i48/n38 ),
    .B2(\i48/n44 ),
    .Y(\i48/n175 ));
 AOI21xp33_ASAP7_75t_SL \i48/i282  (.A1(\i48/n54 ),
    .A2(\i48/n63 ),
    .B(\i48/n64 ),
    .Y(\i48/n174 ));
 AO21x1_ASAP7_75t_SL \i48/i283  (.A1(\i48/n34 ),
    .A2(\i48/n53 ),
    .B(\i48/n503 ),
    .Y(\i48/n173 ));
 OAI21xp5_ASAP7_75t_SL \i48/i284  (.A1(\i48/n34 ),
    .A2(\i48/n41 ),
    .B(\i48/n39 ),
    .Y(\i48/n172 ));
 OAI22xp33_ASAP7_75t_SL \i48/i285  (.A1(\i48/n16 ),
    .A2(\i48/n47 ),
    .B1(\i48/n63 ),
    .B2(\i48/n66 ),
    .Y(\i48/n171 ));
 OAI22xp5_ASAP7_75t_SL \i48/i286  (.A1(\i48/n484 ),
    .A2(\i48/n564 ),
    .B1(\i48/n66 ),
    .B2(\i48/n60 ),
    .Y(\i48/n170 ));
 OAI22xp33_ASAP7_75t_SL \i48/i287  (.A1(\i48/n40 ),
    .A2(\i48/n47 ),
    .B1(\i48/n44 ),
    .B2(\i48/n42 ),
    .Y(\i48/n169 ));
 AOI22xp5_ASAP7_75t_SL \i48/i288  (.A1(\i48/n49 ),
    .A2(\i48/n560 ),
    .B1(\i48/n37 ),
    .B2(\i48/n65 ),
    .Y(\i48/n168 ));
 OAI22xp5_ASAP7_75t_SL \i48/i289  (.A1(\i48/n47 ),
    .A2(\i48/n69 ),
    .B1(\i48/n51 ),
    .B2(\i48/n44 ),
    .Y(\i48/n167 ));
 NOR5xp2_ASAP7_75t_SL \i48/i29  (.A(\i48/n374 ),
    .B(\i48/n323 ),
    .C(\i48/n365 ),
    .D(\i48/n289 ),
    .E(\i48/n293 ),
    .Y(\i48/n432 ));
 OAI21xp5_ASAP7_75t_SL \i48/i290  (.A1(\i48/n36 ),
    .A2(\i48/n45 ),
    .B(\i48/n96 ),
    .Y(\i48/n193 ));
 AOI22xp5_ASAP7_75t_SL \i48/i291  (.A1(\i48/n34 ),
    .A2(\i48/n50 ),
    .B1(\i48/n37 ),
    .B2(\i48/n470 ),
    .Y(\i48/n191 ));
 AOI22xp5_ASAP7_75t_SL \i48/i292  (.A1(\i48/n39 ),
    .A2(\i48/n41 ),
    .B1(\i48/n457 ),
    .B2(\i48/n49 ),
    .Y(\i48/n189 ));
 OAI22xp5_ASAP7_75t_R \i48/i293  (.A1(\i48/n35 ),
    .A2(\i48/n552 ),
    .B1(\i48/n47 ),
    .B2(\i48/n56 ),
    .Y(\i48/n166 ));
 NAND2xp33_ASAP7_75t_SL \i48/i294  (.A(\i48/n163 ),
    .B(\i48/n164 ),
    .Y(\i48/n165 ));
 OAI22x1_ASAP7_75t_SL \i48/i295  (.A1(\i48/n15 ),
    .A2(\i48/n69 ),
    .B1(\i48/n38 ),
    .B2(\i48/n58 ),
    .Y(\i48/n187 ));
 AOI22xp5_ASAP7_75t_SL \i48/i296  (.A1(\i48/n39 ),
    .A2(\i48/n457 ),
    .B1(\i48/n37 ),
    .B2(\i48/n559 ),
    .Y(\i48/n185 ));
 AO22x2_ASAP7_75t_SL \i48/i297  (.A1(\i48/n71 ),
    .A2(\i48/n68 ),
    .B1(\i48/n43 ),
    .B2(\i48/n65 ),
    .Y(\i48/n184 ));
 OAI21xp5_ASAP7_75t_SL \i48/i298  (.A1(\i48/n62 ),
    .A2(\i48/n40 ),
    .B(\i48/n541 ),
    .Y(\i48/n183 ));
 OAI22xp33_ASAP7_75t_SL \i48/i299  (.A1(\i48/n64 ),
    .A2(\i48/n35 ),
    .B1(\i48/n36 ),
    .B2(\i48/n63 ),
    .Y(\i48/n181 ));
 INVx2_ASAP7_75t_SL \i48/i3  (.A(\i48/n506 ),
    .Y(\i48/n3 ));
 NOR3xp33_ASAP7_75t_SL \i48/i30  (.A(\i48/n370 ),
    .B(\i48/n387 ),
    .C(\i48/n419 ),
    .Y(\i48/n431 ));
 OAI22xp5_ASAP7_75t_SL \i48/i300  (.A1(\i48/n484 ),
    .A2(\i48/n40 ),
    .B1(\i48/n51 ),
    .B2(\i48/n63 ),
    .Y(\i48/n179 ));
 AOI22xp5_ASAP7_75t_SL \i48/i301  (.A1(\i48/n34 ),
    .A2(\i48/n39 ),
    .B1(\i48/n53 ),
    .B2(\i48/n65 ),
    .Y(\i48/n178 ));
 OAI22x1_ASAP7_75t_SL \i48/i302  (.A1(\i48/n60 ),
    .A2(\i48/n47 ),
    .B1(\i48/n56 ),
    .B2(\i48/n524 ),
    .Y(\i48/n177 ));
 INVxp67_ASAP7_75t_SL \i48/i303  (.A(\i48/n158 ),
    .Y(\i48/n159 ));
 INVx1_ASAP7_75t_SL \i48/i304  (.A(\i48/n500 ),
    .Y(\i48/n157 ));
 INVxp67_ASAP7_75t_SL \i48/i305  (.A(\i48/n155 ),
    .Y(\i48/n156 ));
 INVxp67_ASAP7_75t_SL \i48/i306  (.A(\i48/n153 ),
    .Y(\i48/n154 ));
 INVxp67_ASAP7_75t_SL \i48/i307  (.A(\i48/n487 ),
    .Y(\i48/n152 ));
 INVxp67_ASAP7_75t_R \i48/i308  (.A(\i48/n519 ),
    .Y(\i48/n150 ));
 INVxp67_ASAP7_75t_SL \i48/i309  (.A(\i48/n529 ),
    .Y(\i48/n147 ));
 NOR2x1_ASAP7_75t_SL \i48/i31  (.A(\i48/n416 ),
    .B(\i48/n375 ),
    .Y(\i48/n430 ));
 INVxp67_ASAP7_75t_SL \i48/i310  (.A(\i48/n571 ),
    .Y(\i48/n146 ));
 INVxp67_ASAP7_75t_SL \i48/i311  (.A(\i48/n471 ),
    .Y(\i48/n144 ));
 INVxp67_ASAP7_75t_SL \i48/i312  (.A(\i48/n142 ),
    .Y(\i48/n143 ));
 INVxp67_ASAP7_75t_SL \i48/i313  (.A(\i48/n140 ),
    .Y(\i48/n141 ));
 INVxp67_ASAP7_75t_SL \i48/i314  (.A(\i48/n138 ),
    .Y(\i48/n139 ));
 INVxp67_ASAP7_75t_SL \i48/i315  (.A(\i48/n491 ),
    .Y(\i48/n137 ));
 INVx1_ASAP7_75t_SL \i48/i316  (.A(\i48/n530 ),
    .Y(\i48/n136 ));
 NAND2xp5_ASAP7_75t_SL \i48/i317  (.A(\i48/n50 ),
    .B(\i48/n478 ),
    .Y(\i48/n164 ));
 AND2x2_ASAP7_75t_SL \i48/i318  (.A(\i48/n43 ),
    .B(\i48/n57 ),
    .Y(\i48/n135 ));
 NAND2xp5_ASAP7_75t_SL \i48/i319  (.A(\i48/n546 ),
    .B(\i48/n65 ),
    .Y(\i48/n134 ));
 NAND2xp5_ASAP7_75t_SL \i48/i32  (.A(\i48/n373 ),
    .B(\i48/n394 ),
    .Y(\i48/n429 ));
 NAND2xp5_ASAP7_75t_SL \i48/i320  (.A(\i48/n66 ),
    .B(\i48/n64 ),
    .Y(\i48/n133 ));
 NAND2xp5_ASAP7_75t_SL \i48/i321  (.A(\i48/n37 ),
    .B(\i48/n68 ),
    .Y(\i48/n132 ));
 NAND2xp33_ASAP7_75t_SL \i48/i322  (.A(\i48/n484 ),
    .B(\i48/n535 ),
    .Y(\i48/n131 ));
 NAND2xp5_ASAP7_75t_SL \i48/i323  (.A(\i48/n46 ),
    .B(\i48/n48 ),
    .Y(\i48/n130 ));
 NAND2xp5_ASAP7_75t_SL \i48/i324  (.A(\i48/n46 ),
    .B(\i48/n49 ),
    .Y(\i48/n163 ));
 NAND2xp5_ASAP7_75t_SL \i48/i325  (.A(\i48/n48 ),
    .B(\i48/n55 ),
    .Y(\i48/n162 ));
 NAND2xp5_ASAP7_75t_SL \i48/i326  (.A(\i48/n49 ),
    .B(\i48/n478 ),
    .Y(\i48/n129 ));
 NAND2xp5_ASAP7_75t_SL \i48/i327  (.A(\i48/n4 ),
    .B(\i48/n48 ),
    .Y(\i48/n128 ));
 NAND2xp5_ASAP7_75t_SL \i48/i328  (.A(\i48/n559 ),
    .B(\i48/n546 ),
    .Y(\i48/n127 ));
 NAND2xp5_ASAP7_75t_SL \i48/i329  (.A(\i48/n50 ),
    .B(\i48/n4 ),
    .Y(\i48/n126 ));
 NOR3x1_ASAP7_75t_SL \i48/i33  (.A(\i48/n23 ),
    .B(\i48/n389 ),
    .C(\i48/n315 ),
    .Y(\i48/n437 ));
 NAND2xp5_ASAP7_75t_SL \i48/i330  (.A(\i48/n57 ),
    .B(\i48/n53 ),
    .Y(\i48/n125 ));
 NAND2xp5_ASAP7_75t_SL \i48/i331  (.A(\i48/n49 ),
    .B(\i48/n57 ),
    .Y(\i48/n124 ));
 NAND2xp5_ASAP7_75t_SL \i48/i332  (.A(\i48/n34 ),
    .B(\i48/n43 ),
    .Y(\i48/n123 ));
 NAND2xp5_ASAP7_75t_SL \i48/i333  (.A(\i48/n43 ),
    .B(\i48/n55 ),
    .Y(\i48/n122 ));
 NAND2xp5_ASAP7_75t_SL \i48/i334  (.A(\i48/n50 ),
    .B(\i48/n559 ),
    .Y(\i48/n121 ));
 NAND2xp5_ASAP7_75t_SL \i48/i335  (.A(\i48/n34 ),
    .B(\i48/n549 ),
    .Y(\i48/n161 ));
 AND2x2_ASAP7_75t_SL \i48/i336  (.A(\i48/n43 ),
    .B(\i48/n59 ),
    .Y(\i48/n160 ));
 AND2x2_ASAP7_75t_SL \i48/i337  (.A(\i48/n546 ),
    .B(\i48/n55 ),
    .Y(\i48/n158 ));
 NAND2xp5_ASAP7_75t_SL \i48/i338  (.A(\i48/n57 ),
    .B(\i48/n5 ),
    .Y(\i48/n19 ));
 NAND2xp5_ASAP7_75t_SL \i48/i339  (.A(\i48/n549 ),
    .B(\i48/n559 ),
    .Y(\i48/n155 ));
 NOR3xp33_ASAP7_75t_SL \i48/i34  (.A(\i48/n333 ),
    .B(\i48/n23 ),
    .C(\i48/n413 ),
    .Y(\i48/n427 ));
 NAND2xp5_ASAP7_75t_SL \i48/i340  (.A(\i48/n71 ),
    .B(\i48/n41 ),
    .Y(\i48/n153 ));
 AND2x2_ASAP7_75t_SL \i48/i341  (.A(\i48/n50 ),
    .B(\i48/n457 ),
    .Y(\i48/n151 ));
 NOR2xp67_ASAP7_75t_SL \i48/i342  (.A(\i48/n524 ),
    .B(\i48/n54 ),
    .Y(\i48/n18 ));
 NOR2xp33_ASAP7_75t_SL \i48/i343  (.A(\i48/n52 ),
    .B(\i48/n63 ),
    .Y(\i48/n120 ));
 NAND2xp5_ASAP7_75t_SL \i48/i344  (.A(\i48/n457 ),
    .B(\i48/n48 ),
    .Y(\i48/n119 ));
 NOR2xp33_ASAP7_75t_SL \i48/i345  (.A(\i48/n47 ),
    .B(\i48/n63 ),
    .Y(\i48/n149 ));
 AND2x2_ASAP7_75t_SL \i48/i346  (.A(\i48/n49 ),
    .B(\i48/n4 ),
    .Y(\i48/n148 ));
 NOR2xp33_ASAP7_75t_SL \i48/i347  (.A(\i48/n15 ),
    .B(\i48/n44 ),
    .Y(\i48/n118 ));
 NOR2xp33_ASAP7_75t_SL \i48/i348  (.A(\i48/n47 ),
    .B(\i48/n67 ),
    .Y(\i48/n117 ));
 NOR2xp33_ASAP7_75t_L \i48/i349  (.A(\i48/n71 ),
    .B(\i48/n39 ),
    .Y(\i48/n145 ));
 NOR2xp67_ASAP7_75t_SL \i48/i35  (.A(\i48/n395 ),
    .B(\i48/n23 ),
    .Y(\i48/n426 ));
 NAND2xp5_ASAP7_75t_SL \i48/i350  (.A(\i48/n559 ),
    .B(\i48/n49 ),
    .Y(\i48/n142 ));
 NAND2xp5_ASAP7_75t_SL \i48/i351  (.A(\i48/n71 ),
    .B(\i48/n57 ),
    .Y(\i48/n140 ));
 NAND2xp5_ASAP7_75t_SL \i48/i352  (.A(\i48/n50 ),
    .B(\i48/n61 ),
    .Y(\i48/n116 ));
 NOR2xp33_ASAP7_75t_SL \i48/i353  (.A(\i48/n50 ),
    .B(\i48/n546 ),
    .Y(\i48/n138 ));
 NOR2xp33_ASAP7_75t_SL \i48/i354  (.A(\i48/n45 ),
    .B(\i48/n66 ),
    .Y(\i48/n115 ));
 INVxp67_ASAP7_75t_SL \i48/i355  (.A(\i48/n501 ),
    .Y(\i48/n114 ));
 INVxp67_ASAP7_75t_SL \i48/i356  (.A(\i48/n111 ),
    .Y(\i48/n112 ));
 INVx1_ASAP7_75t_SL \i48/i357  (.A(\i48/n109 ),
    .Y(\i48/n110 ));
 INVxp67_ASAP7_75t_SL \i48/i358  (.A(\i48/n103 ),
    .Y(\i48/n104 ));
 INVxp67_ASAP7_75t_SL \i48/i359  (.A(\i48/n101 ),
    .Y(\i48/n102 ));
 NOR3xp33_ASAP7_75t_SL \i48/i36  (.A(\i48/n371 ),
    .B(\i48/n366 ),
    .C(\i48/n8 ),
    .Y(\i48/n425 ));
 INVxp67_ASAP7_75t_SL \i48/i360  (.A(\i48/n462 ),
    .Y(\i48/n100 ));
 INVxp67_ASAP7_75t_SL \i48/i361  (.A(\i48/n98 ),
    .Y(\i48/n99 ));
 INVxp67_ASAP7_75t_SL \i48/i362  (.A(\i48/n502 ),
    .Y(\i48/n97 ));
 INVxp67_ASAP7_75t_SL \i48/i363  (.A(\i48/n95 ),
    .Y(\i48/n96 ));
 INVxp67_ASAP7_75t_SL \i48/i364  (.A(\i48/n534 ),
    .Y(\i48/n91 ));
 INVx1_ASAP7_75t_SL \i48/i365  (.A(\i48/n543 ),
    .Y(\i48/n89 ));
 NAND2xp5_ASAP7_75t_SL \i48/i366  (.A(\i48/n548 ),
    .B(\i48/n59 ),
    .Y(\i48/n88 ));
 NAND2xp5_ASAP7_75t_SL \i48/i367  (.A(\i48/n39 ),
    .B(\i48/n61 ),
    .Y(\i48/n87 ));
 NAND2xp5_ASAP7_75t_SL \i48/i368  (.A(\i48/n62 ),
    .B(\i48/n52 ),
    .Y(\i48/n86 ));
 NAND2xp5_ASAP7_75t_SL \i48/i369  (.A(\i48/n61 ),
    .B(\i48/n37 ),
    .Y(\i48/n85 ));
 NAND3xp33_ASAP7_75t_SL \i48/i37  (.A(\i48/n335 ),
    .B(\i48/n381 ),
    .C(\i48/n367 ),
    .Y(\i48/n424 ));
 NAND2xp5_ASAP7_75t_SL \i48/i370  (.A(\i48/n549 ),
    .B(\i48/n457 ),
    .Y(\i48/n84 ));
 NAND2xp5_ASAP7_75t_SL \i48/i371  (.A(\i48/n53 ),
    .B(\i48/n470 ),
    .Y(\i48/n83 ));
 NAND2xp5_ASAP7_75t_SL \i48/i372  (.A(\i48/n37 ),
    .B(\i48/n55 ),
    .Y(\i48/n82 ));
 NAND2xp5_ASAP7_75t_L \i48/i373  (.A(\i48/n16 ),
    .B(\i48/n35 ),
    .Y(\i48/n81 ));
 NAND2xp5_ASAP7_75t_SL \i48/i374  (.A(\i48/n5 ),
    .B(\i48/n46 ),
    .Y(\i48/n80 ));
 NAND2xp5_ASAP7_75t_SL \i48/i375  (.A(\i48/n548 ),
    .B(\i48/n46 ),
    .Y(\i48/n79 ));
 NOR2xp33_ASAP7_75t_SL \i48/i376  (.A(\i48/n45 ),
    .B(\i48/n535 ),
    .Y(\i48/n78 ));
 AND2x2_ASAP7_75t_SL \i48/i377  (.A(\i48/n5 ),
    .B(\i48/n61 ),
    .Y(\i48/n113 ));
 NAND2xp5_ASAP7_75t_SL \i48/i378  (.A(\i48/n546 ),
    .B(\i48/n457 ),
    .Y(\i48/n111 ));
 NOR2x1_ASAP7_75t_SL \i48/i379  (.A(\i48/n55 ),
    .B(\i48/n65 ),
    .Y(\i48/n109 ));
 NAND2xp5_ASAP7_75t_L \i48/i38  (.A(\i48/n576 ),
    .B(\i48/n414 ),
    .Y(\i48/n423 ));
 NAND2xp5_ASAP7_75t_SL \i48/i380  (.A(\i48/n5 ),
    .B(\i48/n560 ),
    .Y(\i48/n108 ));
 NAND2xp5_ASAP7_75t_SL \i48/i381  (.A(\i48/n549 ),
    .B(\i48/n470 ),
    .Y(\i48/n107 ));
 NAND2xp5_ASAP7_75t_SL \i48/i382  (.A(\i48/n37 ),
    .B(\i48/n59 ),
    .Y(\i48/n77 ));
 NAND2xp5_ASAP7_75t_SL \i48/i383  (.A(\i48/n43 ),
    .B(\i48/n46 ),
    .Y(\i48/n106 ));
 AND2x2_ASAP7_75t_SL \i48/i384  (.A(\i48/n5 ),
    .B(\i48/n41 ),
    .Y(\i48/n105 ));
 NOR2xp33_ASAP7_75t_SL \i48/i385  (.A(\i48/n55 ),
    .B(\i48/n46 ),
    .Y(\i48/n76 ));
 NAND2xp5_ASAP7_75t_SL \i48/i386  (.A(\i48/n548 ),
    .B(\i48/n559 ),
    .Y(\i48/n103 ));
 NAND2xp5_ASAP7_75t_SL \i48/i387  (.A(\i48/n548 ),
    .B(\i48/n41 ),
    .Y(\i48/n101 ));
 NAND2xp5_ASAP7_75t_SL \i48/i388  (.A(\i48/n37 ),
    .B(\i48/n41 ),
    .Y(\i48/n98 ));
 NAND2xp33_ASAP7_75t_L \i48/i389  (.A(\i48/n40 ),
    .B(\i48/n58 ),
    .Y(\i48/n75 ));
 NAND2xp33_ASAP7_75t_SL \i48/i39  (.A(\i48/n378 ),
    .B(\i48/n396 ),
    .Y(\i48/n422 ));
 NOR2xp67_ASAP7_75t_L \i48/i390  (.A(\i48/n35 ),
    .B(\i48/n535 ),
    .Y(\i48/n95 ));
 NAND2xp5_ASAP7_75t_SL \i48/i391  (.A(\i48/n39 ),
    .B(\i48/n560 ),
    .Y(\i48/n17 ));
 NAND2xp5_ASAP7_75t_SL \i48/i392  (.A(\i48/n39 ),
    .B(\i48/n65 ),
    .Y(\i48/n94 ));
 NAND2xp5_ASAP7_75t_L \i48/i393  (.A(\i48/n44 ),
    .B(\i48/n16 ),
    .Y(\i48/n93 ));
 NOR2xp67_ASAP7_75t_SL \i48/i394  (.A(\i48/n59 ),
    .B(\i48/n511 ),
    .Y(\i48/n92 ));
 NAND2xp5_ASAP7_75t_SL \i48/i395  (.A(\i48/n5 ),
    .B(\i48/n65 ),
    .Y(\i48/n74 ));
 NAND2xp5_ASAP7_75t_SL \i48/i396  (.A(\i48/n549 ),
    .B(\i48/n65 ),
    .Y(\i48/n90 ));
 NOR2xp33_ASAP7_75t_SL \i48/i397  (.A(\i48/n498 ),
    .B(\i48/n44 ),
    .Y(\i48/n73 ));
 NOR2xp33_ASAP7_75t_SL \i48/i398  (.A(\i48/n498 ),
    .B(\i48/n45 ),
    .Y(\i48/n72 ));
 INVx1_ASAP7_75t_SL \i48/i399  (.A(\i48/n71 ),
    .Y(\i48/n70 ));
 INVx2_ASAP7_75t_SL \i48/i4  (.A(\i48/n564 ),
    .Y(\i48/n4 ));
 NOR2x1_ASAP7_75t_SL \i48/i40  (.A(\i48/n452 ),
    .B(\i48/n404 ),
    .Y(\i48/n428 ));
 INVx3_ASAP7_75t_SL \i48/i400  (.A(\i48/n69 ),
    .Y(\i48/n68 ));
 INVx2_ASAP7_75t_SL \i48/i401  (.A(\i48/n559 ),
    .Y(\i48/n67 ));
 INVx3_ASAP7_75t_SL \i48/i402  (.A(\i48/n546 ),
    .Y(\i48/n66 ));
 INVx2_ASAP7_75t_SL \i48/i403  (.A(\i48/n548 ),
    .Y(\i48/n64 ));
 INVx4_ASAP7_75t_SL \i48/i404  (.A(\i48/n560 ),
    .Y(\i48/n63 ));
 INVx2_ASAP7_75t_SL \i48/i405  (.A(\i48/n549 ),
    .Y(\i48/n62 ));
 INVx3_ASAP7_75t_SL \i48/i406  (.A(\i48/n61 ),
    .Y(\i48/n60 ));
 INVx2_ASAP7_75t_SL \i48/i407  (.A(\i48/n59 ),
    .Y(\i48/n58 ));
 INVx2_ASAP7_75t_SL \i48/i408  (.A(\i48/n57 ),
    .Y(\i48/n56 ));
 INVx4_ASAP7_75t_SL \i48/i409  (.A(\i48/n55 ),
    .Y(\i48/n54 ));
 NAND2xp33_ASAP7_75t_L \i48/i41  (.A(\i48/n384 ),
    .B(\i48/n356 ),
    .Y(\i48/n419 ));
 INVx3_ASAP7_75t_SL \i48/i410  (.A(\i48/n53 ),
    .Y(\i48/n52 ));
 INVx3_ASAP7_75t_SL \i48/i411  (.A(\i48/n51 ),
    .Y(\i48/n50 ));
 AND2x4_ASAP7_75t_SL \i48/i412  (.A(\i48/n521 ),
    .B(\i48/n493 ),
    .Y(\i48/n71 ));
 OR2x4_ASAP7_75t_SL \i48/i413  (.A(\i48/n26 ),
    .B(\i48/n6 ),
    .Y(\i48/n69 ));
 AND2x4_ASAP7_75t_SL \i48/i414  (.A(\i48/n28 ),
    .B(\i48/n29 ),
    .Y(\i48/n65 ));
 NAND2x1_ASAP7_75t_SL \i48/i415  (.A(\i48/n28 ),
    .B(\i48/n29 ),
    .Y(\i48/n16 ));
 AND2x4_ASAP7_75t_SL \i48/i416  (.A(\i48/n28 ),
    .B(\i48/n468 ),
    .Y(\i48/n61 ));
 AND2x4_ASAP7_75t_SL \i48/i417  (.A(\i48/n454 ),
    .B(\i48/n14 ),
    .Y(\i48/n59 ));
 AND2x4_ASAP7_75t_SL \i48/i418  (.A(\i48/n454 ),
    .B(\i48/n28 ),
    .Y(\i48/n57 ));
 AND2x4_ASAP7_75t_SL \i48/i419  (.A(\i48/n28 ),
    .B(\i48/n27 ),
    .Y(\i48/n55 ));
 NAND2xp33_ASAP7_75t_L \i48/i42  (.A(\i48/n576 ),
    .B(\i48/n361 ),
    .Y(\i48/n418 ));
 AND2x4_ASAP7_75t_SL \i48/i420  (.A(\i48/n521 ),
    .B(\i48/n482 ),
    .Y(\i48/n53 ));
 OR2x6_ASAP7_75t_SL \i48/i421  (.A(\i48/n31 ),
    .B(\i48/n545 ),
    .Y(\i48/n51 ));
 INVx2_ASAP7_75t_SL \i48/i422  (.A(\i48/n49 ),
    .Y(\i48/n15 ));
 INVx3_ASAP7_75t_SL \i48/i423  (.A(\i48/n48 ),
    .Y(\i48/n47 ));
 INVx2_ASAP7_75t_SL \i48/i424  (.A(\i48/n46 ),
    .Y(\i48/n45 ));
 INVx4_ASAP7_75t_SL \i48/i425  (.A(\i48/n470 ),
    .Y(\i48/n44 ));
 INVx4_ASAP7_75t_SL \i48/i426  (.A(\i48/n43 ),
    .Y(\i48/n42 ));
 INVx3_ASAP7_75t_SL \i48/i427  (.A(\i48/n39 ),
    .Y(\i48/n38 ));
 INVx4_ASAP7_75t_SL \i48/i428  (.A(\i48/n37 ),
    .Y(\i48/n36 ));
 INVx11_ASAP7_75t_SL \i48/i429  (.A(\i48/n35 ),
    .Y(\i48/n34 ));
 NOR2xp33_ASAP7_75t_SL \i48/i43  (.A(\i48/n360 ),
    .B(\i48/n386 ),
    .Y(\i48/n417 ));
 AND2x4_ASAP7_75t_SL \i48/i430  (.A(\i48/n493 ),
    .B(\i48/n33 ),
    .Y(\i48/n49 ));
 AND2x4_ASAP7_75t_SL \i48/i431  (.A(\i48/n531 ),
    .B(\i48/n493 ),
    .Y(\i48/n48 ));
 AND2x4_ASAP7_75t_SL \i48/i432  (.A(\i48/n468 ),
    .B(\i48/n14 ),
    .Y(\i48/n46 ));
 AND2x4_ASAP7_75t_SL \i48/i433  (.A(\i48/n32 ),
    .B(\i48/n532 ),
    .Y(\i48/n43 ));
 AND2x4_ASAP7_75t_SL \i48/i434  (.A(\i48/n3 ),
    .B(\i48/n29 ),
    .Y(\i48/n41 ));
 NAND2x1_ASAP7_75t_SL \i48/i435  (.A(\i48/n3 ),
    .B(\i48/n29 ),
    .Y(\i48/n40 ));
 AND2x4_ASAP7_75t_SL \i48/i436  (.A(\i48/n482 ),
    .B(\i48/n531 ),
    .Y(\i48/n39 ));
 AND2x4_ASAP7_75t_SL \i48/i437  (.A(\i48/n33 ),
    .B(\i48/n482 ),
    .Y(\i48/n37 ));
 OR2x6_ASAP7_75t_SL \i48/i438  (.A(\i48/n25 ),
    .B(\i48/n30 ),
    .Y(\i48/n35 ));
 INVx2_ASAP7_75t_SL \i48/i439  (.A(\i48/n550 ),
    .Y(\i48/n33 ));
 NAND3xp33_ASAP7_75t_SL \i48/i44  (.A(\i48/n351 ),
    .B(\i48/n358 ),
    .C(\i48/n326 ),
    .Y(\i48/n416 ));
 NAND2xp5_ASAP7_75t_SL \i48/i440  (.A(\i48/n9 ),
    .B(\i48/n2 ),
    .Y(\i48/n30 ));
 NAND2x1p5_ASAP7_75t_SL \i48/i441  (.A(n25[4]),
    .B(n25[5]),
    .Y(\i48/n31 ));
 INVx2_ASAP7_75t_SL \i48/i442  (.A(\i48/n6 ),
    .Y(\i48/n29 ));
 INVx2_ASAP7_75t_SL \i48/i443  (.A(\i48/n507 ),
    .Y(\i48/n27 ));
 NAND2xp5_ASAP7_75t_SL \i48/i444  (.A(\i48/n24 ),
    .B(\i48/n10 ),
    .Y(\i48/n25 ));
 AND2x4_ASAP7_75t_SL \i48/i445  (.A(n25[2]),
    .B(n25[3]),
    .Y(\i48/n28 ));
 NAND2x1_ASAP7_75t_SL \i48/i446  (.A(n25[3]),
    .B(\i48/n2 ),
    .Y(\i48/n26 ));
 INVx1_ASAP7_75t_SL \i48/i447  (.A(n25[1]),
    .Y(\i48/n24 ));
 INVx2_ASAP7_75t_SL \i48/i448  (.A(\i48/n26 ),
    .Y(\i48/n14 ));
 INVx2_ASAP7_75t_SL \i48/i449  (.A(n25[6]),
    .Y(\i48/n13 ));
 NOR2x1_ASAP7_75t_SL \i48/i45  (.A(\i48/n308 ),
    .B(\i48/n369 ),
    .Y(\i48/n415 ));
 INVx2_ASAP7_75t_SL \i48/i450  (.A(n25[7]),
    .Y(\i48/n11 ));
 INVx3_ASAP7_75t_SL \i48/i451  (.A(n25[0]),
    .Y(\i48/n10 ));
 INVx2_ASAP7_75t_SL \i48/i452  (.A(n25[3]),
    .Y(\i48/n9 ));
 INVx1_ASAP7_75t_SL \i48/i453  (.A(\i48/n381 ),
    .Y(\i48/n8 ));
 OR2x2_ASAP7_75t_SL \i48/i454  (.A(\i48/n105 ),
    .B(\i48/n517 ),
    .Y(\i48/n7 ));
 OR2x2_ASAP7_75t_SL \i48/i455  (.A(n25[0]),
    .B(n25[1]),
    .Y(\i48/n6 ));
 NAND4xp25_ASAP7_75t_SL \i48/i456  (.A(\i48/n354 ),
    .B(\i48/n449 ),
    .C(\i48/n348 ),
    .D(\i48/n380 ),
    .Y(\i48/n450 ));
 NOR2xp67_ASAP7_75t_SL \i48/i457  (.A(\i48/n477 ),
    .B(\i48/n509 ),
    .Y(\i48/n449 ));
 NAND3xp33_ASAP7_75t_L \i48/i458  (.A(\i48/n331 ),
    .B(\i48/n449 ),
    .C(\i48/n398 ),
    .Y(\i48/n451 ));
 NAND4xp25_ASAP7_75t_SL \i48/i459  (.A(\i48/n341 ),
    .B(\i48/n449 ),
    .C(\i48/n353 ),
    .D(\i48/n337 ),
    .Y(\i48/n452 ));
 NOR2xp33_ASAP7_75t_SL \i48/i46  (.A(\i48/n376 ),
    .B(\i48/n289 ),
    .Y(\i48/n414 ));
 OAI221xp5_ASAP7_75t_SL \i48/i460  (.A1(\i48/n467 ),
    .A2(\i48/n62 ),
    .B1(\i48/n54 ),
    .B2(\i48/n52 ),
    .C(\i48/n182 ),
    .Y(\i48/n453 ));
 AND2x2_ASAP7_75t_SL \i48/i461  (.A(n25[0]),
    .B(n25[1]),
    .Y(\i48/n454 ));
 AND2x2_ASAP7_75t_SL \i48/i462  (.A(\i48/n9 ),
    .B(\i48/n2 ),
    .Y(\i48/n455 ));
 INVx4_ASAP7_75t_SL \i48/i463  (.A(\i48/n456 ),
    .Y(\i48/n457 ));
 NAND2x1p5_ASAP7_75t_SL \i48/i464  (.A(\i48/n454 ),
    .B(\i48/n455 ),
    .Y(\i48/n456 ));
 OAI22xp5_ASAP7_75t_SL \i48/i465  (.A1(\i48/n42 ),
    .A2(\i48/n456 ),
    .B1(\i48/n51 ),
    .B2(\i48/n58 ),
    .Y(\i48/n458 ));
 OAI221xp5_ASAP7_75t_SL \i48/i466  (.A1(\i48/n491 ),
    .A2(\i48/n69 ),
    .B1(\i48/n456 ),
    .B2(\i48/n52 ),
    .C(\i48/n142 ),
    .Y(\i48/n459 ));
 NOR2xp33_ASAP7_75t_SL \i48/i467  (.A(\i48/n456 ),
    .B(\i48/n36 ),
    .Y(\i48/n460 ));
 NAND2xp5_ASAP7_75t_SL \i48/i468  (.A(\i48/n37 ),
    .B(\i48/n4 ),
    .Y(\i48/n461 ));
 NOR2xp67_ASAP7_75t_SL \i48/i469  (.A(\i48/n467 ),
    .B(\i48/n42 ),
    .Y(\i48/n462 ));
 NAND2xp5_ASAP7_75t_SL \i48/i47  (.A(\i48/n384 ),
    .B(\i48/n379 ),
    .Y(\i48/n413 ));
 OAI22xp5_ASAP7_75t_SL \i48/i470  (.A1(\i48/n70 ),
    .A2(\i48/n564 ),
    .B1(\i48/n552 ),
    .B2(\i48/n467 ),
    .Y(\i48/n463 ));
 OAI22xp33_ASAP7_75t_SL \i48/i471  (.A1(\i48/n47 ),
    .A2(\i48/n35 ),
    .B1(\i48/n467 ),
    .B2(\i48/n484 ),
    .Y(\i48/n464 ));
 OAI22xp5_ASAP7_75t_SL \i48/i472  (.A1(\i48/n47 ),
    .A2(\i48/n467 ),
    .B1(\i48/n498 ),
    .B2(\i48/n44 ),
    .Y(\i48/n465 ));
 OAI221xp5_ASAP7_75t_SL \i48/i473  (.A1(\i48/n467 ),
    .A2(\i48/n64 ),
    .B1(\i48/n16 ),
    .B2(\i48/n15 ),
    .C(\i48/n216 ),
    .Y(\i48/n466 ));
 AND2x4_ASAP7_75t_SL \i48/i474  (.A(n25[0]),
    .B(\i48/n24 ),
    .Y(\i48/n468 ));
 NAND2xp33_ASAP7_75t_SL \i48/i475  (.A(\i48/n456 ),
    .B(\i48/n564 ),
    .Y(\i48/n469 ));
 NAND2xp5_ASAP7_75t_SL \i48/i476  (.A(\i48/n71 ),
    .B(\i48/n470 ),
    .Y(\i48/n471 ));
 OAI21xp5_ASAP7_75t_SL \i48/i477  (.A1(\i48/n59 ),
    .A2(\i48/n470 ),
    .B(\i48/n50 ),
    .Y(\i48/n472 ));
 OAI21xp5_ASAP7_75t_SL \i48/i478  (.A1(\i48/n511 ),
    .A2(\i48/n470 ),
    .B(\i48/n546 ),
    .Y(\i48/n473 ));
 AOI21x1_ASAP7_75t_SL \i48/i479  (.A1(\i48/n470 ),
    .A2(\i48/n48 ),
    .B(\i48/n465 ),
    .Y(\i48/n474 ));
 NOR2x1_ASAP7_75t_SL \i48/i48  (.A(\i48/n293 ),
    .B(\i48/n386 ),
    .Y(\i48/n412 ));
 INVx2_ASAP7_75t_L \i48/i480  (.A(\i48/n468 ),
    .Y(\i48/n475 ));
 INVx2_ASAP7_75t_SL \i48/i481  (.A(\i48/n455 ),
    .Y(\i48/n476 ));
 OAI22xp5_ASAP7_75t_SL \i48/i482  (.A1(\i48/n524 ),
    .A2(\i48/n63 ),
    .B1(\i48/n52 ),
    .B2(\i48/n467 ),
    .Y(\i48/n477 ));
 INVx4_ASAP7_75t_SL \i48/i483  (.A(\i48/n467 ),
    .Y(\i48/n478 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i48/i484  (.A1(\i48/n467 ),
    .A2(\i48/n40 ),
    .B(\i48/n52 ),
    .C(\i48/n94 ),
    .Y(\i48/n479 ));
 AOI21xp5_ASAP7_75t_L \i48/i485  (.A1(\i48/n484 ),
    .A2(\i48/n145 ),
    .B(\i48/n467 ),
    .Y(\i48/n480 ));
 OAI222xp33_ASAP7_75t_SL \i48/i486  (.A1(\i48/n467 ),
    .A2(\i48/n36 ),
    .B1(\i48/n40 ),
    .B2(\i48/n15 ),
    .C1(\i48/n56 ),
    .C2(\i48/n51 ),
    .Y(\i48/n481 ));
 AND2x2_ASAP7_75t_SL \i48/i487  (.A(n25[7]),
    .B(\i48/n13 ),
    .Y(\i48/n482 ));
 INVx3_ASAP7_75t_SL \i48/i488  (.A(\i48/n483 ),
    .Y(\i48/n484 ));
 AND2x4_ASAP7_75t_SL \i48/i489  (.A(\i48/n32 ),
    .B(\i48/n482 ),
    .Y(\i48/n483 ));
 NOR2x1_ASAP7_75t_SL \i48/i49  (.A(\i48/n359 ),
    .B(\i48/n370 ),
    .Y(\i48/n411 ));
 OAI31xp33_ASAP7_75t_SL \i48/i490  (.A1(\i48/n457 ),
    .A2(\i48/n511 ),
    .A3(\i48/n68 ),
    .B(\i48/n483 ),
    .Y(\i48/n485 ));
 AOI21xp5_ASAP7_75t_SL \i48/i491  (.A1(\i48/n59 ),
    .A2(\i48/n483 ),
    .B(\i48/n223 ),
    .Y(\i48/n486 ));
 NAND2xp5_ASAP7_75t_SL \i48/i492  (.A(\i48/n483 ),
    .B(\i48/n55 ),
    .Y(\i48/n487 ));
 NAND2xp5_ASAP7_75t_SL \i48/i493  (.A(\i48/n483 ),
    .B(\i48/n46 ),
    .Y(\i48/n488 ));
 NOR2xp33_ASAP7_75t_SL \i48/i494  (.A(\i48/n483 ),
    .B(\i48/n546 ),
    .Y(\i48/n489 ));
 NAND2xp5_ASAP7_75t_SL \i48/i495  (.A(\i48/n483 ),
    .B(\i48/n560 ),
    .Y(\i48/n490 ));
 NOR2x1_ASAP7_75t_SL \i48/i496  (.A(\i48/n483 ),
    .B(\i48/n548 ),
    .Y(\i48/n491 ));
 OAI221xp5_ASAP7_75t_SL \i48/i497  (.A1(\i48/n70 ),
    .A2(\i48/n92 ),
    .B1(\i48/n92 ),
    .B2(\i48/n552 ),
    .C(\i48/n525 ),
    .Y(\i48/n492 ));
 AND2x2_ASAP7_75t_SL \i48/i498  (.A(\i48/n11 ),
    .B(\i48/n13 ),
    .Y(\i48/n493 ));
 INVx3_ASAP7_75t_SL \i48/i499  (.A(\i48/n31 ),
    .Y(\i48/n32 ));
 INVx3_ASAP7_75t_SL \i48/i5  (.A(\i48/n552 ),
    .Y(\i48/n5 ));
 NAND2xp5_ASAP7_75t_SL \i48/i50  (.A(\i48/n325 ),
    .B(\i48/n364 ),
    .Y(\i48/n410 ));
 AOI22xp5_ASAP7_75t_SL \i48/i500  (.A1(\i48/n494 ),
    .A2(\i48/n41 ),
    .B1(\i48/n483 ),
    .B2(\i48/n57 ),
    .Y(\i48/n495 ));
 AND2x4_ASAP7_75t_SL \i48/i501  (.A(\i48/n493 ),
    .B(\i48/n32 ),
    .Y(\i48/n494 ));
 AOI22xp5_ASAP7_75t_SL \i48/i502  (.A1(\i48/n494 ),
    .A2(\i48/n478 ),
    .B1(\i48/n546 ),
    .B2(\i48/n470 ),
    .Y(\i48/n496 ));
 AOI22xp5_ASAP7_75t_SL \i48/i503  (.A1(\i48/n559 ),
    .A2(\i48/n494 ),
    .B1(\i48/n548 ),
    .B2(\i48/n57 ),
    .Y(\i48/n497 ));
 INVx2_ASAP7_75t_SL \i48/i504  (.A(\i48/n494 ),
    .Y(\i48/n498 ));
 AOI22xp5_ASAP7_75t_SL \i48/i505  (.A1(\i48/n34 ),
    .A2(\i48/n37 ),
    .B1(\i48/n494 ),
    .B2(\i48/n59 ),
    .Y(\i48/n499 ));
 AND2x2_ASAP7_75t_SL \i48/i506  (.A(\i48/n494 ),
    .B(\i48/n57 ),
    .Y(\i48/n500 ));
 NAND2xp5_ASAP7_75t_SL \i48/i507  (.A(\i48/n494 ),
    .B(\i48/n511 ),
    .Y(\i48/n501 ));
 NAND2xp5_ASAP7_75t_SL \i48/i508  (.A(\i48/n34 ),
    .B(\i48/n494 ),
    .Y(\i48/n502 ));
 AND2x2_ASAP7_75t_SL \i48/i509  (.A(\i48/n494 ),
    .B(\i48/n65 ),
    .Y(\i48/n503 ));
 NOR5xp2_ASAP7_75t_SL \i48/i51  (.A(\i48/n254 ),
    .B(\i48/n512 ),
    .C(\i48/n265 ),
    .D(\i48/n22 ),
    .E(\i48/n453 ),
    .Y(\i48/n409 ));
 AND2x2_ASAP7_75t_SL \i48/i510  (.A(\i48/n494 ),
    .B(\i48/n457 ),
    .Y(\i48/n504 ));
 NAND2xp5_ASAP7_75t_SL \i48/i511  (.A(\i48/n494 ),
    .B(\i48/n61 ),
    .Y(\i48/n505 ));
 OR2x2_ASAP7_75t_SL \i48/i512  (.A(\i48/n2 ),
    .B(n25[3]),
    .Y(\i48/n506 ));
 NAND2x1_ASAP7_75t_SL \i48/i513  (.A(\i48/n10 ),
    .B(n25[1]),
    .Y(\i48/n507 ));
 OAI221xp5_ASAP7_75t_SL \i48/i514  (.A1(\i48/n535 ),
    .A2(\i48/n40 ),
    .B1(\i48/n508 ),
    .B2(\i48/n36 ),
    .C(\i48/n502 ),
    .Y(\i48/n509 ));
 OR2x4_ASAP7_75t_SL \i48/i515  (.A(\i48/n506 ),
    .B(\i48/n507 ),
    .Y(\i48/n508 ));
 OAI21xp5_ASAP7_75t_SL \i48/i516  (.A1(\i48/n62 ),
    .A2(\i48/n508 ),
    .B(\i48/n106 ),
    .Y(\i48/n510 ));
 INVx4_ASAP7_75t_SL \i48/i517  (.A(\i48/n508 ),
    .Y(\i48/n511 ));
 OAI221xp5_ASAP7_75t_SL \i48/i518  (.A1(\i48/n45 ),
    .A2(\i48/n524 ),
    .B1(\i48/n42 ),
    .B2(\i48/n508 ),
    .C(\i48/n540 ),
    .Y(\i48/n512 ));
 AO21x1_ASAP7_75t_SL \i48/i519  (.A1(\i48/n508 ),
    .A2(\i48/n134 ),
    .B(\i48/n489 ),
    .Y(\i48/n513 ));
 NOR2x1_ASAP7_75t_SL \i48/i52  (.A(\i48/n8 ),
    .B(\i48/n371 ),
    .Y(\i48/n408 ));
 AOI31xp33_ASAP7_75t_SL \i48/i520  (.A1(\i48/n42 ),
    .A2(\i48/n64 ),
    .A3(\i48/n52 ),
    .B(\i48/n508 ),
    .Y(\i48/n514 ));
 OAI22xp33_ASAP7_75t_SL \i48/i521  (.A1(\i48/n38 ),
    .A2(\i48/n69 ),
    .B1(\i48/n508 ),
    .B2(\i48/n47 ),
    .Y(\i48/n515 ));
 OA21x2_ASAP7_75t_SL \i48/i522  (.A1(\i48/n42 ),
    .A2(\i48/n508 ),
    .B(\i48/n540 ),
    .Y(\i48/n516 ));
 OAI22xp5_ASAP7_75t_SL \i48/i523  (.A1(\i48/n42 ),
    .A2(\i48/n63 ),
    .B1(\i48/n51 ),
    .B2(\i48/n508 ),
    .Y(\i48/n517 ));
 OAI22xp5_ASAP7_75t_SL \i48/i524  (.A1(\i48/n42 ),
    .A2(\i48/n40 ),
    .B1(\i48/n508 ),
    .B2(\i48/n38 ),
    .Y(\i48/n518 ));
 NOR2xp33_ASAP7_75t_SL \i48/i525  (.A(\i48/n508 ),
    .B(\i48/n524 ),
    .Y(\i48/n519 ));
 NOR2xp33_ASAP7_75t_SL \i48/i526  (.A(\i48/n508 ),
    .B(\i48/n38 ),
    .Y(\i48/n520 ));
 AND2x4_ASAP7_75t_SL \i48/i527  (.A(\i48/n0 ),
    .B(\i48/n1 ),
    .Y(\i48/n521 ));
 AOI22xp33_ASAP7_75t_SL \i48/i528  (.A1(\i48/n522 ),
    .A2(\i48/n457 ),
    .B1(\i48/n494 ),
    .B2(\i48/n46 ),
    .Y(\i48/n523 ));
 AND2x4_ASAP7_75t_SL \i48/i529  (.A(\i48/n521 ),
    .B(\i48/n532 ),
    .Y(\i48/n522 ));
 NAND2x1_ASAP7_75t_SL \i48/i53  (.A(\i48/n368 ),
    .B(\i48/n349 ),
    .Y(\i48/n421 ));
 INVx3_ASAP7_75t_SL \i48/i530  (.A(\i48/n522 ),
    .Y(\i48/n524 ));
 AOI211x1_ASAP7_75t_SL \i48/i531  (.A1(\i48/n81 ),
    .A2(\i48/n522 ),
    .B(\i48/n158 ),
    .C(\i48/n160 ),
    .Y(\i48/n525 ));
 AOI22xp5_ASAP7_75t_SL \i48/i532  (.A1(\i48/n522 ),
    .A2(\i48/n68 ),
    .B1(\i48/n5 ),
    .B2(\i48/n65 ),
    .Y(\i48/n526 ));
 NAND2xp5_ASAP7_75t_SL \i48/i533  (.A(\i48/n522 ),
    .B(\i48/n4 ),
    .Y(\i48/n527 ));
 NAND2xp5_ASAP7_75t_SL \i48/i534  (.A(\i48/n61 ),
    .B(\i48/n522 ),
    .Y(\i48/n528 ));
 NAND2xp5_ASAP7_75t_SL \i48/i535  (.A(\i48/n522 ),
    .B(\i48/n41 ),
    .Y(\i48/n529 ));
 OR2x2_ASAP7_75t_SL \i48/i536  (.A(\i48/n39 ),
    .B(\i48/n522 ),
    .Y(\i48/n530 ));
 AND2x2_ASAP7_75t_SL \i48/i537  (.A(\i48/n0 ),
    .B(n25[4]),
    .Y(\i48/n531 ));
 AND2x2_ASAP7_75t_L \i48/i538  (.A(\i48/n11 ),
    .B(n25[6]),
    .Y(\i48/n532 ));
 NAND2xp5_ASAP7_75t_SL \i48/i539  (.A(\i48/n533 ),
    .B(\i48/n470 ),
    .Y(\i48/n534 ));
 NOR2x1_ASAP7_75t_SL \i48/i54  (.A(\i48/n387 ),
    .B(\i48/n370 ),
    .Y(\i48/n407 ));
 AND2x4_ASAP7_75t_SL \i48/i540  (.A(\i48/n531 ),
    .B(\i48/n532 ),
    .Y(\i48/n533 ));
 INVx4_ASAP7_75t_SL \i48/i541  (.A(\i48/n533 ),
    .Y(\i48/n535 ));
 OAI21xp33_ASAP7_75t_SL \i48/i542  (.A1(\i48/n511 ),
    .A2(\i48/n41 ),
    .B(\i48/n533 ),
    .Y(\i48/n536 ));
 OAI21xp5_ASAP7_75t_SL \i48/i543  (.A1(\i48/n533 ),
    .A2(\i48/n53 ),
    .B(\i48/n55 ),
    .Y(\i48/n537 ));
 OAI21xp5_ASAP7_75t_SL \i48/i544  (.A1(\i48/n548 ),
    .A2(\i48/n533 ),
    .B(\i48/n511 ),
    .Y(\i48/n538 ));
 AOI22xp5_ASAP7_75t_SL \i48/i545  (.A1(\i48/n533 ),
    .A2(\i48/n65 ),
    .B1(\i48/n37 ),
    .B2(\i48/n457 ),
    .Y(\i48/n539 ));
 NAND2xp5_ASAP7_75t_SL \i48/i546  (.A(\i48/n533 ),
    .B(\i48/n59 ),
    .Y(\i48/n540 ));
 NAND2xp5_ASAP7_75t_SL \i48/i547  (.A(\i48/n533 ),
    .B(\i48/n61 ),
    .Y(\i48/n541 ));
 NAND2xp5_ASAP7_75t_SL \i48/i548  (.A(\i48/n533 ),
    .B(\i48/n560 ),
    .Y(\i48/n542 ));
 NAND2xp5_ASAP7_75t_SL \i48/i549  (.A(\i48/n533 ),
    .B(\i48/n478 ),
    .Y(\i48/n543 ));
 NOR2x1_ASAP7_75t_SL \i48/i55  (.A(\i48/n307 ),
    .B(\i48/n369 ),
    .Y(\i48/n420 ));
 INVx2_ASAP7_75t_SL \i48/i550  (.A(\i48/n544 ),
    .Y(\i48/n545 ));
 AND2x2_ASAP7_75t_SL \i48/i551  (.A(n25[7]),
    .B(n25[6]),
    .Y(\i48/n544 ));
 AND2x4_ASAP7_75t_SL \i48/i552  (.A(\i48/n544 ),
    .B(\i48/n33 ),
    .Y(\i48/n546 ));
 AOI211xp5_ASAP7_75t_R \i48/i553  (.A1(\i48/n68 ),
    .A2(\i48/n544 ),
    .B(\i48/n503 ),
    .C(\i48/n99 ),
    .Y(\i48/n547 ));
 AND2x4_ASAP7_75t_SL \i48/i554  (.A(\i48/n544 ),
    .B(\i48/n521 ),
    .Y(\i48/n548 ));
 AND2x4_ASAP7_75t_SL \i48/i555  (.A(\i48/n544 ),
    .B(\i48/n531 ),
    .Y(\i48/n549 ));
 NAND2xp5_ASAP7_75t_SL \i48/i556  (.A(\i48/n1 ),
    .B(n25[5]),
    .Y(\i48/n550 ));
 NAND2xp5_ASAP7_75t_SL \i48/i557  (.A(\i48/n51 ),
    .B(\i48/n552 ),
    .Y(\i48/n553 ));
 OR2x2_ASAP7_75t_SL \i48/i558  (.A(\i48/n551 ),
    .B(\i48/n550 ),
    .Y(\i48/n552 ));
 NAND2xp5_ASAP7_75t_SL \i48/i559  (.A(\i48/n11 ),
    .B(n25[6]),
    .Y(\i48/n551 ));
 INVxp67_ASAP7_75t_SL \i48/i56  (.A(\i48/n405 ),
    .Y(\i48/n406 ));
 OAI21xp5_ASAP7_75t_SL \i48/i560  (.A1(\i48/n552 ),
    .A2(\i48/n564 ),
    .B(\i48/n98 ),
    .Y(\i48/n554 ));
 AND2x4_ASAP7_75t_SL \i48/i561  (.A(\i48/n27 ),
    .B(\i48/n14 ),
    .Y(\i48/n470 ));
 NAND4xp25_ASAP7_75t_SL \i48/i562  (.A(\i48/n178 ),
    .B(\i48/n191 ),
    .C(\i48/n277 ),
    .D(\i48/n555 ),
    .Y(\i48/n556 ));
 NAND2x1p5_ASAP7_75t_SL \i48/i563  (.A(\i48/n5 ),
    .B(\i48/n470 ),
    .Y(\i48/n555 ));
 INVx1_ASAP7_75t_SL \i48/i564  (.A(\i48/n555 ),
    .Y(\i48/n557 ));
 NAND2xp5_ASAP7_75t_L \i48/i565  (.A(\i48/n555 ),
    .B(\i48/n132 ),
    .Y(\i48/n558 ));
 AND2x4_ASAP7_75t_SL \i48/i566  (.A(\i48/n454 ),
    .B(\i48/n3 ),
    .Y(\i48/n559 ));
 AND2x4_ASAP7_75t_SL \i48/i567  (.A(\i48/n455 ),
    .B(\i48/n27 ),
    .Y(\i48/n560 ));
 OA21x2_ASAP7_75t_SL \i48/i568  (.A1(\i48/n36 ),
    .A2(\i48/n561 ),
    .B(\i48/n101 ),
    .Y(\i48/n562 ));
 NOR2xp33_ASAP7_75t_SL \i48/i569  (.A(\i48/n559 ),
    .B(\i48/n560 ),
    .Y(\i48/n561 ));
 INVxp67_ASAP7_75t_SL \i48/i57  (.A(\i48/n401 ),
    .Y(\i48/n402 ));
 OAI21xp33_ASAP7_75t_SL \i48/i570  (.A1(\i48/n42 ),
    .A2(\i48/n561 ),
    .B(\i48/n161 ),
    .Y(\i48/n563 ));
 NAND2x1p5_ASAP7_75t_SL \i48/i571  (.A(\i48/n3 ),
    .B(\i48/n468 ),
    .Y(\i48/n564 ));
 NAND2xp5_ASAP7_75t_SL \i48/i572  (.A(\i48/n4 ),
    .B(\i48/n533 ),
    .Y(\i48/n565 ));
 AOI22xp33_ASAP7_75t_SL \i48/i573  (.A1(\i48/n71 ),
    .A2(\i48/n511 ),
    .B1(\i48/n522 ),
    .B2(\i48/n4 ),
    .Y(\i48/n566 ));
 NAND2xp5_ASAP7_75t_SL \i48/i574  (.A(\i48/n494 ),
    .B(\i48/n4 ),
    .Y(\i48/n567 ));
 AOI22xp5_ASAP7_75t_SL \i48/i575  (.A1(\i48/n494 ),
    .A2(\i48/n560 ),
    .B1(\i48/n549 ),
    .B2(\i48/n4 ),
    .Y(\i48/n568 ));
 NAND2xp33_ASAP7_75t_L \i48/i576  (.A(\i48/n4 ),
    .B(\i48/n549 ),
    .Y(\i48/n569 ));
 AO21x2_ASAP7_75t_SL \i48/i577  (.A1(\i48/n548 ),
    .A2(\i48/n4 ),
    .B(\i48/n177 ),
    .Y(\i48/n570 ));
 NAND2xp5_ASAP7_75t_SL \i48/i578  (.A(\i48/n546 ),
    .B(\i48/n4 ),
    .Y(\i48/n571 ));
 NOR2xp33_ASAP7_75t_SL \i48/i579  (.A(\i48/n559 ),
    .B(\i48/n4 ),
    .Y(\i48/n572 ));
 AND5x1_ASAP7_75t_SL \i48/i58  (.A(\i48/n321 ),
    .B(\i48/n302 ),
    .C(\i48/n313 ),
    .D(\i48/n242 ),
    .E(\i48/n222 ),
    .Y(\i48/n400 ));
 AOI22xp5_ASAP7_75t_SL \i48/i580  (.A1(\i48/n548 ),
    .A2(\i48/n457 ),
    .B1(\i48/n39 ),
    .B2(\i48/n4 ),
    .Y(\i48/n573 ));
 OAI31xp33_ASAP7_75t_SL \i48/i581  (.A1(\i48/n57 ),
    .A2(\i48/n4 ),
    .A3(\i48/n470 ),
    .B(\i48/n39 ),
    .Y(\i48/n574 ));
 OR2x6_ASAP7_75t_SL \i48/i582  (.A(\i48/n475 ),
    .B(\i48/n476 ),
    .Y(\i48/n467 ));
 AND4x1_ASAP7_75t_SL \i48/i583  (.A(\i48/n253 ),
    .B(\i48/n291 ),
    .C(\i48/n302 ),
    .D(\i48/n231 ),
    .Y(\i48/n575 ));
 AND4x1_ASAP7_75t_SL \i48/i584  (.A(\i48/n243 ),
    .B(\i48/n486 ),
    .C(\i48/n264 ),
    .D(\i48/n253 ),
    .Y(\i48/n576 ));
 AO221x1_ASAP7_75t_SL \i48/i585  (.A1(\i48/n522 ),
    .A2(\i48/n59 ),
    .B1(\i48/n5 ),
    .B2(\i48/n511 ),
    .C(\i48/n229 ),
    .Y(\i48/n577 ));
 NAND3xp33_ASAP7_75t_SL \i48/i586  (.A(\i48/n578 ),
    .B(\i48/n526 ),
    .C(\i48/n283 ),
    .Y(\i48/n579 ));
 AO21x1_ASAP7_75t_SL \i48/i587  (.A1(\i48/n524 ),
    .A2(\i48/n42 ),
    .B(\i48/n67 ),
    .Y(\i48/n578 ));
 NOR3xp33_ASAP7_75t_SL \i48/i588  (.A(\i48/n580 ),
    .B(\i48/n563 ),
    .C(\i48/n177 ),
    .Y(\i48/n581 ));
 OAI21xp5_ASAP7_75t_SL \i48/i589  (.A1(\i48/n51 ),
    .A2(\i48/n16 ),
    .B(\i48/n565 ),
    .Y(\i48/n580 ));
 NOR3xp33_ASAP7_75t_SL \i48/i59  (.A(\i48/n332 ),
    .B(\i48/n312 ),
    .C(\i48/n294 ),
    .Y(\i48/n399 ));
 NOR2x2_ASAP7_75t_SL \i48/i6  (.A(\i48/n444 ),
    .B(\i48/n443 ),
    .Y(n24[4]));
 NOR3xp33_ASAP7_75t_SL \i48/i60  (.A(\i48/n556 ),
    .B(\i48/n295 ),
    .C(\i48/n252 ),
    .Y(\i48/n398 ));
 AND5x1_ASAP7_75t_SL \i48/i61  (.A(\i48/n285 ),
    .B(\i48/n298 ),
    .C(\i48/n547 ),
    .D(\i48/n288 ),
    .E(\i48/n228 ),
    .Y(\i48/n397 ));
 NOR2xp33_ASAP7_75t_SL \i48/i62  (.A(\i48/n357 ),
    .B(\i48/n362 ),
    .Y(\i48/n396 ));
 NAND5xp2_ASAP7_75t_SL \i48/i63  (.A(\i48/n320 ),
    .B(\i48/n279 ),
    .C(\i48/n194 ),
    .D(\i48/n180 ),
    .E(\i48/n12 ),
    .Y(\i48/n395 ));
 NOR4xp25_ASAP7_75t_SL \i48/i64  (.A(\i48/n310 ),
    .B(\i48/n512 ),
    .C(\i48/n266 ),
    .D(\i48/n245 ),
    .Y(\i48/n394 ));
 NAND4xp25_ASAP7_75t_SL \i48/i65  (.A(\i48/n329 ),
    .B(\i48/n346 ),
    .C(\i48/n343 ),
    .D(\i48/n348 ),
    .Y(\i48/n393 ));
 NAND4xp25_ASAP7_75t_SL \i48/i66  (.A(\i48/n355 ),
    .B(\i48/n353 ),
    .C(\i48/n516 ),
    .D(\i48/n221 ),
    .Y(\i48/n392 ));
 NOR2x1_ASAP7_75t_SL \i48/i67  (.A(\i48/n173 ),
    .B(\i48/n383 ),
    .Y(\i48/n391 ));
 NAND3xp33_ASAP7_75t_SL \i48/i68  (.A(\i48/n348 ),
    .B(\i48/n319 ),
    .C(\i48/n17 ),
    .Y(\i48/n405 ));
 NAND4xp75_ASAP7_75t_SL \i48/i69  (.A(\i48/n525 ),
    .B(\i48/n234 ),
    .C(\i48/n306 ),
    .D(\i48/n19 ),
    .Y(\i48/n404 ));
 NOR2x1p5_ASAP7_75t_SL \i48/i7  (.A(\i48/n439 ),
    .B(\i48/n445 ),
    .Y(n24[3]));
 NAND2xp33_ASAP7_75t_SL \i48/i70  (.A(\i48/n328 ),
    .B(\i48/n388 ),
    .Y(\i48/n390 ));
 AND2x2_ASAP7_75t_SL \i48/i71  (.A(\i48/n331 ),
    .B(\i48/n377 ),
    .Y(\i48/n403 ));
 NAND2x1p5_ASAP7_75t_SL \i48/i72  (.A(\i48/n385 ),
    .B(\i48/n342 ),
    .Y(\i48/n401 ));
 INVxp67_ASAP7_75t_SL \i48/i73  (.A(\i48/n388 ),
    .Y(\i48/n389 ));
 INVxp67_ASAP7_75t_SL \i48/i74  (.A(\i48/n382 ),
    .Y(\i48/n383 ));
 NOR5xp2_ASAP7_75t_SL \i48/i75  (.A(\i48/n480 ),
    .B(\i48/n251 ),
    .C(\i48/n187 ),
    .D(\i48/n500 ),
    .E(\i48/n520 ),
    .Y(\i48/n380 ));
 NOR3xp33_ASAP7_75t_SL \i48/i76  (.A(\i48/n352 ),
    .B(\i48/n270 ),
    .C(\i48/n263 ),
    .Y(\i48/n379 ));
 NOR2xp33_ASAP7_75t_SL \i48/i77  (.A(\i48/n309 ),
    .B(\i48/n330 ),
    .Y(\i48/n378 ));
 NOR2xp33_ASAP7_75t_SL \i48/i78  (.A(\i48/n350 ),
    .B(\i48/n300 ),
    .Y(\i48/n377 ));
 NOR2x1_ASAP7_75t_SL \i48/i79  (.A(\i48/n314 ),
    .B(\i48/n286 ),
    .Y(\i48/n388 ));
 AND5x2_ASAP7_75t_SL \i48/i8  (.A(\i48/n437 ),
    .B(\i48/n417 ),
    .C(\i48/n430 ),
    .D(\i48/n428 ),
    .E(\i48/n409 ),
    .Y(n24[6]));
 NAND3xp33_ASAP7_75t_SL \i48/i80  (.A(\i48/n260 ),
    .B(\i48/n574 ),
    .C(\i48/n497 ),
    .Y(\i48/n376 ));
 NAND2xp5_ASAP7_75t_L \i48/i81  (.A(\i48/n349 ),
    .B(\i48/n318 ),
    .Y(\i48/n375 ));
 NAND2xp5_ASAP7_75t_SL \i48/i82  (.A(\i48/n299 ),
    .B(\i48/n340 ),
    .Y(\i48/n374 ));
 NAND3xp33_ASAP7_75t_SL \i48/i83  (.A(\i48/n302 ),
    .B(\i48/n246 ),
    .C(\i48/n231 ),
    .Y(\i48/n387 ));
 NOR3xp33_ASAP7_75t_SL \i48/i84  (.A(\i48/n492 ),
    .B(\i48/n7 ),
    .C(\i48/n466 ),
    .Y(\i48/n373 ));
 NAND2xp5_ASAP7_75t_SL \i48/i85  (.A(\i48/n490 ),
    .B(\i48/n329 ),
    .Y(\i48/n386 ));
 OR3x1_ASAP7_75t_SL \i48/i86  (.A(\i48/n254 ),
    .B(\i48/n265 ),
    .C(\i48/n22 ),
    .Y(\i48/n372 ));
 NOR2x1_ASAP7_75t_SL \i48/i87  (.A(\i48/n263 ),
    .B(\i48/n352 ),
    .Y(\i48/n385 ));
 NOR2xp33_ASAP7_75t_L \i48/i88  (.A(\i48/n311 ),
    .B(\i48/n297 ),
    .Y(\i48/n384 ));
 NOR2xp33_ASAP7_75t_SL \i48/i89  (.A(\i48/n339 ),
    .B(\i48/n459 ),
    .Y(\i48/n382 ));
 AND3x4_ASAP7_75t_SL \i48/i9  (.A(\i48/n437 ),
    .B(\i48/n446 ),
    .C(\i48/n425 ),
    .Y(n24[1]));
 NOR3x1_ASAP7_75t_SL \i48/i90  (.A(\i48/n259 ),
    .B(\i48/n170 ),
    .C(\i48/n303 ),
    .Y(\i48/n381 ));
 NOR3xp33_ASAP7_75t_SL \i48/i91  (.A(\i48/n267 ),
    .B(\i48/n193 ),
    .C(\i48/n257 ),
    .Y(\i48/n368 ));
 NOR2xp33_ASAP7_75t_SL \i48/i92  (.A(\i48/n579 ),
    .B(\i48/n324 ),
    .Y(\i48/n367 ));
 NAND3xp33_ASAP7_75t_SL \i48/i93  (.A(\i48/n253 ),
    .B(\i48/n316 ),
    .C(\i48/n264 ),
    .Y(\i48/n366 ));
 NAND4xp25_ASAP7_75t_SL \i48/i94  (.A(\i48/n562 ),
    .B(\i48/n250 ),
    .C(\i48/n275 ),
    .D(\i48/n485 ),
    .Y(\i48/n365 ));
 NAND2xp5_ASAP7_75t_SL \i48/i95  (.A(\i48/n338 ),
    .B(\i48/n351 ),
    .Y(\i48/n371 ));
 NOR5xp2_ASAP7_75t_SL \i48/i96  (.A(\i48/n347 ),
    .B(\i48/n479 ),
    .C(\i48/n104 ),
    .D(\i48/n207 ),
    .E(\i48/n143 ),
    .Y(\i48/n364 ));
 NAND3xp33_ASAP7_75t_SL \i48/i97  (.A(\i48/n301 ),
    .B(\i48/n322 ),
    .C(\i48/n496 ),
    .Y(\i48/n363 ));
 NAND2xp33_ASAP7_75t_SL \i48/i98  (.A(\i48/n247 ),
    .B(\i48/n344 ),
    .Y(\i48/n362 ));
 NOR5xp2_ASAP7_75t_SL \i48/i99  (.A(\i48/n287 ),
    .B(\i48/n459 ),
    .C(\i48/n274 ),
    .D(\i48/n229 ),
    .E(\i48/n184 ),
    .Y(\i48/n361 ));
 XOR2xp5_ASAP7_75t_SL i480 (.A(n799),
    .B(n597),
    .Y(n992));
 XNOR2xp5_ASAP7_75t_SL i481 (.A(n598),
    .B(n596),
    .Y(n991));
 XOR2xp5_ASAP7_75t_SL i482 (.A(n491),
    .B(n600),
    .Y(n990));
 AOI22xp5_ASAP7_75t_SL i483 (.A1(n839),
    .A2(n781),
    .B1(n840),
    .B2(n782),
    .Y(n989));
 XOR2xp5_ASAP7_75t_SL i484 (.A(n601),
    .B(n604),
    .Y(n988));
 XOR2xp5_ASAP7_75t_SL i485 (.A(n607),
    .B(n608),
    .Y(n987));
 XNOR2xp5_ASAP7_75t_SL i486 (.A(n610),
    .B(n609),
    .Y(n986));
 AOI22xp5_ASAP7_75t_SL i487 (.A1(n509),
    .A2(n855),
    .B1(n508),
    .B2(n856),
    .Y(n985));
 XOR2xp5_ASAP7_75t_SL i488 (.A(n625),
    .B(n622),
    .Y(n984));
 XOR2xp5_ASAP7_75t_SL i489 (.A(n1173),
    .B(n615),
    .Y(n983));
 INVx2_ASAP7_75t_SL \i49/i0  (.A(n23[2]),
    .Y(\i49/n0 ));
 INVx2_ASAP7_75t_SL \i49/i1  (.A(n23[0]),
    .Y(\i49/n1 ));
 NOR2x1p5_ASAP7_75t_SL \i49/i10  (.A(\i49/n516 ),
    .B(\i49/n507 ),
    .Y(n22[5]));
 NAND2xp33_ASAP7_75t_SL \i49/i100  (.A(\i49/n304 ),
    .B(\i49/n409 ),
    .Y(\i49/n429 ));
 NOR5xp2_ASAP7_75t_SL \i49/i101  (.A(\i49/n350 ),
    .B(\i49/n554 ),
    .C(\i49/n334 ),
    .D(\i49/n278 ),
    .E(\i49/n225 ),
    .Y(\i49/n428 ));
 NAND5xp2_ASAP7_75t_SL \i49/i102  (.A(\i49/n570 ),
    .B(\i49/n365 ),
    .C(\i49/n567 ),
    .D(\i49/n332 ),
    .E(\i49/n274 ),
    .Y(\i49/n427 ));
 NAND3xp33_ASAP7_75t_L \i49/i103  (.A(\i49/n283 ),
    .B(\i49/n317 ),
    .C(\i49/n392 ),
    .Y(\i49/n426 ));
 NOR5xp2_ASAP7_75t_SL \i49/i104  (.A(\i49/n281 ),
    .B(\i49/n295 ),
    .C(\i49/n272 ),
    .D(\i49/n118 ),
    .E(\i49/n556 ),
    .Y(\i49/n425 ));
 NAND5xp2_ASAP7_75t_SL \i49/i105  (.A(\i49/n26 ),
    .B(\i49/n366 ),
    .C(\i49/n567 ),
    .D(\i49/n540 ),
    .E(\i49/n195 ),
    .Y(\i49/n424 ));
 NAND4xp25_ASAP7_75t_SL \i49/i106  (.A(\i49/n219 ),
    .B(\i49/n233 ),
    .C(\i49/n338 ),
    .D(\i49/n19 ),
    .Y(\i49/n423 ));
 NOR5xp2_ASAP7_75t_SL \i49/i107  (.A(\i49/n239 ),
    .B(\i49/n286 ),
    .C(\i49/n224 ),
    .D(\i49/n189 ),
    .E(\i49/n188 ),
    .Y(\i49/n422 ));
 NOR2xp33_ASAP7_75t_SL \i49/i108  (.A(\i49/n382 ),
    .B(\i49/n416 ),
    .Y(\i49/n421 ));
 NOR2xp33_ASAP7_75t_SL \i49/i109  (.A(\i49/n370 ),
    .B(\i49/n401 ),
    .Y(\i49/n420 ));
 AND2x2_ASAP7_75t_SL \i49/i11  (.A(\i49/n517 ),
    .B(\i49/n500 ),
    .Y(n22[0]));
 NAND3x2_ASAP7_75t_SL \i49/i110  (.B(\i49/n365 ),
    .C(\i49/n399 ),
    .Y(\i49/n437 ),
    .A(\i49/n237 ));
 NAND3x1_ASAP7_75t_SL \i49/i111  (.A(\i49/n360 ),
    .B(\i49/n339 ),
    .C(\i49/n305 ),
    .Y(\i49/n436 ));
 AOI21xp5_ASAP7_75t_L \i49/i112  (.A1(\i49/n74 ),
    .A2(\i49/n242 ),
    .B(\i49/n166 ),
    .Y(\i49/n412 ));
 NOR2xp33_ASAP7_75t_SL \i49/i113  (.A(\i49/n309 ),
    .B(\i49/n350 ),
    .Y(\i49/n411 ));
 NAND2xp5_ASAP7_75t_SL \i49/i114  (.A(\i49/n337 ),
    .B(\i49/n369 ),
    .Y(\i49/n410 ));
 NOR2xp33_ASAP7_75t_SL \i49/i115  (.A(\i49/n368 ),
    .B(\i49/n28 ),
    .Y(\i49/n409 ));
 NOR2xp33_ASAP7_75t_SL \i49/i116  (.A(\i49/n345 ),
    .B(\i49/n355 ),
    .Y(\i49/n408 ));
 NOR2xp67_ASAP7_75t_SL \i49/i117  (.A(\i49/n175 ),
    .B(\i49/n352 ),
    .Y(\i49/n407 ));
 NOR2xp33_ASAP7_75t_SL \i49/i118  (.A(\i49/n22 ),
    .B(\i49/n350 ),
    .Y(\i49/n406 ));
 NOR4xp25_ASAP7_75t_SL \i49/i119  (.A(\i49/n320 ),
    .B(\i49/n24 ),
    .C(\i49/n22 ),
    .D(\i49/n184 ),
    .Y(\i49/n405 ));
 NOR3xp33_ASAP7_75t_SL \i49/i12  (.A(\i49/n489 ),
    .B(\i49/n485 ),
    .C(\i49/n492 ),
    .Y(\i49/n517 ));
 NAND2xp5_ASAP7_75t_SL \i49/i120  (.A(\i49/n560 ),
    .B(\i49/n329 ),
    .Y(\i49/n404 ));
 NOR4xp25_ASAP7_75t_SL \i49/i121  (.A(\i49/n115 ),
    .B(\i49/n261 ),
    .C(\i49/n227 ),
    .D(\i49/n243 ),
    .Y(\i49/n403 ));
 NOR3xp33_ASAP7_75t_SL \i49/i122  (.A(\i49/n266 ),
    .B(\i49/n553 ),
    .C(\i49/n265 ),
    .Y(\i49/n402 ));
 NAND2xp33_ASAP7_75t_SL \i49/i123  (.A(\i49/n316 ),
    .B(\i49/n23 ),
    .Y(\i49/n401 ));
 NOR2xp33_ASAP7_75t_SL \i49/i124  (.A(\i49/n309 ),
    .B(\i49/n311 ),
    .Y(\i49/n400 ));
 NOR2x1p5_ASAP7_75t_SL \i49/i125  (.A(\i49/n290 ),
    .B(\i49/n315 ),
    .Y(\i49/n399 ));
 NAND2xp33_ASAP7_75t_SL \i49/i126  (.A(\i49/n367 ),
    .B(\i49/n349 ),
    .Y(\i49/n398 ));
 NAND3xp33_ASAP7_75t_SL \i49/i127  (.A(\i49/n25 ),
    .B(\i49/n525 ),
    .C(\i49/n249 ),
    .Y(\i49/n397 ));
 NOR3xp33_ASAP7_75t_SL \i49/i128  (.A(\i49/n220 ),
    .B(\i49/n234 ),
    .C(\i49/n205 ),
    .Y(\i49/n419 ));
 NAND2xp5_ASAP7_75t_SL \i49/i129  (.A(\i49/n13 ),
    .B(\i49/n219 ),
    .Y(\i49/n418 ));
 NOR2x2_ASAP7_75t_SL \i49/i13  (.A(\i49/n509 ),
    .B(\i49/n510 ),
    .Y(n22[2]));
 NOR2x1_ASAP7_75t_SL \i49/i130  (.A(\i49/n289 ),
    .B(\i49/n313 ),
    .Y(\i49/n417 ));
 NAND2xp5_ASAP7_75t_SL \i49/i131  (.A(\i49/n567 ),
    .B(\i49/n321 ),
    .Y(\i49/n416 ));
 NOR2x1_ASAP7_75t_SL \i49/i132  (.A(\i49/n291 ),
    .B(\i49/n353 ),
    .Y(\i49/n415 ));
 NOR2x1_ASAP7_75t_SL \i49/i133  (.A(\i49/n24 ),
    .B(\i49/n309 ),
    .Y(\i49/n414 ));
 NOR3x1_ASAP7_75t_SL \i49/i134  (.A(\i49/n224 ),
    .B(\i49/n215 ),
    .C(\i49/n186 ),
    .Y(\i49/n413 ));
 INVx1_ASAP7_75t_SL \i49/i135  (.A(\i49/n394 ),
    .Y(\i49/n395 ));
 INVx1_ASAP7_75t_SL \i49/i136  (.A(\i49/n29 ),
    .Y(\i49/n393 ));
 NOR4xp25_ASAP7_75t_SL \i49/i137  (.A(\i49/n208 ),
    .B(\i49/n246 ),
    .C(\i49/n232 ),
    .D(\i49/n201 ),
    .Y(\i49/n392 ));
 AOI211xp5_ASAP7_75t_SL \i49/i138  (.A1(\i49/n536 ),
    .A2(\i49/n69 ),
    .B(\i49/n315 ),
    .C(\i49/n180 ),
    .Y(\i49/n391 ));
 AOI211xp5_ASAP7_75t_SL \i49/i139  (.A1(\i49/n121 ),
    .A2(\i49/n56 ),
    .B(\i49/n333 ),
    .C(\i49/n264 ),
    .Y(\i49/n390 ));
 NAND4xp75_ASAP7_75t_SL \i49/i14  (.A(\i49/n475 ),
    .B(\i49/n495 ),
    .C(\i49/n473 ),
    .D(\i49/n573 ),
    .Y(\i49/n516 ));
 NAND2xp33_ASAP7_75t_L \i49/i140  (.A(\i49/n306 ),
    .B(\i49/n331 ),
    .Y(\i49/n389 ));
 NAND5xp2_ASAP7_75t_SL \i49/i141  (.A(\i49/n244 ),
    .B(\i49/n259 ),
    .C(\i49/n270 ),
    .D(\i49/n182 ),
    .E(\i49/n116 ),
    .Y(\i49/n388 ));
 OAI221xp5_ASAP7_75t_SL \i49/i142  (.A1(\i49/n119 ),
    .A2(\i49/n90 ),
    .B1(\i49/n119 ),
    .B2(\i49/n17 ),
    .C(\i49/n316 ),
    .Y(\i49/n387 ));
 NOR2xp33_ASAP7_75t_SL \i49/i143  (.A(\i49/n296 ),
    .B(\i49/n300 ),
    .Y(\i49/n386 ));
 AOI211xp5_ASAP7_75t_SL \i49/i144  (.A1(\i49/n170 ),
    .A2(\i49/n532 ),
    .B(\i49/n280 ),
    .C(\i49/n191 ),
    .Y(\i49/n385 ));
 OA21x2_ASAP7_75t_SL \i49/i145  (.A1(\i49/n522 ),
    .A2(\i49/n74 ),
    .B(\i49/n366 ),
    .Y(\i49/n384 ));
 NOR4xp25_ASAP7_75t_SL \i49/i146  (.A(\i49/n273 ),
    .B(\i49/n179 ),
    .C(\i49/n212 ),
    .D(\i49/n186 ),
    .Y(\i49/n383 ));
 NAND5xp2_ASAP7_75t_SL \i49/i147  (.A(\i49/n149 ),
    .B(\i49/n105 ),
    .C(\i49/n160 ),
    .D(\i49/n151 ),
    .E(\i49/n97 ),
    .Y(\i49/n382 ));
 NOR3xp33_ASAP7_75t_SL \i49/i148  (.A(\i49/n314 ),
    .B(\i49/n181 ),
    .C(\i49/n95 ),
    .Y(\i49/n381 ));
 NAND2xp5_ASAP7_75t_SL \i49/i149  (.A(\i49/n294 ),
    .B(\i49/n26 ),
    .Y(\i49/n380 ));
 NOR3xp33_ASAP7_75t_SL \i49/i15  (.A(\i49/n493 ),
    .B(\i49/n458 ),
    .C(\i49/n503 ),
    .Y(\i49/n515 ));
 NAND5xp2_ASAP7_75t_SL \i49/i150  (.A(\i49/n542 ),
    .B(\i49/n111 ),
    .C(\i49/n524 ),
    .D(\i49/n200 ),
    .E(\i49/n199 ),
    .Y(\i49/n379 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i49/i151  (.A1(\i49/n537 ),
    .A2(\i49/n100 ),
    .B(\i49/n79 ),
    .C(\i49/n285 ),
    .Y(\i49/n378 ));
 NAND4xp25_ASAP7_75t_SL \i49/i152  (.A(\i49/n327 ),
    .B(\i49/n260 ),
    .C(\i49/n117 ),
    .D(\i49/n183 ),
    .Y(\i49/n377 ));
 NAND5xp2_ASAP7_75t_SL \i49/i153  (.A(\i49/n171 ),
    .B(\i49/n150 ),
    .C(\i49/n251 ),
    .D(\i49/n113 ),
    .E(\i49/n108 ),
    .Y(\i49/n376 ));
 NAND2xp5_ASAP7_75t_SL \i49/i154  (.A(\i49/n293 ),
    .B(\i49/n319 ),
    .Y(\i49/n375 ));
 NAND3xp33_ASAP7_75t_SL \i49/i155  (.A(\i49/n312 ),
    .B(\i49/n96 ),
    .C(\i49/n102 ),
    .Y(\i49/n374 ));
 NAND2xp5_ASAP7_75t_SL \i49/i156  (.A(\i49/n237 ),
    .B(\i49/n365 ),
    .Y(\i49/n373 ));
 NOR2xp33_ASAP7_75t_L \i49/i157  (.A(\i49/n343 ),
    .B(\i49/n355 ),
    .Y(\i49/n396 ));
 NAND2xp5_ASAP7_75t_SL \i49/i158  (.A(\i49/n238 ),
    .B(\i49/n367 ),
    .Y(\i49/n372 ));
 NOR2x1_ASAP7_75t_SL \i49/i159  (.A(\i49/n298 ),
    .B(\i49/n347 ),
    .Y(\i49/n394 ));
 NAND4xp75_ASAP7_75t_SL \i49/i16  (.A(\i49/n474 ),
    .B(\i49/n505 ),
    .C(\i49/n479 ),
    .D(\i49/n469 ),
    .Y(\i49/n514 ));
 NAND3x1_ASAP7_75t_SL \i49/i160  (.A(\i49/n277 ),
    .B(\i49/n142 ),
    .C(\i49/n154 ),
    .Y(\i49/n29 ));
 INVxp67_ASAP7_75t_SL \i49/i161  (.A(\i49/n370 ),
    .Y(\i49/n371 ));
 INVxp67_ASAP7_75t_SL \i49/i162  (.A(\i49/n7 ),
    .Y(\i49/n369 ));
 INVxp67_ASAP7_75t_SL \i49/i163  (.A(\i49/n363 ),
    .Y(\i49/n364 ));
 INVxp67_ASAP7_75t_SL \i49/i164  (.A(\i49/n361 ),
    .Y(\i49/n362 ));
 INVx1_ASAP7_75t_SL \i49/i165  (.A(\i49/n359 ),
    .Y(\i49/n360 ));
 INVxp67_ASAP7_75t_SL \i49/i166  (.A(\i49/n357 ),
    .Y(\i49/n358 ));
 INVxp67_ASAP7_75t_SL \i49/i167  (.A(\i49/n353 ),
    .Y(\i49/n354 ));
 INVxp67_ASAP7_75t_SL \i49/i168  (.A(\i49/n27 ),
    .Y(\i49/n351 ));
 OAI31xp33_ASAP7_75t_SL \i49/i169  (.A1(\i49/n532 ),
    .A2(\i49/n3 ),
    .A3(\i49/n57 ),
    .B(\i49/n53 ),
    .Y(\i49/n348 ));
 AND3x2_ASAP7_75t_SL \i49/i17  (.A(\i49/n496 ),
    .B(\i49/n511 ),
    .C(\i49/n501 ),
    .Y(n22[7]));
 NAND2xp5_ASAP7_75t_SL \i49/i170  (.A(\i49/n564 ),
    .B(\i49/n229 ),
    .Y(\i49/n347 ));
 NOR2xp33_ASAP7_75t_SL \i49/i171  (.A(\i49/n271 ),
    .B(\i49/n266 ),
    .Y(\i49/n346 ));
 NAND2xp33_ASAP7_75t_SL \i49/i172  (.A(\i49/n525 ),
    .B(\i49/n567 ),
    .Y(\i49/n345 ));
 OAI21xp5_ASAP7_75t_SL \i49/i173  (.A1(\i49/n55 ),
    .A2(\i49/n546 ),
    .B(\i49/n197 ),
    .Y(\i49/n344 ));
 NAND2xp5_ASAP7_75t_SL \i49/i174  (.A(\i49/n185 ),
    .B(\i49/n525 ),
    .Y(\i49/n343 ));
 AOI211xp5_ASAP7_75t_SL \i49/i175  (.A1(\i49/n88 ),
    .A2(\i49/n33 ),
    .B(\i49/n122 ),
    .C(\i49/n128 ),
    .Y(\i49/n342 ));
 AOI31xp33_ASAP7_75t_SL \i49/i176  (.A1(\i49/n55 ),
    .A2(\i49/n18 ),
    .A3(\i49/n64 ),
    .B(\i49/n49 ),
    .Y(\i49/n341 ));
 NOR3xp33_ASAP7_75t_SL \i49/i177  (.A(\i49/n553 ),
    .B(\i49/n139 ),
    .C(\i49/n127 ),
    .Y(\i49/n340 ));
 NOR3xp33_ASAP7_75t_SL \i49/i178  (.A(\i49/n120 ),
    .B(\i49/n569 ),
    .C(\i49/n271 ),
    .Y(\i49/n339 ));
 OAI31xp33_ASAP7_75t_SL \i49/i179  (.A1(\i49/n51 ),
    .A2(\i49/n53 ),
    .A3(\i49/n72 ),
    .B(\i49/n88 ),
    .Y(\i49/n338 ));
 NAND4xp75_ASAP7_75t_SL \i49/i18  (.A(\i49/n572 ),
    .B(\i49/n478 ),
    .C(\i49/n487 ),
    .D(\i49/n504 ),
    .Y(\i49/n513 ));
 AOI221xp5_ASAP7_75t_SL \i49/i180  (.A1(\i49/n537 ),
    .A2(\i49/n91 ),
    .B1(\i49/n58 ),
    .B2(\i49/n66 ),
    .C(\i49/n202 ),
    .Y(\i49/n337 ));
 OAI31xp33_ASAP7_75t_R \i49/i181  (.A1(\i49/n532 ),
    .A2(\i49/n76 ),
    .A3(\i49/n537 ),
    .B(\i49/n72 ),
    .Y(\i49/n336 ));
 AOI21xp5_ASAP7_75t_SL \i49/i182  (.A1(\i49/n166 ),
    .A2(\i49/n64 ),
    .B(\i49/n86 ),
    .Y(\i49/n370 ));
 AOI21xp5_ASAP7_75t_L \i49/i183  (.A1(\i49/n64 ),
    .A2(\i49/n176 ),
    .B(\i49/n85 ),
    .Y(\i49/n335 ));
 OAI221xp5_ASAP7_75t_SL \i49/i184  (.A1(\i49/n534 ),
    .A2(\i49/n90 ),
    .B1(\i49/n52 ),
    .B2(\i49/n60 ),
    .C(\i49/n226 ),
    .Y(\i49/n334 ));
 AOI21xp33_ASAP7_75t_SL \i49/i185  (.A1(\i49/n176 ),
    .A2(\i49/n50 ),
    .B(\i49/n77 ),
    .Y(\i49/n333 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i49/i186  (.A1(\i49/n83 ),
    .A2(\i49/n5 ),
    .B(\i49/n87 ),
    .C(\i49/n20 ),
    .Y(\i49/n332 ));
 NOR3xp33_ASAP7_75t_SL \i49/i187  (.A(\i49/n240 ),
    .B(\i49/n120 ),
    .C(\i49/n146 ),
    .Y(\i49/n331 ));
 NAND3xp33_ASAP7_75t_SL \i49/i188  (.A(\i49/n548 ),
    .B(\i49/n545 ),
    .C(\i49/n174 ),
    .Y(\i49/n330 ));
 AOI22xp5_ASAP7_75t_SL \i49/i189  (.A1(\i49/n552 ),
    .A2(\i49/n162 ),
    .B1(\i49/n66 ),
    .B2(\i49/n57 ),
    .Y(\i49/n329 ));
 NAND2x1_ASAP7_75t_SL \i49/i19  (.A(\i49/n466 ),
    .B(\i49/n497 ),
    .Y(\i49/n512 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i49/i190  (.A1(\i49/n85 ),
    .A2(\i49/n54 ),
    .B(\i49/n71 ),
    .C(\i49/n123 ),
    .Y(\i49/n328 ));
 OAI21xp33_ASAP7_75t_SL \i49/i191  (.A1(\i49/n63 ),
    .A2(\i49/n168 ),
    .B(\i49/n532 ),
    .Y(\i49/n327 ));
 NAND4xp25_ASAP7_75t_SL \i49/i192  (.A(\i49/n562 ),
    .B(\i49/n183 ),
    .C(\i49/n152 ),
    .D(\i49/n155 ),
    .Y(\i49/n326 ));
 NAND2xp33_ASAP7_75t_SL \i49/i193  (.A(\i49/n254 ),
    .B(\i49/n145 ),
    .Y(\i49/n325 ));
 OAI211xp5_ASAP7_75t_SL \i49/i194  (.A1(\i49/n70 ),
    .A2(\i49/n77 ),
    .B(\i49/n157 ),
    .C(\i49/n161 ),
    .Y(\i49/n368 ));
 NOR2xp67_ASAP7_75t_SL \i49/i195  (.A(\i49/n216 ),
    .B(\i49/n272 ),
    .Y(\i49/n367 ));
 AO21x1_ASAP7_75t_SL \i49/i196  (.A1(\i49/n59 ),
    .A2(\i49/n165 ),
    .B(\i49/n147 ),
    .Y(\i49/n366 ));
 AOI21x1_ASAP7_75t_SL \i49/i197  (.A1(\i49/n57 ),
    .A2(\i49/n63 ),
    .B(\i49/n280 ),
    .Y(\i49/n365 ));
 NAND2xp5_ASAP7_75t_SL \i49/i198  (.A(\i49/n256 ),
    .B(\i49/n231 ),
    .Y(\i49/n28 ));
 NOR2xp33_ASAP7_75t_SL \i49/i199  (.A(\i49/n257 ),
    .B(\i49/n273 ),
    .Y(\i49/n363 ));
 INVx1_ASAP7_75t_SL \i49/i2  (.A(\i49/n448 ),
    .Y(\i49/n2 ));
 NOR2xp33_ASAP7_75t_SL \i49/i20  (.A(\i49/n498 ),
    .B(\i49/n459 ),
    .Y(\i49/n511 ));
 OAI211xp5_ASAP7_75t_SL \i49/i200  (.A1(\i49/n64 ),
    .A2(\i49/n77 ),
    .B(\i49/n197 ),
    .C(\i49/n198 ),
    .Y(\i49/n361 ));
 OR2x2_ASAP7_75t_SL \i49/i201  (.A(\i49/n210 ),
    .B(\i49/n230 ),
    .Y(\i49/n359 ));
 AOI21xp5_ASAP7_75t_SL \i49/i202  (.A1(\i49/n76 ),
    .A2(\i49/n65 ),
    .B(\i49/n269 ),
    .Y(\i49/n357 ));
 OAI211xp5_ASAP7_75t_SL \i49/i203  (.A1(\i49/n90 ),
    .A2(\i49/n541 ),
    .B(\i49/n193 ),
    .C(\i49/n135 ),
    .Y(\i49/n356 ));
 NAND2xp5_ASAP7_75t_SL \i49/i204  (.A(\i49/n274 ),
    .B(\i49/n275 ),
    .Y(\i49/n355 ));
 NAND2xp5_ASAP7_75t_SL \i49/i205  (.A(\i49/n25 ),
    .B(\i49/n544 ),
    .Y(\i49/n353 ));
 NAND2xp5_ASAP7_75t_SL \i49/i206  (.A(\i49/n253 ),
    .B(\i49/n543 ),
    .Y(\i49/n352 ));
 OAI221xp5_ASAP7_75t_SL \i49/i207  (.A1(\i49/n60 ),
    .A2(\i49/n67 ),
    .B1(\i49/n55 ),
    .B2(\i49/n59 ),
    .C(\i49/n526 ),
    .Y(\i49/n27 ));
 NAND2xp5_ASAP7_75t_SL \i49/i208  (.A(\i49/n190 ),
    .B(\i49/n214 ),
    .Y(\i49/n350 ));
 NOR2x1_ASAP7_75t_SL \i49/i209  (.A(\i49/n255 ),
    .B(\i49/n225 ),
    .Y(\i49/n349 ));
 NAND4xp75_ASAP7_75t_SL \i49/i21  (.A(\i49/n470 ),
    .B(\i49/n482 ),
    .C(\i49/n464 ),
    .D(\i49/n467 ),
    .Y(\i49/n510 ));
 INVxp67_ASAP7_75t_SL \i49/i210  (.A(\i49/n320 ),
    .Y(\i49/n321 ));
 INVx1_ASAP7_75t_SL \i49/i211  (.A(\i49/n317 ),
    .Y(\i49/n318 ));
 INVx1_ASAP7_75t_SL \i49/i212  (.A(\i49/n312 ),
    .Y(\i49/n313 ));
 NAND4xp25_ASAP7_75t_SL \i49/i213  (.A(\i49/n529 ),
    .B(\i49/n547 ),
    .C(\i49/n123 ),
    .D(\i49/n528 ),
    .Y(\i49/n308 ));
 AOI31xp33_ASAP7_75t_SL \i49/i214  (.A1(\i49/n136 ),
    .A2(\i49/n74 ),
    .A3(\i49/n49 ),
    .B(\i49/n50 ),
    .Y(\i49/n307 ));
 NOR4xp25_ASAP7_75t_SL \i49/i215  (.A(\i49/n115 ),
    .B(\i49/n129 ),
    .C(\i49/n196 ),
    .D(\i49/n94 ),
    .Y(\i49/n306 ));
 AOI211xp5_ASAP7_75t_SL \i49/i216  (.A1(\i49/n137 ),
    .A2(\i49/n81 ),
    .B(\i49/n181 ),
    .C(\i49/n103 ),
    .Y(\i49/n305 ));
 AOI21xp5_ASAP7_75t_SL \i49/i217  (.A1(\i49/n167 ),
    .A2(\i49/n87 ),
    .B(\i49/n245 ),
    .Y(\i49/n304 ));
 NOR2xp33_ASAP7_75t_L \i49/i218  (.A(\i49/n204 ),
    .B(\i49/n267 ),
    .Y(\i49/n303 ));
 OAI31xp33_ASAP7_75t_SL \i49/i219  (.A1(\i49/n552 ),
    .A2(\i49/n58 ),
    .A3(\i49/n88 ),
    .B(\i49/n65 ),
    .Y(\i49/n302 ));
 OR3x1_ASAP7_75t_SL \i49/i22  (.A(\i49/n490 ),
    .B(\i49/n488 ),
    .C(\i49/n471 ),
    .Y(\i49/n509 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i49/i220  (.A1(\i49/n77 ),
    .A2(\i49/n54 ),
    .B(\i49/n82 ),
    .C(\i49/n241 ),
    .Y(\i49/n301 ));
 OAI22xp5_ASAP7_75t_SL \i49/i221  (.A1(\i49/n541 ),
    .A2(\i49/n169 ),
    .B1(\i49/n70 ),
    .B2(\i49/n101 ),
    .Y(\i49/n300 ));
 NOR2xp33_ASAP7_75t_SL \i49/i222  (.A(\i49/n222 ),
    .B(\i49/n206 ),
    .Y(\i49/n299 ));
 OAI222xp33_ASAP7_75t_SL \i49/i223  (.A1(\i49/n85 ),
    .A2(\i49/n50 ),
    .B1(\i49/n54 ),
    .B2(\i49/n18 ),
    .C1(\i49/n74 ),
    .C2(\i49/n70 ),
    .Y(\i49/n298 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i49/i224  (.A1(\i49/n552 ),
    .A2(\i49/n61 ),
    .B(\i49/n5 ),
    .C(\i49/n178 ),
    .Y(\i49/n297 ));
 NAND2xp33_ASAP7_75t_L \i49/i225  (.A(\i49/n530 ),
    .B(\i49/n559 ),
    .Y(\i49/n296 ));
 NAND2xp33_ASAP7_75t_SL \i49/i226  (.A(\i49/n263 ),
    .B(\i49/n134 ),
    .Y(\i49/n295 ));
 AOI22xp5_ASAP7_75t_SL \i49/i227  (.A1(\i49/n76 ),
    .A2(\i49/n112 ),
    .B1(\i49/n81 ),
    .B2(\i49/n537 ),
    .Y(\i49/n294 ));
 OAI21xp33_ASAP7_75t_L \i49/i228  (.A1(\i49/n121 ),
    .A2(\i49/n76 ),
    .B(\i49/n81 ),
    .Y(\i49/n293 ));
 OA21x2_ASAP7_75t_SL \i49/i229  (.A1(\i49/n50 ),
    .A2(\i49/n546 ),
    .B(\i49/n565 ),
    .Y(\i49/n292 ));
 OR3x1_ASAP7_75t_SL \i49/i23  (.A(\i49/n491 ),
    .B(\i49/n457 ),
    .C(\i49/n430 ),
    .Y(\i49/n508 ));
 NAND2xp5_ASAP7_75t_SL \i49/i230  (.A(\i49/n211 ),
    .B(\i49/n279 ),
    .Y(\i49/n291 ));
 NAND4xp25_ASAP7_75t_SL \i49/i231  (.A(\i49/n132 ),
    .B(\i49/n156 ),
    .C(\i49/n110 ),
    .D(\i49/n107 ),
    .Y(\i49/n290 ));
 OAI221xp5_ASAP7_75t_SL \i49/i232  (.A1(\i49/n89 ),
    .A2(\i49/n82 ),
    .B1(\i49/n73 ),
    .B2(\i49/n17 ),
    .C(\i49/n114 ),
    .Y(\i49/n324 ));
 OAI222xp33_ASAP7_75t_SL \i49/i233  (.A1(\i49/n8 ),
    .A2(\i49/n55 ),
    .B1(\i49/n60 ),
    .B2(\i49/n70 ),
    .C1(\i49/n73 ),
    .C2(\i49/n78 ),
    .Y(\i49/n289 ));
 OAI221xp5_ASAP7_75t_SL \i49/i234  (.A1(\i49/n85 ),
    .A2(\i49/n78 ),
    .B1(\i49/n73 ),
    .B2(\i49/n71 ),
    .C(\i49/n223 ),
    .Y(\i49/n288 ));
 AND3x1_ASAP7_75t_SL \i49/i235  (.A(\i49/n130 ),
    .B(\i49/n547 ),
    .C(\i49/n247 ),
    .Y(\i49/n287 ));
 AOI22xp5_ASAP7_75t_SL \i49/i236  (.A1(\i49/n84 ),
    .A2(\i49/n164 ),
    .B1(\i49/n63 ),
    .B2(\i49/n87 ),
    .Y(\i49/n323 ));
 AOI31xp33_ASAP7_75t_SL \i49/i237  (.A1(\i49/n55 ),
    .A2(\i49/n80 ),
    .A3(\i49/n71 ),
    .B(\i49/n59 ),
    .Y(\i49/n286 ));
 NAND2xp33_ASAP7_75t_SL \i49/i238  (.A(\i49/n563 ),
    .B(\i49/n248 ),
    .Y(\i49/n285 ));
 OAI221xp5_ASAP7_75t_SL \i49/i239  (.A1(\i49/n85 ),
    .A2(\i49/n80 ),
    .B1(\i49/n534 ),
    .B2(\i49/n18 ),
    .C(\i49/n262 ),
    .Y(\i49/n284 ));
 NAND3xp33_ASAP7_75t_SL \i49/i24  (.A(\i49/n502 ),
    .B(\i49/n487 ),
    .C(\i49/n470 ),
    .Y(\i49/n507 ));
 OAI222xp33_ASAP7_75t_SL \i49/i240  (.A1(\i49/n541 ),
    .A2(\i49/n80 ),
    .B1(\i49/n89 ),
    .B2(\i49/n78 ),
    .C1(\i49/n534 ),
    .C2(\i49/n64 ),
    .Y(\i49/n322 ));
 NAND3x1_ASAP7_75t_SL \i49/i241  (.A(\i49/n523 ),
    .B(\i49/n159 ),
    .C(\i49/n153 ),
    .Y(\i49/n320 ));
 AOI22x1_ASAP7_75t_SL \i49/i242  (.A1(\i49/n158 ),
    .A2(\i49/n88 ),
    .B1(\i49/n58 ),
    .B2(\i49/n72 ),
    .Y(\i49/n13 ));
 AOI22xp5_ASAP7_75t_SL \i49/i243  (.A1(\i49/n91 ),
    .A2(\i49/n555 ),
    .B1(\i49/n51 ),
    .B2(\i49/n532 ),
    .Y(\i49/n319 ));
 AOI221x1_ASAP7_75t_SL \i49/i244  (.A1(\i49/n88 ),
    .A2(\i49/n72 ),
    .B1(\i49/n537 ),
    .B2(\i49/n79 ),
    .C(\i49/n250 ),
    .Y(\i49/n317 ));
 AOI211x1_ASAP7_75t_SL \i49/i245  (.A1(\i49/n106 ),
    .A2(\i49/n68 ),
    .B(\i49/n194 ),
    .C(\i49/n196 ),
    .Y(\i49/n316 ));
 AO21x2_ASAP7_75t_SL \i49/i246  (.A1(\i49/n81 ),
    .A2(\i49/n3 ),
    .B(\i49/n218 ),
    .Y(\i49/n315 ));
 OAI21xp5_ASAP7_75t_SL \i49/i247  (.A1(\i49/n49 ),
    .A2(\i49/n82 ),
    .B(\i49/n258 ),
    .Y(\i49/n314 ));
 NOR2x1_ASAP7_75t_SL \i49/i248  (.A(\i49/n131 ),
    .B(\i49/n209 ),
    .Y(\i49/n312 ));
 OAI211xp5_ASAP7_75t_SL \i49/i249  (.A1(\i49/n71 ),
    .A2(\i49/n109 ),
    .B(\i49/n117 ),
    .C(\i49/n141 ),
    .Y(\i49/n311 ));
 NOR2x1_ASAP7_75t_SL \i49/i25  (.A(\i49/n410 ),
    .B(\i49/n488 ),
    .Y(\i49/n505 ));
 NOR2xp33_ASAP7_75t_SL \i49/i250  (.A(\i49/n140 ),
    .B(\i49/n213 ),
    .Y(\i49/n26 ));
 NOR2xp33_ASAP7_75t_SL \i49/i251  (.A(\i49/n143 ),
    .B(\i49/n276 ),
    .Y(\i49/n283 ));
 AOI222xp33_ASAP7_75t_SL \i49/i252  (.A1(\i49/n537 ),
    .A2(\i49/n66 ),
    .B1(\i49/n5 ),
    .B2(\i49/n48 ),
    .C1(\i49/n532 ),
    .C2(\i49/n63 ),
    .Y(\i49/n310 ));
 OAI221xp5_ASAP7_75t_SL \i49/i253  (.A1(\i49/n522 ),
    .A2(\i49/n54 ),
    .B1(\i49/n59 ),
    .B2(\i49/n50 ),
    .C(\i49/n126 ),
    .Y(\i49/n309 ));
 INVx1_ASAP7_75t_SL \i49/i254  (.A(\i49/n543 ),
    .Y(\i49/n281 ));
 INVx1_ASAP7_75t_SL \i49/i255  (.A(\i49/n278 ),
    .Y(\i49/n279 ));
 INVx1_ASAP7_75t_SL \i49/i256  (.A(\i49/n276 ),
    .Y(\i49/n277 ));
 INVxp67_ASAP7_75t_SL \i49/i257  (.A(\i49/n269 ),
    .Y(\i49/n270 ));
 INVx1_ASAP7_75t_SL \i49/i258  (.A(\i49/n267 ),
    .Y(\i49/n268 ));
 OAI21xp33_ASAP7_75t_SL \i49/i259  (.A1(\i49/n75 ),
    .A2(\i49/n62 ),
    .B(\i49/n187 ),
    .Y(\i49/n265 ));
 NOR2x1_ASAP7_75t_SL \i49/i26  (.A(\i49/n472 ),
    .B(\i49/n468 ),
    .Y(\i49/n504 ));
 NAND2xp5_ASAP7_75t_SL \i49/i260  (.A(\i49/n99 ),
    .B(\i49/n135 ),
    .Y(\i49/n264 ));
 OAI21xp5_ASAP7_75t_SL \i49/i261  (.A1(\i49/n58 ),
    .A2(\i49/n57 ),
    .B(\i49/n83 ),
    .Y(\i49/n263 ));
 NOR2xp33_ASAP7_75t_SL \i49/i262  (.A(\i49/n144 ),
    .B(\i49/n180 ),
    .Y(\i49/n262 ));
 NAND2xp33_ASAP7_75t_L \i49/i263  (.A(\i49/n177 ),
    .B(\i49/n104 ),
    .Y(\i49/n261 ));
 OAI21xp5_ASAP7_75t_SL \i49/i264  (.A1(\i49/n536 ),
    .A2(\i49/n61 ),
    .B(\i49/n53 ),
    .Y(\i49/n260 ));
 NOR2xp33_ASAP7_75t_SL \i49/i265  (.A(\i49/n20 ),
    .B(\i49/n124 ),
    .Y(\i49/n259 ));
 OAI21xp5_ASAP7_75t_SL \i49/i266  (.A1(\i49/n76 ),
    .A2(\i49/n533 ),
    .B(\i49/n66 ),
    .Y(\i49/n258 ));
 OAI21xp5_ASAP7_75t_SL \i49/i267  (.A1(\i49/n522 ),
    .A2(\i49/n86 ),
    .B(\i49/n568 ),
    .Y(\i49/n257 ));
 AOI22xp5_ASAP7_75t_SL \i49/i268  (.A1(\i49/n83 ),
    .A2(\i49/n61 ),
    .B1(\i49/n79 ),
    .B2(\i49/n532 ),
    .Y(\i49/n256 ));
 OAI21xp5_ASAP7_75t_SL \i49/i269  (.A1(\i49/n18 ),
    .A2(\i49/n73 ),
    .B(\i49/n138 ),
    .Y(\i49/n255 ));
 NAND3xp33_ASAP7_75t_SL \i49/i27  (.A(\i49/n452 ),
    .B(\i49/n581 ),
    .C(\i49/n449 ),
    .Y(\i49/n503 ));
 OAI21xp5_ASAP7_75t_SL \i49/i270  (.A1(\i49/n76 ),
    .A2(\i49/n57 ),
    .B(\i49/n69 ),
    .Y(\i49/n254 ));
 AOI22xp5_ASAP7_75t_R \i49/i271  (.A1(\i49/n48 ),
    .A2(\i49/n91 ),
    .B1(\i49/n51 ),
    .B2(\i49/n76 ),
    .Y(\i49/n253 ));
 OA21x2_ASAP7_75t_SL \i49/i272  (.A1(\i49/n67 ),
    .A2(\i49/n16 ),
    .B(\i49/n182 ),
    .Y(\i49/n282 ));
 AOI21xp33_ASAP7_75t_SL \i49/i273  (.A1(\i49/n70 ),
    .A2(\i49/n67 ),
    .B(\i49/n49 ),
    .Y(\i49/n252 ));
 OAI21xp5_ASAP7_75t_SL \i49/i274  (.A1(\i49/n79 ),
    .A2(\i49/n91 ),
    .B(\i49/n84 ),
    .Y(\i49/n251 ));
 OA21x2_ASAP7_75t_SL \i49/i275  (.A1(\i49/n5 ),
    .A2(\i49/n91 ),
    .B(\i49/n87 ),
    .Y(\i49/n250 ));
 AOI22xp33_ASAP7_75t_SL \i49/i276  (.A1(\i49/n91 ),
    .A2(\i49/n58 ),
    .B1(\i49/n68 ),
    .B2(\i49/n3 ),
    .Y(\i49/n249 ));
 OAI21xp5_ASAP7_75t_SL \i49/i277  (.A1(\i49/n69 ),
    .A2(\i49/n51 ),
    .B(\i49/n84 ),
    .Y(\i49/n248 ));
 OAI21xp5_ASAP7_75t_SL \i49/i278  (.A1(\i49/n76 ),
    .A2(\i49/n536 ),
    .B(\i49/n91 ),
    .Y(\i49/n247 ));
 AOI21xp33_ASAP7_75t_SL \i49/i279  (.A1(\i49/n64 ),
    .A2(\i49/n82 ),
    .B(\i49/n49 ),
    .Y(\i49/n246 ));
 NOR2xp33_ASAP7_75t_L \i49/i28  (.A(\i49/n477 ),
    .B(\i49/n439 ),
    .Y(\i49/n502 ));
 OAI21xp5_ASAP7_75t_SL \i49/i280  (.A1(\i49/n522 ),
    .A2(\i49/n73 ),
    .B(\i49/n23 ),
    .Y(\i49/n245 ));
 AOI22xp5_ASAP7_75t_SL \i49/i281  (.A1(\i49/n63 ),
    .A2(\i49/n552 ),
    .B1(\i49/n79 ),
    .B2(\i49/n61 ),
    .Y(\i49/n244 ));
 AOI21xp33_ASAP7_75t_SL \i49/i282  (.A1(\i49/n77 ),
    .A2(\i49/n49 ),
    .B(\i49/n71 ),
    .Y(\i49/n243 ));
 OAI21xp5_ASAP7_75t_SL \i49/i283  (.A1(\i49/n87 ),
    .A2(\i49/n76 ),
    .B(\i49/n53 ),
    .Y(\i49/n242 ));
 OAI21xp5_ASAP7_75t_SL \i49/i284  (.A1(\i49/n536 ),
    .A2(\i49/n552 ),
    .B(\i49/n79 ),
    .Y(\i49/n241 ));
 NAND2xp5_ASAP7_75t_SL \i49/i285  (.A(\i49/n84 ),
    .B(\i49/n167 ),
    .Y(\i49/n25 ));
 NAND2xp5_ASAP7_75t_L \i49/i286  (.A(\i49/n197 ),
    .B(\i49/n198 ),
    .Y(\i49/n240 ));
 OAI22xp5_ASAP7_75t_SL \i49/i287  (.A1(\i49/n62 ),
    .A2(\i49/n85 ),
    .B1(\i49/n92 ),
    .B2(\i49/n16 ),
    .Y(\i49/n280 ));
 OAI22xp5_ASAP7_75t_SL \i49/i288  (.A1(\i49/n92 ),
    .A2(\i49/n73 ),
    .B1(\i49/n534 ),
    .B2(\i49/n70 ),
    .Y(\i49/n278 ));
 OAI22xp5_ASAP7_75t_SL \i49/i289  (.A1(\i49/n90 ),
    .A2(\i49/n60 ),
    .B1(\i49/n522 ),
    .B2(\i49/n541 ),
    .Y(\i49/n276 ));
 NOR5xp2_ASAP7_75t_SL \i49/i29  (.A(\i49/n441 ),
    .B(\i49/n432 ),
    .C(\i49/n388 ),
    .D(\i49/n352 ),
    .E(\i49/n356 ),
    .Y(\i49/n501 ));
 AOI22xp5_ASAP7_75t_SL \i49/i290  (.A1(\i49/n68 ),
    .A2(\i49/n88 ),
    .B1(\i49/n5 ),
    .B2(\i49/n533 ),
    .Y(\i49/n275 ));
 AOI22xp5_ASAP7_75t_SL \i49/i291  (.A1(\i49/n68 ),
    .A2(\i49/n552 ),
    .B1(\i49/n93 ),
    .B2(\i49/n61 ),
    .Y(\i49/n274 ));
 OAI22xp5_ASAP7_75t_SL \i49/i292  (.A1(\i49/n71 ),
    .A2(\i49/n541 ),
    .B1(\i49/n73 ),
    .B2(\i49/n52 ),
    .Y(\i49/n273 ));
 OAI22xp33_ASAP7_75t_SL \i49/i293  (.A1(\i49/n92 ),
    .A2(\i49/n89 ),
    .B1(\i49/n50 ),
    .B2(\i49/n8 ),
    .Y(\i49/n272 ));
 NAND2xp5_ASAP7_75t_L \i49/i294  (.A(\i49/n19 ),
    .B(\i49/n163 ),
    .Y(\i49/n271 ));
 OAI22xp5_ASAP7_75t_SL \i49/i295  (.A1(\i49/n522 ),
    .A2(\i49/n89 ),
    .B1(\i49/n70 ),
    .B2(\i49/n86 ),
    .Y(\i49/n269 ));
 NOR2xp33_ASAP7_75t_L \i49/i296  (.A(\i49/n16 ),
    .B(\i49/n21 ),
    .Y(\i49/n267 ));
 NAND2xp33_ASAP7_75t_L \i49/i297  (.A(\i49/n117 ),
    .B(\i49/n141 ),
    .Y(\i49/n239 ));
 OAI21xp5_ASAP7_75t_SL \i49/i298  (.A1(\i49/n71 ),
    .A2(\i49/n60 ),
    .B(\i49/n116 ),
    .Y(\i49/n266 ));
 INVxp67_ASAP7_75t_SL \i49/i299  (.A(\i49/n235 ),
    .Y(\i49/n236 ));
 INVx2_ASAP7_75t_SL \i49/i3  (.A(\i49/n8 ),
    .Y(\i49/n3 ));
 NOR3xp33_ASAP7_75t_SL \i49/i30  (.A(\i49/n437 ),
    .B(\i49/n454 ),
    .C(\i49/n486 ),
    .Y(\i49/n500 ));
 INVxp67_ASAP7_75t_SL \i49/i300  (.A(\i49/n233 ),
    .Y(\i49/n234 ));
 INVx1_ASAP7_75t_SL \i49/i301  (.A(\i49/n564 ),
    .Y(\i49/n232 ));
 INVx1_ASAP7_75t_SL \i49/i302  (.A(\i49/n228 ),
    .Y(\i49/n229 ));
 INVxp67_ASAP7_75t_SL \i49/i303  (.A(\i49/n226 ),
    .Y(\i49/n227 ));
 INVxp67_ASAP7_75t_SL \i49/i304  (.A(\i49/n222 ),
    .Y(\i49/n223 ));
 INVxp67_ASAP7_75t_SL \i49/i305  (.A(\i49/n220 ),
    .Y(\i49/n221 ));
 OAI22xp33_ASAP7_75t_SL \i49/i306  (.A1(\i49/n52 ),
    .A2(\i49/n89 ),
    .B1(\i49/n59 ),
    .B2(\i49/n62 ),
    .Y(\i49/n216 ));
 OAI21xp5_ASAP7_75t_SL \i49/i307  (.A1(\i49/n17 ),
    .A2(\i49/n8 ),
    .B(\i49/n566 ),
    .Y(\i49/n215 ));
 AOI22xp5_ASAP7_75t_SL \i49/i308  (.A1(\i49/n81 ),
    .A2(\i49/n552 ),
    .B1(\i49/n53 ),
    .B2(\i49/n3 ),
    .Y(\i49/n214 ));
 OAI22xp5_ASAP7_75t_SL \i49/i309  (.A1(\i49/n89 ),
    .A2(\i49/n55 ),
    .B1(\i49/n52 ),
    .B2(\i49/n16 ),
    .Y(\i49/n213 ));
 NOR2x1_ASAP7_75t_SL \i49/i31  (.A(\i49/n483 ),
    .B(\i49/n442 ),
    .Y(\i49/n499 ));
 AOI21xp33_ASAP7_75t_SL \i49/i310  (.A1(\i49/n73 ),
    .A2(\i49/n541 ),
    .B(\i49/n80 ),
    .Y(\i49/n212 ));
 AOI22xp33_ASAP7_75t_SL \i49/i311  (.A1(\i49/n68 ),
    .A2(\i49/n76 ),
    .B1(\i49/n5 ),
    .B2(\i49/n58 ),
    .Y(\i49/n211 ));
 OAI22xp33_ASAP7_75t_SL \i49/i312  (.A1(\i49/n62 ),
    .A2(\i49/n49 ),
    .B1(\i49/n85 ),
    .B2(\i49/n64 ),
    .Y(\i49/n210 ));
 AOI22xp5_ASAP7_75t_SL \i49/i313  (.A1(\i49/n93 ),
    .A2(\i49/n84 ),
    .B1(\i49/n83 ),
    .B2(\i49/n57 ),
    .Y(\i49/n238 ));
 OAI22xp33_ASAP7_75t_SL \i49/i314  (.A1(\i49/n534 ),
    .A2(\i49/n62 ),
    .B1(\i49/n541 ),
    .B2(\i49/n82 ),
    .Y(\i49/n209 ));
 OAI22xp5_ASAP7_75t_SL \i49/i315  (.A1(\i49/n90 ),
    .A2(\i49/n8 ),
    .B1(\i49/n17 ),
    .B2(\i49/n85 ),
    .Y(\i49/n208 ));
 OAI22xp5_ASAP7_75t_SL \i49/i316  (.A1(\i49/n64 ),
    .A2(\i49/n8 ),
    .B1(\i49/n82 ),
    .B2(\i49/n77 ),
    .Y(\i49/n207 ));
 AOI22xp5_ASAP7_75t_SL \i49/i317  (.A1(\i49/n48 ),
    .A2(\i49/n51 ),
    .B1(\i49/n93 ),
    .B2(\i49/n76 ),
    .Y(\i49/n237 ));
 OAI22xp33_ASAP7_75t_SL \i49/i318  (.A1(\i49/n54 ),
    .A2(\i49/n62 ),
    .B1(\i49/n16 ),
    .B2(\i49/n55 ),
    .Y(\i49/n206 ));
 OAI22xp5_ASAP7_75t_SL \i49/i319  (.A1(\i49/n62 ),
    .A2(\i49/n89 ),
    .B1(\i49/n70 ),
    .B2(\i49/n16 ),
    .Y(\i49/n205 ));
 NAND2xp5_ASAP7_75t_SL \i49/i32  (.A(\i49/n440 ),
    .B(\i49/n460 ),
    .Y(\i49/n498 ));
 OAI21xp5_ASAP7_75t_SL \i49/i320  (.A1(\i49/n78 ),
    .A2(\i49/n59 ),
    .B(\i49/n134 ),
    .Y(\i49/n204 ));
 OAI21xp5_ASAP7_75t_SL \i49/i321  (.A1(\i49/n50 ),
    .A2(\i49/n60 ),
    .B(\i49/n125 ),
    .Y(\i49/n235 ));
 AOI22xp5_ASAP7_75t_SL \i49/i322  (.A1(\i49/n48 ),
    .A2(\i49/n69 ),
    .B1(\i49/n51 ),
    .B2(\i49/n57 ),
    .Y(\i49/n233 ));
 OA21x2_ASAP7_75t_SL \i49/i323  (.A1(\i49/n55 ),
    .A2(\i49/n59 ),
    .B(\i49/n526 ),
    .Y(\i49/n203 ));
 AOI22xp5_ASAP7_75t_SL \i49/i324  (.A1(\i49/n87 ),
    .A2(\i49/n93 ),
    .B1(\i49/n81 ),
    .B2(\i49/n532 ),
    .Y(\i49/n231 ));
 OAI22xp5_ASAP7_75t_SL \i49/i325  (.A1(\i49/n55 ),
    .A2(\i49/n541 ),
    .B1(\i49/n70 ),
    .B2(\i49/n59 ),
    .Y(\i49/n230 ));
 OAI22xp5_ASAP7_75t_SL \i49/i326  (.A1(\i49/n49 ),
    .A2(\i49/n17 ),
    .B1(\i49/n62 ),
    .B2(\i49/n74 ),
    .Y(\i49/n202 ));
 NAND2xp33_ASAP7_75t_SL \i49/i327  (.A(\i49/n199 ),
    .B(\i49/n200 ),
    .Y(\i49/n201 ));
 OAI22x1_ASAP7_75t_SL \i49/i328  (.A1(\i49/n18 ),
    .A2(\i49/n89 ),
    .B1(\i49/n52 ),
    .B2(\i49/n75 ),
    .Y(\i49/n228 ));
 AOI22xp5_ASAP7_75t_SL \i49/i329  (.A1(\i49/n53 ),
    .A2(\i49/n552 ),
    .B1(\i49/n51 ),
    .B2(\i49/n87 ),
    .Y(\i49/n226 ));
 NOR3x1_ASAP7_75t_SL \i49/i33  (.A(\i49/n29 ),
    .B(\i49/n456 ),
    .C(\i49/n380 ),
    .Y(\i49/n506 ));
 AO22x2_ASAP7_75t_SL \i49/i330  (.A1(\i49/n91 ),
    .A2(\i49/n88 ),
    .B1(\i49/n56 ),
    .B2(\i49/n533 ),
    .Y(\i49/n225 ));
 OAI21xp5_ASAP7_75t_SL \i49/i331  (.A1(\i49/n78 ),
    .A2(\i49/n54 ),
    .B(\i49/n527 ),
    .Y(\i49/n224 ));
 OAI22xp33_ASAP7_75t_SL \i49/i332  (.A1(\i49/n80 ),
    .A2(\i49/n49 ),
    .B1(\i49/n50 ),
    .B2(\i49/n541 ),
    .Y(\i49/n222 ));
 OAI22xp5_ASAP7_75t_SL \i49/i333  (.A1(\i49/n64 ),
    .A2(\i49/n54 ),
    .B1(\i49/n70 ),
    .B2(\i49/n541 ),
    .Y(\i49/n220 ));
 AOI22xp5_ASAP7_75t_SL \i49/i334  (.A1(\i49/n48 ),
    .A2(\i49/n53 ),
    .B1(\i49/n72 ),
    .B2(\i49/n533 ),
    .Y(\i49/n219 ));
 OAI22xp5_ASAP7_75t_SL \i49/i335  (.A1(\i49/n77 ),
    .A2(\i49/n62 ),
    .B1(\i49/n74 ),
    .B2(\i49/n67 ),
    .Y(\i49/n218 ));
 OAI22xp5_ASAP7_75t_SL \i49/i336  (.A1(\i49/n67 ),
    .A2(\i49/n541 ),
    .B1(\i49/n71 ),
    .B2(\i49/n85 ),
    .Y(\i49/n24 ));
 OAI22xp5_ASAP7_75t_SL \i49/i337  (.A1(\i49/n55 ),
    .A2(\i49/n54 ),
    .B1(\i49/n59 ),
    .B2(\i49/n52 ),
    .Y(\i49/n217 ));
 INVxp67_ASAP7_75t_SL \i49/i338  (.A(\i49/n194 ),
    .Y(\i49/n195 ));
 INVx1_ASAP7_75t_SL \i49/i339  (.A(\i49/n192 ),
    .Y(\i49/n193 ));
 NOR3xp33_ASAP7_75t_SL \i49/i34  (.A(\i49/n480 ),
    .B(\i49/n29 ),
    .C(\i49/n398 ),
    .Y(\i49/n496 ));
 INVxp67_ASAP7_75t_SL \i49/i340  (.A(\i49/n190 ),
    .Y(\i49/n191 ));
 INVxp67_ASAP7_75t_SL \i49/i341  (.A(\i49/n562 ),
    .Y(\i49/n189 ));
 INVxp67_ASAP7_75t_SL \i49/i342  (.A(\i49/n187 ),
    .Y(\i49/n188 ));
 INVxp67_ASAP7_75t_SL \i49/i343  (.A(\i49/n184 ),
    .Y(\i49/n185 ));
 INVxp67_ASAP7_75t_SL \i49/i344  (.A(\i49/n568 ),
    .Y(\i49/n179 ));
 INVxp67_ASAP7_75t_SL \i49/i345  (.A(\i49/n177 ),
    .Y(\i49/n178 ));
 INVxp67_ASAP7_75t_SL \i49/i346  (.A(\i49/n174 ),
    .Y(\i49/n175 ));
 INVxp67_ASAP7_75t_SL \i49/i347  (.A(\i49/n172 ),
    .Y(\i49/n173 ));
 INVxp67_ASAP7_75t_SL \i49/i348  (.A(\i49/n169 ),
    .Y(\i49/n170 ));
 INVxp67_ASAP7_75t_SL \i49/i349  (.A(\i49/n21 ),
    .Y(\i49/n168 ));
 NOR2xp67_ASAP7_75t_SL \i49/i35  (.A(\i49/n461 ),
    .B(\i49/n29 ),
    .Y(\i49/n495 ));
 INVx1_ASAP7_75t_SL \i49/i350  (.A(\i49/n167 ),
    .Y(\i49/n166 ));
 NAND2xp5_ASAP7_75t_SL \i49/i351  (.A(\i49/n69 ),
    .B(\i49/n84 ),
    .Y(\i49/n200 ));
 NAND2xp5_ASAP7_75t_SL \i49/i352  (.A(\i49/n83 ),
    .B(\i49/n533 ),
    .Y(\i49/n165 ));
 NAND2xp5_ASAP7_75t_SL \i49/i353  (.A(\i49/n82 ),
    .B(\i49/n80 ),
    .Y(\i49/n164 ));
 NAND2xp5_ASAP7_75t_SL \i49/i354  (.A(\i49/n51 ),
    .B(\i49/n88 ),
    .Y(\i49/n163 ));
 NAND2xp33_ASAP7_75t_SL \i49/i355  (.A(\i49/n64 ),
    .B(\i49/n522 ),
    .Y(\i49/n162 ));
 NAND2xp5_ASAP7_75t_SL \i49/i356  (.A(\i49/n61 ),
    .B(\i49/n63 ),
    .Y(\i49/n161 ));
 NAND2xp5_ASAP7_75t_SL \i49/i357  (.A(\i49/n61 ),
    .B(\i49/n66 ),
    .Y(\i49/n199 ));
 NAND2xp5_ASAP7_75t_SL \i49/i358  (.A(\i49/n63 ),
    .B(\i49/n536 ),
    .Y(\i49/n198 ));
 NAND2xp5_ASAP7_75t_SL \i49/i359  (.A(\i49/n66 ),
    .B(\i49/n84 ),
    .Y(\i49/n160 ));
 NOR3xp33_ASAP7_75t_SL \i49/i36  (.A(\i49/n438 ),
    .B(\i49/n433 ),
    .C(\i49/n2 ),
    .Y(\i49/n494 ));
 NAND2xp5_ASAP7_75t_SL \i49/i360  (.A(\i49/n3 ),
    .B(\i49/n63 ),
    .Y(\i49/n159 ));
 NAND2xp5_ASAP7_75t_SL \i49/i361  (.A(\i49/n70 ),
    .B(\i49/n17 ),
    .Y(\i49/n158 ));
 NAND2xp5_ASAP7_75t_SL \i49/i362  (.A(\i49/n83 ),
    .B(\i49/n87 ),
    .Y(\i49/n157 ));
 NAND2xp5_ASAP7_75t_SL \i49/i363  (.A(\i49/n69 ),
    .B(\i49/n3 ),
    .Y(\i49/n156 ));
 NAND2xp33_ASAP7_75t_SL \i49/i364  (.A(\i49/n532 ),
    .B(\i49/n72 ),
    .Y(\i49/n155 ));
 NAND2xp5_ASAP7_75t_SL \i49/i365  (.A(\i49/n66 ),
    .B(\i49/n532 ),
    .Y(\i49/n154 ));
 NAND2xp5_ASAP7_75t_SL \i49/i366  (.A(\i49/n48 ),
    .B(\i49/n56 ),
    .Y(\i49/n153 ));
 NAND2xp5_ASAP7_75t_SL \i49/i367  (.A(\i49/n56 ),
    .B(\i49/n536 ),
    .Y(\i49/n152 ));
 NAND2xp5_ASAP7_75t_SL \i49/i368  (.A(\i49/n69 ),
    .B(\i49/n87 ),
    .Y(\i49/n151 ));
 NAND2xp5_ASAP7_75t_SL \i49/i369  (.A(\i49/n48 ),
    .B(\i49/n79 ),
    .Y(\i49/n197 ));
 NAND4xp25_ASAP7_75t_SL \i49/i37  (.A(\i49/n420 ),
    .B(\i49/n414 ),
    .C(\i49/n413 ),
    .D(\i49/n447 ),
    .Y(\i49/n493 ));
 AND2x2_ASAP7_75t_SL \i49/i370  (.A(\i49/n56 ),
    .B(\i49/n76 ),
    .Y(\i49/n196 ));
 AND2x2_ASAP7_75t_SL \i49/i371  (.A(\i49/n83 ),
    .B(\i49/n536 ),
    .Y(\i49/n194 ));
 AND2x2_ASAP7_75t_SL \i49/i372  (.A(\i49/n93 ),
    .B(\i49/n532 ),
    .Y(\i49/n192 ));
 NAND2xp5_ASAP7_75t_SL \i49/i373  (.A(\i49/n532 ),
    .B(\i49/n5 ),
    .Y(\i49/n23 ));
 NAND2xp5_ASAP7_75t_SL \i49/i374  (.A(\i49/n79 ),
    .B(\i49/n87 ),
    .Y(\i49/n190 ));
 NAND2xp5_ASAP7_75t_SL \i49/i375  (.A(\i49/n65 ),
    .B(\i49/n536 ),
    .Y(\i49/n187 ));
 AND2x2_ASAP7_75t_SL \i49/i376  (.A(\i49/n69 ),
    .B(\i49/n552 ),
    .Y(\i49/n186 ));
 NOR2xp67_ASAP7_75t_SL \i49/i377  (.A(\i49/n67 ),
    .B(\i49/n73 ),
    .Y(\i49/n22 ));
 NOR2xp33_ASAP7_75t_SL \i49/i378  (.A(\i49/n59 ),
    .B(\i49/n67 ),
    .Y(\i49/n184 ));
 NAND2xp5_ASAP7_75t_SL \i49/i379  (.A(\i49/n68 ),
    .B(\i49/n3 ),
    .Y(\i49/n150 ));
 NAND3xp33_ASAP7_75t_L \i49/i38  (.A(\i49/n396 ),
    .B(\i49/n414 ),
    .C(\i49/n465 ),
    .Y(\i49/n492 ));
 NAND2xp5_ASAP7_75t_SL \i49/i380  (.A(\i49/n537 ),
    .B(\i49/n68 ),
    .Y(\i49/n183 ));
 NAND2xp5_ASAP7_75t_SL \i49/i381  (.A(\i49/n65 ),
    .B(\i49/n61 ),
    .Y(\i49/n182 ));
 NAND2xp5_ASAP7_75t_SL \i49/i382  (.A(\i49/n552 ),
    .B(\i49/n63 ),
    .Y(\i49/n149 ));
 NOR2xp33_ASAP7_75t_SL \i49/i383  (.A(\i49/n62 ),
    .B(\i49/n541 ),
    .Y(\i49/n181 ));
 AND2x2_ASAP7_75t_SL \i49/i384  (.A(\i49/n66 ),
    .B(\i49/n3 ),
    .Y(\i49/n180 ));
 NOR2xp33_ASAP7_75t_SL \i49/i385  (.A(\i49/n18 ),
    .B(\i49/n16 ),
    .Y(\i49/n148 ));
 NOR2xp33_ASAP7_75t_SL \i49/i386  (.A(\i49/n65 ),
    .B(\i49/n83 ),
    .Y(\i49/n147 ));
 NOR2xp33_ASAP7_75t_SL \i49/i387  (.A(\i49/n62 ),
    .B(\i49/n86 ),
    .Y(\i49/n146 ));
 NAND2xp5_ASAP7_75t_SL \i49/i388  (.A(\i49/n83 ),
    .B(\i49/n3 ),
    .Y(\i49/n177 ));
 NOR2xp33_ASAP7_75t_L \i49/i389  (.A(\i49/n91 ),
    .B(\i49/n53 ),
    .Y(\i49/n176 ));
 NAND3xp33_ASAP7_75t_SL \i49/i39  (.A(\i49/n400 ),
    .B(\i49/n448 ),
    .C(\i49/n434 ),
    .Y(\i49/n491 ));
 NAND2xp5_ASAP7_75t_SL \i49/i390  (.A(\i49/n91 ),
    .B(\i49/n57 ),
    .Y(\i49/n174 ));
 NAND2xp5_ASAP7_75t_SL \i49/i391  (.A(\i49/n87 ),
    .B(\i49/n66 ),
    .Y(\i49/n172 ));
 NAND2xp5_ASAP7_75t_SL \i49/i392  (.A(\i49/n91 ),
    .B(\i49/n532 ),
    .Y(\i49/n171 ));
 NAND2xp5_ASAP7_75t_SL \i49/i393  (.A(\i49/n69 ),
    .B(\i49/n537 ),
    .Y(\i49/n145 ));
 NOR2xp67_ASAP7_75t_SL \i49/i394  (.A(\i49/n83 ),
    .B(\i49/n69 ),
    .Y(\i49/n169 ));
 NOR2xp33_ASAP7_75t_SL \i49/i395  (.A(\i49/n60 ),
    .B(\i49/n82 ),
    .Y(\i49/n144 ));
 NOR2x1_ASAP7_75t_SL \i49/i396  (.A(\i49/n65 ),
    .B(\i49/n81 ),
    .Y(\i49/n21 ));
 OR2x2_ASAP7_75t_SL \i49/i397  (.A(\i49/n53 ),
    .B(\i49/n68 ),
    .Y(\i49/n167 ));
 INVxp67_ASAP7_75t_SL \i49/i398  (.A(\i49/n142 ),
    .Y(\i49/n143 ));
 INVxp67_ASAP7_75t_SL \i49/i399  (.A(\i49/n138 ),
    .Y(\i49/n139 ));
 INVx1_ASAP7_75t_SL \i49/i4  (.A(\i49/n35 ),
    .Y(\i49/n4 ));
 NAND2xp5_ASAP7_75t_L \i49/i40  (.A(\i49/n574 ),
    .B(\i49/n481 ),
    .Y(\i49/n490 ));
 INVx1_ASAP7_75t_SL \i49/i400  (.A(\i49/n136 ),
    .Y(\i49/n137 ));
 INVxp67_ASAP7_75t_SL \i49/i401  (.A(\i49/n132 ),
    .Y(\i49/n133 ));
 INVxp67_ASAP7_75t_SL \i49/i402  (.A(\i49/n565 ),
    .Y(\i49/n131 ));
 INVxp67_ASAP7_75t_SL \i49/i403  (.A(\i49/n129 ),
    .Y(\i49/n130 ));
 INVxp67_ASAP7_75t_SL \i49/i404  (.A(\i49/n566 ),
    .Y(\i49/n128 ));
 INVxp67_ASAP7_75t_SL \i49/i405  (.A(\i49/n126 ),
    .Y(\i49/n127 ));
 INVxp67_ASAP7_75t_SL \i49/i406  (.A(\i49/n124 ),
    .Y(\i49/n125 ));
 INVxp67_ASAP7_75t_SL \i49/i407  (.A(\i49/n529 ),
    .Y(\i49/n118 ));
 INVx1_ASAP7_75t_SL \i49/i408  (.A(\i49/n530 ),
    .Y(\i49/n115 ));
 INVx1_ASAP7_75t_SL \i49/i409  (.A(\i49/n19 ),
    .Y(\i49/n20 ));
 NAND2xp33_ASAP7_75t_SL \i49/i41  (.A(\i49/n445 ),
    .B(\i49/n463 ),
    .Y(\i49/n489 ));
 NAND2xp5_ASAP7_75t_SL \i49/i410  (.A(\i49/n81 ),
    .B(\i49/n76 ),
    .Y(\i49/n114 ));
 NAND2xp5_ASAP7_75t_SL \i49/i411  (.A(\i49/n53 ),
    .B(\i49/n537 ),
    .Y(\i49/n113 ));
 NAND2xp5_ASAP7_75t_SL \i49/i412  (.A(\i49/n78 ),
    .B(\i49/n71 ),
    .Y(\i49/n112 ));
 NAND2xp5_ASAP7_75t_SL \i49/i413  (.A(\i49/n537 ),
    .B(\i49/n51 ),
    .Y(\i49/n111 ));
 NAND2xp5_ASAP7_75t_SL \i49/i414  (.A(\i49/n79 ),
    .B(\i49/n552 ),
    .Y(\i49/n110 ));
 NOR2xp33_ASAP7_75t_SL \i49/i415  (.A(\i49/n87 ),
    .B(\i49/n3 ),
    .Y(\i49/n109 ));
 NAND2xp5_ASAP7_75t_SL \i49/i416  (.A(\i49/n72 ),
    .B(\i49/n57 ),
    .Y(\i49/n108 ));
 NAND2xp5_ASAP7_75t_SL \i49/i417  (.A(\i49/n51 ),
    .B(\i49/n536 ),
    .Y(\i49/n107 ));
 NAND2xp5_ASAP7_75t_L \i49/i418  (.A(\i49/n534 ),
    .B(\i49/n49 ),
    .Y(\i49/n106 ));
 NAND2xp5_ASAP7_75t_SL \i49/i419  (.A(\i49/n5 ),
    .B(\i49/n61 ),
    .Y(\i49/n105 ));
 NOR2x1_ASAP7_75t_SL \i49/i42  (.A(\i49/n462 ),
    .B(\i49/n471 ),
    .Y(\i49/n497 ));
 NAND2xp5_ASAP7_75t_SL \i49/i420  (.A(\i49/n93 ),
    .B(\i49/n58 ),
    .Y(\i49/n142 ));
 NAND2xp5_ASAP7_75t_SL \i49/i421  (.A(\i49/n81 ),
    .B(\i49/n61 ),
    .Y(\i49/n104 ));
 NOR2xp33_ASAP7_75t_SL \i49/i422  (.A(\i49/n60 ),
    .B(\i49/n522 ),
    .Y(\i49/n103 ));
 NAND2xp5_ASAP7_75t_SL \i49/i423  (.A(\i49/n3 ),
    .B(\i49/n93 ),
    .Y(\i49/n141 ));
 AND2x2_ASAP7_75t_SL \i49/i424  (.A(\i49/n5 ),
    .B(\i49/n537 ),
    .Y(\i49/n140 ));
 NAND2xp5_ASAP7_75t_SL \i49/i425  (.A(\i49/n83 ),
    .B(\i49/n552 ),
    .Y(\i49/n138 ));
 NOR2x1_ASAP7_75t_SL \i49/i426  (.A(\i49/n536 ),
    .B(\i49/n533 ),
    .Y(\i49/n136 ));
 NAND2xp5_ASAP7_75t_SL \i49/i427  (.A(\i49/n79 ),
    .B(\i49/n57 ),
    .Y(\i49/n135 ));
 NAND2xp5_ASAP7_75t_SL \i49/i428  (.A(\i49/n51 ),
    .B(\i49/n76 ),
    .Y(\i49/n102 ));
 NAND2xp5_ASAP7_75t_SL \i49/i429  (.A(\i49/n56 ),
    .B(\i49/n61 ),
    .Y(\i49/n134 ));
 NAND2xp33_ASAP7_75t_L \i49/i43  (.A(\i49/n451 ),
    .B(\i49/n422 ),
    .Y(\i49/n486 ));
 NOR2xp33_ASAP7_75t_SL \i49/i430  (.A(\i49/n536 ),
    .B(\i49/n61 ),
    .Y(\i49/n101 ));
 NAND2xp5_ASAP7_75t_SL \i49/i431  (.A(\i49/n81 ),
    .B(\i49/n87 ),
    .Y(\i49/n132 ));
 NOR2xp67_ASAP7_75t_SL \i49/i432  (.A(\i49/n55 ),
    .B(\i49/n85 ),
    .Y(\i49/n129 ));
 NAND2xp33_ASAP7_75t_L \i49/i433  (.A(\i49/n54 ),
    .B(\i49/n75 ),
    .Y(\i49/n100 ));
 NAND2xp5_ASAP7_75t_SL \i49/i434  (.A(\i49/n48 ),
    .B(\i49/n93 ),
    .Y(\i49/n126 ));
 NOR2xp33_ASAP7_75t_SL \i49/i435  (.A(\i49/n49 ),
    .B(\i49/n522 ),
    .Y(\i49/n124 ));
 NAND2xp5_ASAP7_75t_SL \i49/i436  (.A(\i49/n53 ),
    .B(\i49/n533 ),
    .Y(\i49/n123 ));
 AND2x2_ASAP7_75t_SL \i49/i437  (.A(\i49/n93 ),
    .B(\i49/n533 ),
    .Y(\i49/n122 ));
 NAND2xp5_ASAP7_75t_L \i49/i438  (.A(\i49/n16 ),
    .B(\i49/n534 ),
    .Y(\i49/n121 ));
 NAND2xp33_ASAP7_75t_L \i49/i439  (.A(\i49/n3 ),
    .B(\i49/n79 ),
    .Y(\i49/n99 ));
 NAND2xp33_ASAP7_75t_L \i49/i44  (.A(\i49/n574 ),
    .B(\i49/n428 ),
    .Y(\i49/n485 ));
 AND2x2_ASAP7_75t_SL \i49/i440  (.A(\i49/n93 ),
    .B(\i49/n552 ),
    .Y(\i49/n120 ));
 NOR2xp33_ASAP7_75t_SL \i49/i441  (.A(\i49/n59 ),
    .B(\i49/n52 ),
    .Y(\i49/n98 ));
 NOR2xp33_ASAP7_75t_SL \i49/i442  (.A(\i49/n58 ),
    .B(\i49/n76 ),
    .Y(\i49/n119 ));
 NAND2xp5_ASAP7_75t_SL \i49/i443  (.A(\i49/n5 ),
    .B(\i49/n533 ),
    .Y(\i49/n97 ));
 NAND2xp5_ASAP7_75t_SL \i49/i444  (.A(\i49/n51 ),
    .B(\i49/n3 ),
    .Y(\i49/n96 ));
 NAND2xp5_ASAP7_75t_SL \i49/i445  (.A(\i49/n79 ),
    .B(\i49/n533 ),
    .Y(\i49/n117 ));
 NAND2xp5_ASAP7_75t_SL \i49/i446  (.A(\i49/n93 ),
    .B(\i49/n537 ),
    .Y(\i49/n116 ));
 NOR2xp33_ASAP7_75t_SL \i49/i447  (.A(\i49/n92 ),
    .B(\i49/n16 ),
    .Y(\i49/n95 ));
 NOR2xp33_ASAP7_75t_SL \i49/i448  (.A(\i49/n92 ),
    .B(\i49/n60 ),
    .Y(\i49/n94 ));
 NAND2xp5_ASAP7_75t_SL \i49/i449  (.A(\i49/n5 ),
    .B(\i49/n57 ),
    .Y(\i49/n19 ));
 NOR2xp33_ASAP7_75t_SL \i49/i45  (.A(\i49/n427 ),
    .B(\i49/n453 ),
    .Y(\i49/n484 ));
 INVx2_ASAP7_75t_SL \i49/i450  (.A(\i49/n93 ),
    .Y(\i49/n92 ));
 INVx1_ASAP7_75t_SL \i49/i451  (.A(\i49/n91 ),
    .Y(\i49/n90 ));
 INVx3_ASAP7_75t_SL \i49/i452  (.A(\i49/n89 ),
    .Y(\i49/n88 ));
 INVx2_ASAP7_75t_SL \i49/i453  (.A(\i49/n87 ),
    .Y(\i49/n86 ));
 INVx4_ASAP7_75t_SL \i49/i454  (.A(\i49/n85 ),
    .Y(\i49/n84 ));
 INVx3_ASAP7_75t_SL \i49/i455  (.A(\i49/n83 ),
    .Y(\i49/n82 ));
 INVx2_ASAP7_75t_SL \i49/i456  (.A(\i49/n81 ),
    .Y(\i49/n80 ));
 INVx2_ASAP7_75t_SL \i49/i457  (.A(\i49/n79 ),
    .Y(\i49/n78 ));
 INVx3_ASAP7_75t_SL \i49/i458  (.A(\i49/n537 ),
    .Y(\i49/n77 ));
 INVx2_ASAP7_75t_SL \i49/i459  (.A(\i49/n76 ),
    .Y(\i49/n75 ));
 NAND3xp33_ASAP7_75t_SL \i49/i46  (.A(\i49/n417 ),
    .B(\i49/n425 ),
    .C(\i49/n391 ),
    .Y(\i49/n483 ));
 INVx2_ASAP7_75t_SL \i49/i460  (.A(\i49/n532 ),
    .Y(\i49/n74 ));
 INVx3_ASAP7_75t_SL \i49/i461  (.A(\i49/n536 ),
    .Y(\i49/n73 ));
 INVx3_ASAP7_75t_SL \i49/i462  (.A(\i49/n72 ),
    .Y(\i49/n71 ));
 INVx3_ASAP7_75t_SL \i49/i463  (.A(\i49/n70 ),
    .Y(\i49/n69 ));
 AND2x4_ASAP7_75t_SL \i49/i464  (.A(\i49/n40 ),
    .B(\i49/n44 ),
    .Y(\i49/n93 ));
 AND2x4_ASAP7_75t_SL \i49/i465  (.A(\i49/n42 ),
    .B(\i49/n40 ),
    .Y(\i49/n91 ));
 OR2x2_ASAP7_75t_SL \i49/i466  (.A(\i49/n6 ),
    .B(\i49/n34 ),
    .Y(\i49/n89 ));
 AND2x4_ASAP7_75t_SL \i49/i467  (.A(\i49/n4 ),
    .B(\i49/n549 ),
    .Y(\i49/n87 ));
 OR2x6_ASAP7_75t_SL \i49/i468  (.A(\i49/n37 ),
    .B(\i49/n47 ),
    .Y(\i49/n85 ));
 AND2x4_ASAP7_75t_SL \i49/i469  (.A(\i49/n33 ),
    .B(\i49/n46 ),
    .Y(\i49/n83 ));
 NOR2x1_ASAP7_75t_SL \i49/i47  (.A(\i49/n373 ),
    .B(\i49/n436 ),
    .Y(\i49/n482 ));
 AND2x4_ASAP7_75t_SL \i49/i470  (.A(\i49/n33 ),
    .B(\i49/n42 ),
    .Y(\i49/n81 ));
 AND2x4_ASAP7_75t_SL \i49/i471  (.A(\i49/n33 ),
    .B(\i49/n519 ),
    .Y(\i49/n79 ));
 AND2x4_ASAP7_75t_SL \i49/i472  (.A(\i49/n549 ),
    .B(\i49/n15 ),
    .Y(\i49/n76 ));
 AND2x4_ASAP7_75t_SL \i49/i473  (.A(\i49/n42 ),
    .B(\i49/n41 ),
    .Y(\i49/n72 ));
 OR2x6_ASAP7_75t_SL \i49/i474  (.A(\i49/n43 ),
    .B(\i49/n32 ),
    .Y(\i49/n70 ));
 INVx3_ASAP7_75t_SL \i49/i475  (.A(\i49/n68 ),
    .Y(\i49/n67 ));
 INVx3_ASAP7_75t_SL \i49/i476  (.A(\i49/n66 ),
    .Y(\i49/n18 ));
 INVx3_ASAP7_75t_SL \i49/i477  (.A(\i49/n65 ),
    .Y(\i49/n64 ));
 INVx3_ASAP7_75t_SL \i49/i478  (.A(\i49/n63 ),
    .Y(\i49/n62 ));
 INVx2_ASAP7_75t_SL \i49/i479  (.A(\i49/n61 ),
    .Y(\i49/n60 ));
 NOR2xp33_ASAP7_75t_SL \i49/i48  (.A(\i49/n443 ),
    .B(\i49/n352 ),
    .Y(\i49/n481 ));
 INVx4_ASAP7_75t_SL \i49/i480  (.A(\i49/n59 ),
    .Y(\i49/n58 ));
 INVx4_ASAP7_75t_SL \i49/i481  (.A(\i49/n57 ),
    .Y(\i49/n16 ));
 INVx4_ASAP7_75t_SL \i49/i482  (.A(\i49/n56 ),
    .Y(\i49/n55 ));
 INVx3_ASAP7_75t_SL \i49/i483  (.A(\i49/n53 ),
    .Y(\i49/n52 ));
 INVx3_ASAP7_75t_SL \i49/i484  (.A(\i49/n51 ),
    .Y(\i49/n50 ));
 INVx3_ASAP7_75t_SL \i49/i485  (.A(\i49/n49 ),
    .Y(\i49/n48 ));
 AND2x4_ASAP7_75t_SL \i49/i486  (.A(\i49/n42 ),
    .B(\i49/n520 ),
    .Y(\i49/n68 ));
 AND2x4_ASAP7_75t_SL \i49/i487  (.A(\i49/n40 ),
    .B(\i49/n46 ),
    .Y(\i49/n66 ));
 AND2x4_ASAP7_75t_SL \i49/i488  (.A(\i49/n44 ),
    .B(\i49/n41 ),
    .Y(\i49/n65 ));
 OR2x2_ASAP7_75t_SL \i49/i489  (.A(\i49/n10 ),
    .B(\i49/n45 ),
    .Y(\i49/n17 ));
 NAND2xp5_ASAP7_75t_SL \i49/i49  (.A(\i49/n451 ),
    .B(\i49/n446 ),
    .Y(\i49/n480 ));
 AND2x4_ASAP7_75t_SL \i49/i490  (.A(\i49/n519 ),
    .B(\i49/n40 ),
    .Y(\i49/n63 ));
 NAND2x1p5_ASAP7_75t_SL \i49/i491  (.A(\i49/n4 ),
    .B(\i49/n38 ),
    .Y(\i49/n8 ));
 AND2x4_ASAP7_75t_SL \i49/i492  (.A(\i49/n38 ),
    .B(\i49/n15 ),
    .Y(\i49/n61 ));
 OR2x4_ASAP7_75t_SL \i49/i493  (.A(\i49/n35 ),
    .B(\i49/n36 ),
    .Y(\i49/n59 ));
 AND2x4_ASAP7_75t_SL \i49/i494  (.A(\i49/n538 ),
    .B(\i49/n15 ),
    .Y(\i49/n57 ));
 AND2x4_ASAP7_75t_SL \i49/i495  (.A(\i49/n44 ),
    .B(\i49/n520 ),
    .Y(\i49/n56 ));
 NAND2x1_ASAP7_75t_SL \i49/i496  (.A(\i49/n4 ),
    .B(\i49/n557 ),
    .Y(\i49/n54 ));
 AND2x4_ASAP7_75t_SL \i49/i497  (.A(\i49/n519 ),
    .B(\i49/n41 ),
    .Y(\i49/n53 ));
 AND2x4_ASAP7_75t_SL \i49/i498  (.A(\i49/n46 ),
    .B(\i49/n41 ),
    .Y(\i49/n51 ));
 OR2x6_ASAP7_75t_SL \i49/i499  (.A(\i49/n31 ),
    .B(\i49/n39 ),
    .Y(\i49/n49 ));
 INVx2_ASAP7_75t_SL \i49/i5  (.A(\i49/n17 ),
    .Y(\i49/n5 ));
 NOR2xp33_ASAP7_75t_SL \i49/i50  (.A(\i49/n356 ),
    .B(\i49/n453 ),
    .Y(\i49/n479 ));
 INVx2_ASAP7_75t_SL \i49/i500  (.A(\i49/n550 ),
    .Y(\i49/n47 ));
 INVx2_ASAP7_75t_SL \i49/i501  (.A(\i49/n45 ),
    .Y(\i49/n46 ));
 INVx3_ASAP7_75t_SL \i49/i502  (.A(\i49/n43 ),
    .Y(\i49/n44 ));
 NAND2xp5_ASAP7_75t_SL \i49/i503  (.A(\i49/n11 ),
    .B(\i49/n0 ),
    .Y(\i49/n39 ));
 NAND2xp5_ASAP7_75t_SL \i49/i504  (.A(\i49/n9 ),
    .B(n23[5]),
    .Y(\i49/n45 ));
 NAND2x1p5_ASAP7_75t_SL \i49/i505  (.A(n23[4]),
    .B(n23[5]),
    .Y(\i49/n43 ));
 AND2x2_ASAP7_75t_SL \i49/i506  (.A(\i49/n571 ),
    .B(\i49/n9 ),
    .Y(\i49/n42 ));
 AND2x4_ASAP7_75t_SL \i49/i507  (.A(n23[7]),
    .B(\i49/n14 ),
    .Y(\i49/n41 ));
 AND2x2_ASAP7_75t_SL \i49/i508  (.A(\i49/n12 ),
    .B(\i49/n14 ),
    .Y(\i49/n40 ));
 INVx1_ASAP7_75t_SL \i49/i509  (.A(\i49/n38 ),
    .Y(\i49/n37 ));
 NOR2x1_ASAP7_75t_SL \i49/i51  (.A(\i49/n426 ),
    .B(\i49/n437 ),
    .Y(\i49/n478 ));
 INVx2_ASAP7_75t_SL \i49/i510  (.A(\i49/n33 ),
    .Y(\i49/n32 ));
 NAND2xp5_ASAP7_75t_SL \i49/i511  (.A(\i49/n30 ),
    .B(\i49/n1 ),
    .Y(\i49/n31 ));
 AND2x4_ASAP7_75t_SL \i49/i512  (.A(n23[0]),
    .B(\i49/n30 ),
    .Y(\i49/n38 ));
 NAND2xp5_ASAP7_75t_SL \i49/i513  (.A(\i49/n1 ),
    .B(n23[1]),
    .Y(\i49/n36 ));
 OR2x2_ASAP7_75t_SL \i49/i514  (.A(\i49/n0 ),
    .B(n23[3]),
    .Y(\i49/n35 ));
 NAND2x1_ASAP7_75t_SL \i49/i515  (.A(n23[3]),
    .B(\i49/n0 ),
    .Y(\i49/n34 ));
 AND2x2_ASAP7_75t_SL \i49/i516  (.A(n23[7]),
    .B(n23[6]),
    .Y(\i49/n33 ));
 INVx1_ASAP7_75t_SL \i49/i517  (.A(n23[1]),
    .Y(\i49/n30 ));
 INVx2_ASAP7_75t_SL \i49/i518  (.A(\i49/n34 ),
    .Y(\i49/n15 ));
 INVx2_ASAP7_75t_SL \i49/i519  (.A(n23[6]),
    .Y(\i49/n14 ));
 NAND2xp5_ASAP7_75t_SL \i49/i52  (.A(\i49/n390 ),
    .B(\i49/n431 ),
    .Y(\i49/n477 ));
 INVx2_ASAP7_75t_SL \i49/i520  (.A(n23[7]),
    .Y(\i49/n12 ));
 INVx2_ASAP7_75t_SL \i49/i521  (.A(n23[3]),
    .Y(\i49/n11 ));
 NAND2xp5_ASAP7_75t_SL \i49/i522  (.A(\i49/n12 ),
    .B(n23[6]),
    .Y(\i49/n10 ));
 INVx2_ASAP7_75t_SL \i49/i523  (.A(n23[4]),
    .Y(\i49/n9 ));
 OR2x2_ASAP7_75t_SL \i49/i524  (.A(\i49/n569 ),
    .B(\i49/n230 ),
    .Y(\i49/n7 ));
 OR2x2_ASAP7_75t_SL \i49/i525  (.A(n23[0]),
    .B(n23[1]),
    .Y(\i49/n6 ));
 INVx2_ASAP7_75t_SL \i49/i526  (.A(\i49/n349 ),
    .Y(\i49/n518 ));
 AND2x2_ASAP7_75t_SL \i49/i527  (.A(n23[4]),
    .B(\i49/n571 ),
    .Y(\i49/n519 ));
 AND2x2_ASAP7_75t_L \i49/i528  (.A(\i49/n12 ),
    .B(n23[6]),
    .Y(\i49/n520 ));
 INVx4_ASAP7_75t_SL \i49/i529  (.A(\i49/n521 ),
    .Y(\i49/n522 ));
 NOR5xp2_ASAP7_75t_SL \i49/i53  (.A(\i49/n311 ),
    .B(\i49/n27 ),
    .C(\i49/n324 ),
    .D(\i49/n28 ),
    .E(\i49/n288 ),
    .Y(\i49/n476 ));
 AND2x4_ASAP7_75t_SL \i49/i530  (.A(\i49/n519 ),
    .B(\i49/n520 ),
    .Y(\i49/n521 ));
 OAI21xp5_ASAP7_75t_SL \i49/i531  (.A1(\i49/n521 ),
    .A2(\i49/n72 ),
    .B(\i49/n536 ),
    .Y(\i49/n523 ));
 OAI21xp5_ASAP7_75t_SL \i49/i532  (.A1(\i49/n81 ),
    .A2(\i49/n521 ),
    .B(\i49/n58 ),
    .Y(\i49/n524 ));
 AOI22xp5_ASAP7_75t_SL \i49/i533  (.A1(\i49/n521 ),
    .A2(\i49/n533 ),
    .B1(\i49/n51 ),
    .B2(\i49/n552 ),
    .Y(\i49/n525 ));
 NAND2xp5_ASAP7_75t_SL \i49/i534  (.A(\i49/n521 ),
    .B(\i49/n76 ),
    .Y(\i49/n526 ));
 NAND2xp5_ASAP7_75t_SL \i49/i535  (.A(\i49/n521 ),
    .B(\i49/n537 ),
    .Y(\i49/n527 ));
 NAND2xp5_ASAP7_75t_SL \i49/i536  (.A(\i49/n3 ),
    .B(\i49/n521 ),
    .Y(\i49/n528 ));
 NAND2xp5_ASAP7_75t_SL \i49/i537  (.A(\i49/n521 ),
    .B(\i49/n57 ),
    .Y(\i49/n529 ));
 NAND2xp5_ASAP7_75t_SL \i49/i538  (.A(\i49/n521 ),
    .B(\i49/n84 ),
    .Y(\i49/n530 ));
 AND2x4_ASAP7_75t_SL \i49/i539  (.A(\i49/n549 ),
    .B(\i49/n531 ),
    .Y(\i49/n532 ));
 NOR2x1_ASAP7_75t_SL \i49/i54  (.A(\i49/n2 ),
    .B(\i49/n438 ),
    .Y(\i49/n475 ));
 AND2x4_ASAP7_75t_SL \i49/i540  (.A(n23[2]),
    .B(n23[3]),
    .Y(\i49/n531 ));
 AND2x4_ASAP7_75t_SL \i49/i541  (.A(\i49/n531 ),
    .B(\i49/n557 ),
    .Y(\i49/n533 ));
 NAND2x1_ASAP7_75t_SL \i49/i542  (.A(\i49/n531 ),
    .B(\i49/n557 ),
    .Y(\i49/n534 ));
 AND2x4_ASAP7_75t_SL \i49/i543  (.A(\i49/n535 ),
    .B(\i49/n538 ),
    .Y(\i49/n536 ));
 AND2x2_ASAP7_75t_SL \i49/i544  (.A(n23[2]),
    .B(n23[3]),
    .Y(\i49/n535 ));
 AND2x4_ASAP7_75t_SL \i49/i545  (.A(\i49/n535 ),
    .B(\i49/n38 ),
    .Y(\i49/n537 ));
 INVx2_ASAP7_75t_SL \i49/i546  (.A(\i49/n36 ),
    .Y(\i49/n538 ));
 NAND2xp5_ASAP7_75t_SL \i49/i547  (.A(\i49/n521 ),
    .B(\i49/n539 ),
    .Y(\i49/n540 ));
 AND2x4_ASAP7_75t_SL \i49/i548  (.A(\i49/n550 ),
    .B(\i49/n538 ),
    .Y(\i49/n539 ));
 INVx4_ASAP7_75t_SL \i49/i549  (.A(\i49/n539 ),
    .Y(\i49/n541 ));
 NAND2xp5_ASAP7_75t_SL \i49/i55  (.A(\i49/n435 ),
    .B(\i49/n415 ),
    .Y(\i49/n488 ));
 OAI21xp5_ASAP7_75t_SL \i49/i550  (.A1(\i49/n61 ),
    .A2(\i49/n539 ),
    .B(\i49/n79 ),
    .Y(\i49/n542 ));
 AOI22xp5_ASAP7_75t_SL \i49/i551  (.A1(\i49/n93 ),
    .A2(\i49/n539 ),
    .B1(\i49/n79 ),
    .B2(\i49/n3 ),
    .Y(\i49/n543 ));
 AOI22xp5_ASAP7_75t_SL \i49/i552  (.A1(\i49/n66 ),
    .A2(\i49/n539 ),
    .B1(\i49/n51 ),
    .B2(\i49/n533 ),
    .Y(\i49/n544 ));
 NAND2xp5_ASAP7_75t_SL \i49/i553  (.A(\i49/n65 ),
    .B(\i49/n539 ),
    .Y(\i49/n545 ));
 NOR2xp33_ASAP7_75t_SL \i49/i554  (.A(\i49/n87 ),
    .B(\i49/n539 ),
    .Y(\i49/n546 ));
 NAND2xp5_ASAP7_75t_SL \i49/i555  (.A(\i49/n5 ),
    .B(\i49/n539 ),
    .Y(\i49/n547 ));
 NAND2xp5_ASAP7_75t_SL \i49/i556  (.A(\i49/n53 ),
    .B(\i49/n539 ),
    .Y(\i49/n548 ));
 AND2x2_ASAP7_75t_SL \i49/i557  (.A(n23[0]),
    .B(n23[1]),
    .Y(\i49/n549 ));
 AND2x2_ASAP7_75t_SL \i49/i558  (.A(\i49/n11 ),
    .B(\i49/n0 ),
    .Y(\i49/n550 ));
 INVx4_ASAP7_75t_SL \i49/i559  (.A(\i49/n551 ),
    .Y(\i49/n552 ));
 NOR2x1_ASAP7_75t_SL \i49/i56  (.A(\i49/n454 ),
    .B(\i49/n437 ),
    .Y(\i49/n474 ));
 NAND2x1p5_ASAP7_75t_SL \i49/i560  (.A(\i49/n549 ),
    .B(\i49/n550 ),
    .Y(\i49/n551 ));
 OAI22xp5_ASAP7_75t_SL \i49/i561  (.A1(\i49/n55 ),
    .A2(\i49/n551 ),
    .B1(\i49/n70 ),
    .B2(\i49/n75 ),
    .Y(\i49/n553 ));
 OAI221xp5_ASAP7_75t_SL \i49/i562  (.A1(\i49/n21 ),
    .A2(\i49/n89 ),
    .B1(\i49/n551 ),
    .B2(\i49/n71 ),
    .C(\i49/n172 ),
    .Y(\i49/n554 ));
 NAND2xp33_ASAP7_75t_SL \i49/i563  (.A(\i49/n551 ),
    .B(\i49/n8 ),
    .Y(\i49/n555 ));
 NOR2xp33_ASAP7_75t_SL \i49/i564  (.A(\i49/n551 ),
    .B(\i49/n50 ),
    .Y(\i49/n556 ));
 INVx2_ASAP7_75t_SL \i49/i565  (.A(\i49/n6 ),
    .Y(\i49/n557 ));
 OAI21xp5_ASAP7_75t_SL \i49/i566  (.A1(\i49/n58 ),
    .A2(\i49/n558 ),
    .B(\i49/n521 ),
    .Y(\i49/n559 ));
 AND2x4_ASAP7_75t_SL \i49/i567  (.A(\i49/n4 ),
    .B(\i49/n557 ),
    .Y(\i49/n558 ));
 OAI21xp5_ASAP7_75t_SL \i49/i568  (.A1(\i49/n76 ),
    .A2(\i49/n558 ),
    .B(\i49/n83 ),
    .Y(\i49/n560 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i49/i569  (.A1(\i49/n87 ),
    .A2(\i49/n558 ),
    .B(\i49/n72 ),
    .C(\i49/n140 ),
    .Y(\i49/n561 ));
 NOR2x1_ASAP7_75t_SL \i49/i57  (.A(\i49/n372 ),
    .B(\i49/n436 ),
    .Y(\i49/n487 ));
 NAND2xp5_ASAP7_75t_SL \i49/i570  (.A(\i49/n91 ),
    .B(\i49/n558 ),
    .Y(\i49/n562 ));
 OAI21xp5_ASAP7_75t_SL \i49/i571  (.A1(\i49/n48 ),
    .A2(\i49/n558 ),
    .B(\i49/n53 ),
    .Y(\i49/n563 ));
 AOI22xp5_ASAP7_75t_SL \i49/i572  (.A1(\i49/n53 ),
    .A2(\i49/n558 ),
    .B1(\i49/n552 ),
    .B2(\i49/n66 ),
    .Y(\i49/n564 ));
 NAND2xp5_ASAP7_75t_SL \i49/i573  (.A(\i49/n81 ),
    .B(\i49/n558 ),
    .Y(\i49/n565 ));
 NAND2xp5_ASAP7_75t_SL \i49/i574  (.A(\i49/n51 ),
    .B(\i49/n558 ),
    .Y(\i49/n566 ));
 AOI22xp5_ASAP7_75t_SL \i49/i575  (.A1(\i49/n93 ),
    .A2(\i49/n558 ),
    .B1(\i49/n65 ),
    .B2(\i49/n532 ),
    .Y(\i49/n567 ));
 NAND2xp5_ASAP7_75t_SL \i49/i576  (.A(\i49/n68 ),
    .B(\i49/n558 ),
    .Y(\i49/n568 ));
 AND2x2_ASAP7_75t_SL \i49/i577  (.A(\i49/n5 ),
    .B(\i49/n558 ),
    .Y(\i49/n569 ));
 AOI221xp5_ASAP7_75t_SL \i49/i578  (.A1(\i49/n66 ),
    .A2(\i49/n48 ),
    .B1(\i49/n558 ),
    .B2(\i49/n69 ),
    .C(\i49/n217 ),
    .Y(\i49/n570 ));
 INVx2_ASAP7_75t_SL \i49/i579  (.A(n23[5]),
    .Y(\i49/n571 ));
 INVxp67_ASAP7_75t_SL \i49/i58  (.A(\i49/n472 ),
    .Y(\i49/n473 ));
 AOI211x1_ASAP7_75t_SL \i49/i580  (.A1(\i49/n48 ),
    .A2(\i49/n72 ),
    .B(\i49/n122 ),
    .C(\i49/n450 ),
    .Y(\i49/n572 ));
 AND4x1_ASAP7_75t_SL \i49/i581  (.A(\i49/n310 ),
    .B(\i49/n354 ),
    .C(\i49/n575 ),
    .D(\i49/n282 ),
    .Y(\i49/n573 ));
 AND4x1_ASAP7_75t_SL \i49/i582  (.A(\i49/n299 ),
    .B(\i49/n357 ),
    .C(\i49/n323 ),
    .D(\i49/n310 ),
    .Y(\i49/n574 ));
 AOI21xp5_ASAP7_75t_SL \i49/i583  (.A1(\i49/n56 ),
    .A2(\i49/n532 ),
    .B(\i49/n217 ),
    .Y(\i49/n575 ));
 NOR3xp33_ASAP7_75t_SL \i49/i584  (.A(\i49/n576 ),
    .B(\i49/n341 ),
    .C(\i49/n148 ),
    .Y(\i49/n577 ));
 OAI21xp5_ASAP7_75t_SL \i49/i585  (.A1(\i49/n71 ),
    .A2(\i49/n541 ),
    .B(\i49/n171 ),
    .Y(\i49/n576 ));
 NAND3xp33_ASAP7_75t_SL \i49/i586  (.A(\i49/n578 ),
    .B(\i49/n275 ),
    .C(\i49/n346 ),
    .Y(\i49/n579 ));
 AO21x1_ASAP7_75t_SL \i49/i587  (.A1(\i49/n67 ),
    .A2(\i49/n55 ),
    .B(\i49/n86 ),
    .Y(\i49/n578 ));
 NOR3xp33_ASAP7_75t_SL \i49/i588  (.A(\i49/n580 ),
    .B(\i49/n344 ),
    .C(\i49/n218 ),
    .Y(\i49/n581 ));
 OAI21xp5_ASAP7_75t_SL \i49/i589  (.A1(\i49/n70 ),
    .A2(\i49/n534 ),
    .B(\i49/n528 ),
    .Y(\i49/n580 ));
 INVxp67_ASAP7_75t_SL \i49/i59  (.A(\i49/n468 ),
    .Y(\i49/n469 ));
 NOR2x1p5_ASAP7_75t_SL \i49/i6  (.A(\i49/n513 ),
    .B(\i49/n512 ),
    .Y(n22[4]));
 AND5x1_ASAP7_75t_SL \i49/i60  (.A(\i49/n386 ),
    .B(\i49/n575 ),
    .C(\i49/n378 ),
    .D(\i49/n297 ),
    .E(\i49/n560 ),
    .Y(\i49/n467 ));
 NOR3xp33_ASAP7_75t_SL \i49/i61  (.A(\i49/n397 ),
    .B(\i49/n377 ),
    .C(\i49/n358 ),
    .Y(\i49/n466 ));
 NOR3xp33_ASAP7_75t_SL \i49/i62  (.A(\i49/n423 ),
    .B(\i49/n359 ),
    .C(\i49/n308 ),
    .Y(\i49/n465 ));
 AND5x1_ASAP7_75t_SL \i49/i63  (.A(\i49/n349 ),
    .B(\i49/n362 ),
    .C(\i49/n342 ),
    .D(\i49/n351 ),
    .E(\i49/n277 ),
    .Y(\i49/n464 ));
 NOR2xp33_ASAP7_75t_SL \i49/i64  (.A(\i49/n424 ),
    .B(\i49/n429 ),
    .Y(\i49/n463 ));
 NAND4xp25_ASAP7_75t_SL \i49/i65  (.A(\i49/n406 ),
    .B(\i49/n414 ),
    .C(\i49/n419 ),
    .D(\i49/n402 ),
    .Y(\i49/n462 ));
 NAND5xp2_ASAP7_75t_SL \i49/i66  (.A(\i49/n385 ),
    .B(\i49/n340 ),
    .C(\i49/n236 ),
    .D(\i49/n221 ),
    .E(\i49/n13 ),
    .Y(\i49/n461 ));
 NOR4xp25_ASAP7_75t_SL \i49/i67  (.A(\i49/n375 ),
    .B(\i49/n27 ),
    .C(\i49/n325 ),
    .D(\i49/n301 ),
    .Y(\i49/n460 ));
 NAND4xp25_ASAP7_75t_SL \i49/i68  (.A(\i49/n394 ),
    .B(\i49/n408 ),
    .C(\i49/n411 ),
    .D(\i49/n413 ),
    .Y(\i49/n459 ));
 NAND4xp25_ASAP7_75t_SL \i49/i69  (.A(\i49/n421 ),
    .B(\i49/n419 ),
    .C(\i49/n203 ),
    .D(\i49/n268 ),
    .Y(\i49/n458 ));
 NOR2x2_ASAP7_75t_SL \i49/i7  (.A(\i49/n508 ),
    .B(\i49/n514 ),
    .Y(n22[3]));
 NAND3xp33_ASAP7_75t_SL \i49/i70  (.A(\i49/n413 ),
    .B(\i49/n384 ),
    .C(\i49/n548 ),
    .Y(\i49/n472 ));
 NAND4xp75_ASAP7_75t_SL \i49/i71  (.A(\i49/n316 ),
    .B(\i49/n287 ),
    .C(\i49/n371 ),
    .D(\i49/n23 ),
    .Y(\i49/n471 ));
 NAND2xp33_ASAP7_75t_L \i49/i72  (.A(\i49/n393 ),
    .B(\i49/n455 ),
    .Y(\i49/n457 ));
 AND2x2_ASAP7_75t_SL \i49/i73  (.A(\i49/n396 ),
    .B(\i49/n444 ),
    .Y(\i49/n470 ));
 NAND2x1p5_ASAP7_75t_SL \i49/i74  (.A(\i49/n452 ),
    .B(\i49/n407 ),
    .Y(\i49/n468 ));
 INVxp67_ASAP7_75t_SL \i49/i75  (.A(\i49/n455 ),
    .Y(\i49/n456 ));
 INVxp67_ASAP7_75t_SL \i49/i76  (.A(\i49/n449 ),
    .Y(\i49/n450 ));
 NOR5xp2_ASAP7_75t_SL \i49/i77  (.A(\i49/n335 ),
    .B(\i49/n307 ),
    .C(\i49/n228 ),
    .D(\i49/n192 ),
    .E(\i49/n98 ),
    .Y(\i49/n447 ));
 NOR3xp33_ASAP7_75t_SL \i49/i78  (.A(\i49/n418 ),
    .B(\i49/n330 ),
    .C(\i49/n322 ),
    .Y(\i49/n446 ));
 NOR2xp33_ASAP7_75t_SL \i49/i79  (.A(\i49/n374 ),
    .B(\i49/n395 ),
    .Y(\i49/n445 ));
 AND5x2_ASAP7_75t_SL \i49/i8  (.A(\i49/n506 ),
    .B(\i49/n497 ),
    .C(\i49/n499 ),
    .D(\i49/n484 ),
    .E(\i49/n476 ),
    .Y(n22[6]));
 NOR2xp33_ASAP7_75t_SL \i49/i80  (.A(\i49/n416 ),
    .B(\i49/n364 ),
    .Y(\i49/n444 ));
 NOR2x1_ASAP7_75t_SL \i49/i81  (.A(\i49/n379 ),
    .B(\i49/n518 ),
    .Y(\i49/n455 ));
 NAND3xp33_ASAP7_75t_SL \i49/i82  (.A(\i49/n319 ),
    .B(\i49/n348 ),
    .C(\i49/n231 ),
    .Y(\i49/n443 ));
 NAND2xp5_ASAP7_75t_L \i49/i83  (.A(\i49/n415 ),
    .B(\i49/n383 ),
    .Y(\i49/n442 ));
 NAND2xp5_ASAP7_75t_SL \i49/i84  (.A(\i49/n363 ),
    .B(\i49/n405 ),
    .Y(\i49/n441 ));
 NAND3xp33_ASAP7_75t_SL \i49/i85  (.A(\i49/n575 ),
    .B(\i49/n303 ),
    .C(\i49/n282 ),
    .Y(\i49/n454 ));
 NOR3xp33_ASAP7_75t_SL \i49/i86  (.A(\i49/n387 ),
    .B(\i49/n7 ),
    .C(\i49/n284 ),
    .Y(\i49/n440 ));
 NAND2xp5_ASAP7_75t_SL \i49/i87  (.A(\i49/n545 ),
    .B(\i49/n394 ),
    .Y(\i49/n453 ));
 OR3x1_ASAP7_75t_SL \i49/i88  (.A(\i49/n311 ),
    .B(\i49/n324 ),
    .C(\i49/n28 ),
    .Y(\i49/n439 ));
 NOR2x1_ASAP7_75t_SL \i49/i89  (.A(\i49/n322 ),
    .B(\i49/n418 ),
    .Y(\i49/n452 ));
 AND3x4_ASAP7_75t_SL \i49/i9  (.A(\i49/n506 ),
    .B(\i49/n515 ),
    .C(\i49/n494 ),
    .Y(n22[1]));
 NOR2xp33_ASAP7_75t_L \i49/i90  (.A(\i49/n376 ),
    .B(\i49/n361 ),
    .Y(\i49/n451 ));
 NOR2xp33_ASAP7_75t_SL \i49/i91  (.A(\i49/n554 ),
    .B(\i49/n404 ),
    .Y(\i49/n449 ));
 NOR3x1_ASAP7_75t_SL \i49/i92  (.A(\i49/n318 ),
    .B(\i49/n207 ),
    .C(\i49/n368 ),
    .Y(\i49/n448 ));
 NOR3xp33_ASAP7_75t_SL \i49/i93  (.A(\i49/n326 ),
    .B(\i49/n235 ),
    .C(\i49/n314 ),
    .Y(\i49/n435 ));
 NOR2xp33_ASAP7_75t_SL \i49/i94  (.A(\i49/n579 ),
    .B(\i49/n389 ),
    .Y(\i49/n434 ));
 NAND3xp33_ASAP7_75t_SL \i49/i95  (.A(\i49/n310 ),
    .B(\i49/n381 ),
    .C(\i49/n323 ),
    .Y(\i49/n433 ));
 NAND4xp25_ASAP7_75t_SL \i49/i96  (.A(\i49/n292 ),
    .B(\i49/n561 ),
    .C(\i49/n336 ),
    .D(\i49/n302 ),
    .Y(\i49/n432 ));
 NAND2x1_ASAP7_75t_SL \i49/i97  (.A(\i49/n403 ),
    .B(\i49/n417 ),
    .Y(\i49/n438 ));
 NOR5xp2_ASAP7_75t_SL \i49/i98  (.A(\i49/n412 ),
    .B(\i49/n328 ),
    .C(\i49/n133 ),
    .D(\i49/n252 ),
    .E(\i49/n173 ),
    .Y(\i49/n431 ));
 NAND3xp33_ASAP7_75t_SL \i49/i99  (.A(\i49/n367 ),
    .B(\i49/n577 ),
    .C(\i49/n238 ),
    .Y(\i49/n430 ));
 XOR2xp5_ASAP7_75t_SL i490 (.A(n617),
    .B(n618),
    .Y(n982));
 XNOR2xp5_ASAP7_75t_SL i491 (.A(n347),
    .B(n627),
    .Y(n981));
 XOR2xp5_ASAP7_75t_SL i492 (.A(n346),
    .B(n1224),
    .Y(n980));
 XNOR2xp5_ASAP7_75t_SL i493 (.A(n1178),
    .B(n344),
    .Y(n979));
 XOR2xp5_ASAP7_75t_SL i494 (.A(n815),
    .B(n619),
    .Y(n978));
 XOR2xp5_ASAP7_75t_SL i495 (.A(n343),
    .B(n798),
    .Y(n977));
 XNOR2xp5_ASAP7_75t_SL i496 (.A(n341),
    .B(n512),
    .Y(n976));
 XOR2xp5_ASAP7_75t_SL i497 (.A(n624),
    .B(n342),
    .Y(n975));
 XNOR2xp5_ASAP7_75t_SL i498 (.A(n336),
    .B(n337),
    .Y(n974));
 XOR2xp5_ASAP7_75t_SL i499 (.A(n331),
    .B(n329),
    .Y(n973));
 INVxp33_ASAP7_75t_SL i5 (.A(n30[0]),
    .Y(n88));
 INVx2_ASAP7_75t_SL \i50/i0  (.A(n21[2]),
    .Y(\i50/n0 ));
 INVx2_ASAP7_75t_SL \i50/i1  (.A(n21[0]),
    .Y(\i50/n1 ));
 NOR2x1p5_ASAP7_75t_SL \i50/i10  (.A(\i50/n505 ),
    .B(\i50/n496 ),
    .Y(n20[5]));
 NOR5xp2_ASAP7_75t_SL \i50/i100  (.A(\i50/n345 ),
    .B(\i50/n308 ),
    .C(\i50/n329 ),
    .D(\i50/n279 ),
    .E(\i50/n228 ),
    .Y(\i50/n418 ));
 NAND5xp2_ASAP7_75t_SL \i50/i101  (.A(\i50/n289 ),
    .B(\i50/n358 ),
    .C(\i50/n526 ),
    .D(\i50/n327 ),
    .E(\i50/n522 ),
    .Y(\i50/n417 ));
 NAND3xp33_ASAP7_75t_L \i50/i102  (.A(\i50/n283 ),
    .B(\i50/n312 ),
    .C(\i50/n382 ),
    .Y(\i50/n416 ));
 NOR5xp2_ASAP7_75t_SL \i50/i103  (.A(\i50/n281 ),
    .B(\i50/n293 ),
    .C(\i50/n273 ),
    .D(\i50/n122 ),
    .E(\i50/n101 ),
    .Y(\i50/n415 ));
 NAND4xp25_ASAP7_75t_SL \i50/i104  (.A(\i50/n224 ),
    .B(\i50/n235 ),
    .C(\i50/n333 ),
    .D(\i50/n18 ),
    .Y(\i50/n414 ));
 NOR5xp2_ASAP7_75t_SL \i50/i105  (.A(\i50/n239 ),
    .B(\i50/n556 ),
    .C(\i50/n510 ),
    .D(\i50/n195 ),
    .E(\i50/n193 ),
    .Y(\i50/n413 ));
 NOR2xp33_ASAP7_75t_SL \i50/i106  (.A(\i50/n372 ),
    .B(\i50/n407 ),
    .Y(\i50/n412 ));
 NOR2xp33_ASAP7_75t_SL \i50/i107  (.A(\i50/n362 ),
    .B(\i50/n392 ),
    .Y(\i50/n411 ));
 NAND3x2_ASAP7_75t_SL \i50/i108  (.B(\i50/n390 ),
    .C(\i50/n358 ),
    .Y(\i50/n427 ),
    .A(\i50/n525 ));
 NAND3x1_ASAP7_75t_SL \i50/i109  (.A(\i50/n353 ),
    .B(\i50/n334 ),
    .C(\i50/n301 ),
    .Y(\i50/n426 ));
 AND2x2_ASAP7_75t_SL \i50/i11  (.A(\i50/n506 ),
    .B(\i50/n489 ),
    .Y(n20[0]));
 AOI21xp5_ASAP7_75t_L \i50/i110  (.A1(\i50/n541 ),
    .A2(\i50/n242 ),
    .B(\i50/n170 ),
    .Y(\i50/n403 ));
 NOR2xp33_ASAP7_75t_SL \i50/i111  (.A(\i50/n560 ),
    .B(\i50/n345 ),
    .Y(\i50/n402 ));
 NAND2xp5_ASAP7_75t_SL \i50/i112  (.A(\i50/n332 ),
    .B(\i50/n361 ),
    .Y(\i50/n401 ));
 NOR2xp33_ASAP7_75t_SL \i50/i113  (.A(\i50/n360 ),
    .B(\i50/n28 ),
    .Y(\i50/n400 ));
 NOR2xp33_ASAP7_75t_SL \i50/i114  (.A(\i50/n340 ),
    .B(\i50/n350 ),
    .Y(\i50/n399 ));
 NOR2xp67_ASAP7_75t_SL \i50/i115  (.A(\i50/n180 ),
    .B(\i50/n347 ),
    .Y(\i50/n398 ));
 NOR2xp33_ASAP7_75t_SL \i50/i116  (.A(\i50/n24 ),
    .B(\i50/n345 ),
    .Y(\i50/n397 ));
 NOR4xp25_ASAP7_75t_SL \i50/i117  (.A(\i50/n316 ),
    .B(\i50/n26 ),
    .C(\i50/n24 ),
    .D(\i50/n568 ),
    .Y(\i50/n396 ));
 NAND2xp5_ASAP7_75t_SL \i50/i118  (.A(\i50/n270 ),
    .B(\i50/n324 ),
    .Y(\i50/n395 ));
 NOR4xp25_ASAP7_75t_SL \i50/i119  (.A(\i50/n119 ),
    .B(\i50/n261 ),
    .C(\i50/n230 ),
    .D(\i50/n243 ),
    .Y(\i50/n394 ));
 NOR3xp33_ASAP7_75t_SL \i50/i12  (.A(\i50/n478 ),
    .B(\i50/n474 ),
    .C(\i50/n481 ),
    .Y(\i50/n506 ));
 NOR3xp33_ASAP7_75t_SL \i50/i120  (.A(\i50/n267 ),
    .B(\i50/n223 ),
    .C(\i50/n266 ),
    .Y(\i50/n393 ));
 NAND2xp33_ASAP7_75t_SL \i50/i121  (.A(\i50/n311 ),
    .B(\i50/n25 ),
    .Y(\i50/n392 ));
 NOR2xp33_ASAP7_75t_SL \i50/i122  (.A(\i50/n560 ),
    .B(\i50/n307 ),
    .Y(\i50/n391 ));
 NOR2x1p5_ASAP7_75t_SL \i50/i123  (.A(\i50/n290 ),
    .B(\i50/n544 ),
    .Y(\i50/n390 ));
 NAND2xp33_ASAP7_75t_SL \i50/i124  (.A(\i50/n359 ),
    .B(\i50/n343 ),
    .Y(\i50/n389 ));
 NAND3xp33_ASAP7_75t_SL \i50/i125  (.A(\i50/n27 ),
    .B(\i50/n222 ),
    .C(\i50/n249 ),
    .Y(\i50/n388 ));
 NOR3xp33_ASAP7_75t_SL \i50/i126  (.A(\i50/n514 ),
    .B(\i50/n236 ),
    .C(\i50/n208 ),
    .Y(\i50/n410 ));
 NAND2xp5_ASAP7_75t_SL \i50/i127  (.A(\i50/n315 ),
    .B(\i50/n224 ),
    .Y(\i50/n409 ));
 NOR2x1_ASAP7_75t_SL \i50/i128  (.A(\i50/n288 ),
    .B(\i50/n533 ),
    .Y(\i50/n408 ));
 NAND2xp5_ASAP7_75t_SL \i50/i129  (.A(\i50/n526 ),
    .B(\i50/n317 ),
    .Y(\i50/n407 ));
 NOR2x2_ASAP7_75t_SL \i50/i13  (.A(\i50/n498 ),
    .B(\i50/n499 ),
    .Y(n20[2]));
 NOR2x1_ASAP7_75t_SL \i50/i130  (.A(\i50/n573 ),
    .B(\i50/n348 ),
    .Y(\i50/n406 ));
 NAND2xp5_ASAP7_75t_SL \i50/i131  (.A(\i50/n319 ),
    .B(\i50/n306 ),
    .Y(\i50/n387 ));
 NOR2x1_ASAP7_75t_SL \i50/i132  (.A(\i50/n26 ),
    .B(\i50/n560 ),
    .Y(\i50/n405 ));
 NOR3x1_ASAP7_75t_SL \i50/i133  (.A(\i50/n510 ),
    .B(\i50/n220 ),
    .C(\i50/n191 ),
    .Y(\i50/n404 ));
 INVx1_ASAP7_75t_SL \i50/i134  (.A(\i50/n384 ),
    .Y(\i50/n385 ));
 INVx1_ASAP7_75t_SL \i50/i135  (.A(\i50/n29 ),
    .Y(\i50/n383 ));
 NOR4xp25_ASAP7_75t_SL \i50/i136  (.A(\i50/n211 ),
    .B(\i50/n246 ),
    .C(\i50/n234 ),
    .D(\i50/n206 ),
    .Y(\i50/n382 ));
 AOI211xp5_ASAP7_75t_SL \i50/i137  (.A1(\i50/n76 ),
    .A2(\i50/n71 ),
    .B(\i50/n544 ),
    .C(\i50/n186 ),
    .Y(\i50/n381 ));
 NAND2xp33_ASAP7_75t_L \i50/i138  (.A(\i50/n302 ),
    .B(\i50/n326 ),
    .Y(\i50/n380 ));
 NAND5xp2_ASAP7_75t_SL \i50/i139  (.A(\i50/n244 ),
    .B(\i50/n259 ),
    .C(\i50/n271 ),
    .D(\i50/n188 ),
    .E(\i50/n532 ),
    .Y(\i50/n379 ));
 NAND4xp75_ASAP7_75t_SL \i50/i14  (.A(\i50/n464 ),
    .B(\i50/n484 ),
    .C(\i50/n462 ),
    .D(\i50/n571 ),
    .Y(\i50/n505 ));
 NOR4xp25_ASAP7_75t_SL \i50/i140  (.A(\i50/n336 ),
    .B(\i50/n151 ),
    .C(\i50/n153 ),
    .D(\i50/n176 ),
    .Y(\i50/n378 ));
 OAI221xp5_ASAP7_75t_SL \i50/i141  (.A1(\i50/n123 ),
    .A2(\i50/n95 ),
    .B1(\i50/n123 ),
    .B2(\i50/n16 ),
    .C(\i50/n311 ),
    .Y(\i50/n377 ));
 NOR2xp33_ASAP7_75t_SL \i50/i142  (.A(\i50/n294 ),
    .B(\i50/n297 ),
    .Y(\i50/n376 ));
 AOI211xp5_ASAP7_75t_SL \i50/i143  (.A1(\i50/n174 ),
    .A2(\i50/n77 ),
    .B(\i50/n280 ),
    .C(\i50/n197 ),
    .Y(\i50/n375 ));
 OA21x2_ASAP7_75t_SL \i50/i144  (.A1(\i50/n63 ),
    .A2(\i50/n541 ),
    .B(\i50/n565 ),
    .Y(\i50/n374 ));
 NOR4xp25_ASAP7_75t_SL \i50/i145  (.A(\i50/n274 ),
    .B(\i50/n185 ),
    .C(\i50/n216 ),
    .D(\i50/n191 ),
    .Y(\i50/n373 ));
 NAND5xp2_ASAP7_75t_SL \i50/i146  (.A(\i50/n152 ),
    .B(\i50/n106 ),
    .C(\i50/n164 ),
    .D(\i50/n155 ),
    .E(\i50/n100 ),
    .Y(\i50/n372 ));
 NOR3xp33_ASAP7_75t_SL \i50/i147  (.A(\i50/n310 ),
    .B(\i50/n187 ),
    .C(\i50/n98 ),
    .Y(\i50/n371 ));
 NAND5xp2_ASAP7_75t_SL \i50/i148  (.A(\i50/n221 ),
    .B(\i50/n113 ),
    .C(\i50/n214 ),
    .D(\i50/n205 ),
    .E(\i50/n204 ),
    .Y(\i50/n370 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i50/i149  (.A1(\i50/n79 ),
    .A2(\i50/n515 ),
    .B(\i50/n81 ),
    .C(\i50/n285 ),
    .Y(\i50/n369 ));
 NOR3xp33_ASAP7_75t_SL \i50/i15  (.A(\i50/n482 ),
    .B(\i50/n447 ),
    .C(\i50/n492 ),
    .Y(\i50/n504 ));
 NAND4xp25_ASAP7_75t_SL \i50/i150  (.A(\i50/n323 ),
    .B(\i50/n260 ),
    .C(\i50/n120 ),
    .D(\i50/n189 ),
    .Y(\i50/n368 ));
 NAND5xp2_ASAP7_75t_SL \i50/i151  (.A(\i50/n175 ),
    .B(\i50/n154 ),
    .C(\i50/n251 ),
    .D(\i50/n116 ),
    .E(\i50/n110 ),
    .Y(\i50/n367 ));
 NAND2xp5_ASAP7_75t_SL \i50/i152  (.A(\i50/n537 ),
    .B(\i50/n314 ),
    .Y(\i50/n366 ));
 NAND2xp5_ASAP7_75t_SL \i50/i153  (.A(\i50/n525 ),
    .B(\i50/n358 ),
    .Y(\i50/n365 ));
 NOR2xp33_ASAP7_75t_L \i50/i154  (.A(\i50/n338 ),
    .B(\i50/n350 ),
    .Y(\i50/n386 ));
 NAND2xp5_ASAP7_75t_SL \i50/i155  (.A(\i50/n524 ),
    .B(\i50/n359 ),
    .Y(\i50/n364 ));
 NOR2x1p5_ASAP7_75t_SL \i50/i156  (.A(\i50/n511 ),
    .B(\i50/n341 ),
    .Y(\i50/n384 ));
 NAND3x1_ASAP7_75t_SL \i50/i157  (.A(\i50/n278 ),
    .B(\i50/n528 ),
    .C(\i50/n158 ),
    .Y(\i50/n29 ));
 INVxp67_ASAP7_75t_SL \i50/i158  (.A(\i50/n362 ),
    .Y(\i50/n363 ));
 INVxp67_ASAP7_75t_SL \i50/i159  (.A(\i50/n7 ),
    .Y(\i50/n361 ));
 NAND4xp75_ASAP7_75t_SL \i50/i16  (.A(\i50/n463 ),
    .B(\i50/n494 ),
    .C(\i50/n468 ),
    .D(\i50/n458 ),
    .Y(\i50/n503 ));
 INVxp67_ASAP7_75t_SL \i50/i160  (.A(\i50/n356 ),
    .Y(\i50/n357 ));
 INVxp67_ASAP7_75t_SL \i50/i161  (.A(\i50/n354 ),
    .Y(\i50/n355 ));
 INVx2_ASAP7_75t_SL \i50/i162  (.A(\i50/n352 ),
    .Y(\i50/n353 ));
 INVxp67_ASAP7_75t_SL \i50/i163  (.A(\i50/n348 ),
    .Y(\i50/n349 ));
 INVxp67_ASAP7_75t_SL \i50/i164  (.A(\i50/n564 ),
    .Y(\i50/n346 ));
 INVx1_ASAP7_75t_SL \i50/i165  (.A(\i50/n343 ),
    .Y(\i50/n344 ));
 OAI31xp33_ASAP7_75t_SL \i50/i166  (.A1(\i50/n77 ),
    .A2(\i50/n2 ),
    .A3(\i50/n60 ),
    .B(\i50/n55 ),
    .Y(\i50/n342 ));
 NAND2x1_ASAP7_75t_SL \i50/i167  (.A(\i50/n233 ),
    .B(\i50/n232 ),
    .Y(\i50/n341 ));
 NAND2xp33_ASAP7_75t_SL \i50/i168  (.A(\i50/n222 ),
    .B(\i50/n526 ),
    .Y(\i50/n340 ));
 OAI21xp5_ASAP7_75t_SL \i50/i169  (.A1(\i50/n57 ),
    .A2(\i50/n145 ),
    .B(\i50/n202 ),
    .Y(\i50/n339 ));
 AND3x4_ASAP7_75t_SL \i50/i17  (.A(\i50/n485 ),
    .B(\i50/n500 ),
    .C(\i50/n490 ),
    .Y(n20[7]));
 NAND2xp5_ASAP7_75t_SL \i50/i170  (.A(\i50/n190 ),
    .B(\i50/n222 ),
    .Y(\i50/n338 ));
 AOI211xp5_ASAP7_75t_SL \i50/i171  (.A1(\i50/n93 ),
    .A2(\i50/n34 ),
    .B(\i50/n530 ),
    .C(\i50/n130 ),
    .Y(\i50/n337 ));
 AOI31xp33_ASAP7_75t_SL \i50/i172  (.A1(\i50/n57 ),
    .A2(\i50/n17 ),
    .A3(\i50/n68 ),
    .B(\i50/n51 ),
    .Y(\i50/n336 ));
 NOR3xp33_ASAP7_75t_SL \i50/i173  (.A(\i50/n223 ),
    .B(\i50/n144 ),
    .C(\i50/n128 ),
    .Y(\i50/n335 ));
 NOR3xp33_ASAP7_75t_SL \i50/i174  (.A(\i50/n531 ),
    .B(\i50/n137 ),
    .C(\i50/n272 ),
    .Y(\i50/n334 ));
 OAI31xp33_ASAP7_75t_SL \i50/i175  (.A1(\i50/n53 ),
    .A2(\i50/n55 ),
    .A3(\i50/n74 ),
    .B(\i50/n93 ),
    .Y(\i50/n333 ));
 AOI221xp5_ASAP7_75t_SL \i50/i176  (.A1(\i50/n79 ),
    .A2(\i50/n96 ),
    .B1(\i50/n563 ),
    .B2(\i50/n69 ),
    .C(\i50/n207 ),
    .Y(\i50/n332 ));
 OAI31xp33_ASAP7_75t_R \i50/i177  (.A1(\i50/n77 ),
    .A2(\i50/n550 ),
    .A3(\i50/n79 ),
    .B(\i50/n74 ),
    .Y(\i50/n331 ));
 AOI21xp5_ASAP7_75t_SL \i50/i178  (.A1(\i50/n170 ),
    .A2(\i50/n68 ),
    .B(\i50/n91 ),
    .Y(\i50/n362 ));
 AOI21xp5_ASAP7_75t_L \i50/i179  (.A1(\i50/n68 ),
    .A2(\i50/n181 ),
    .B(\i50/n90 ),
    .Y(\i50/n330 ));
 NAND4xp75_ASAP7_75t_SL \i50/i18  (.A(\i50/n578 ),
    .B(\i50/n467 ),
    .C(\i50/n476 ),
    .D(\i50/n493 ),
    .Y(\i50/n502 ));
 OAI221xp5_ASAP7_75t_SL \i50/i180  (.A1(\i50/n535 ),
    .A2(\i50/n95 ),
    .B1(\i50/n54 ),
    .B2(\i50/n61 ),
    .C(\i50/n229 ),
    .Y(\i50/n329 ));
 AOI21xp33_ASAP7_75t_SL \i50/i181  (.A1(\i50/n181 ),
    .A2(\i50/n52 ),
    .B(\i50/n539 ),
    .Y(\i50/n328 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i50/i182  (.A1(\i50/n88 ),
    .A2(\i50/n4 ),
    .B(\i50/n92 ),
    .C(\i50/n19 ),
    .Y(\i50/n327 ));
 NOR3xp33_ASAP7_75t_SL \i50/i183  (.A(\i50/n240 ),
    .B(\i50/n531 ),
    .C(\i50/n149 ),
    .Y(\i50/n326 ));
 NAND3xp33_ASAP7_75t_SL \i50/i184  (.A(\i50/n20 ),
    .B(\i50/n23 ),
    .C(\i50/n179 ),
    .Y(\i50/n325 ));
 AOI22xp5_ASAP7_75t_SL \i50/i185  (.A1(\i50/n65 ),
    .A2(\i50/n166 ),
    .B1(\i50/n69 ),
    .B2(\i50/n60 ),
    .Y(\i50/n324 ));
 OAI21xp5_ASAP7_75t_SL \i50/i186  (.A1(\i50/n67 ),
    .A2(\i50/n172 ),
    .B(\i50/n77 ),
    .Y(\i50/n323 ));
 NAND4xp25_ASAP7_75t_SL \i50/i187  (.A(\i50/n194 ),
    .B(\i50/n189 ),
    .C(\i50/n156 ),
    .D(\i50/n159 ),
    .Y(\i50/n322 ));
 NAND2xp33_ASAP7_75t_SL \i50/i188  (.A(\i50/n254 ),
    .B(\i50/n148 ),
    .Y(\i50/n321 ));
 OAI211xp5_ASAP7_75t_SL \i50/i189  (.A1(\i50/n72 ),
    .A2(\i50/n539 ),
    .B(\i50/n161 ),
    .C(\i50/n165 ),
    .Y(\i50/n360 ));
 NAND2x1_ASAP7_75t_SL \i50/i19  (.A(\i50/n486 ),
    .B(\i50/n455 ),
    .Y(\i50/n501 ));
 NOR2xp67_ASAP7_75t_SL \i50/i190  (.A(\i50/n566 ),
    .B(\i50/n273 ),
    .Y(\i50/n359 ));
 AOI21x1_ASAP7_75t_SL \i50/i191  (.A1(\i50/n60 ),
    .A2(\i50/n67 ),
    .B(\i50/n280 ),
    .Y(\i50/n358 ));
 NAND2xp5_ASAP7_75t_SL \i50/i192  (.A(\i50/n256 ),
    .B(\i50/n520 ),
    .Y(\i50/n28 ));
 NOR2xp33_ASAP7_75t_SL \i50/i193  (.A(\i50/n257 ),
    .B(\i50/n274 ),
    .Y(\i50/n356 ));
 OAI211xp5_ASAP7_75t_SL \i50/i194  (.A1(\i50/n68 ),
    .A2(\i50/n539 ),
    .B(\i50/n202 ),
    .C(\i50/n203 ),
    .Y(\i50/n354 ));
 OR2x2_ASAP7_75t_SL \i50/i195  (.A(\i50/n213 ),
    .B(\i50/n567 ),
    .Y(\i50/n352 ));
 OAI211xp5_ASAP7_75t_SL \i50/i196  (.A1(\i50/n95 ),
    .A2(\i50/n82 ),
    .B(\i50/n198 ),
    .C(\i50/n139 ),
    .Y(\i50/n351 ));
 NAND2xp5_ASAP7_75t_SL \i50/i197  (.A(\i50/n522 ),
    .B(\i50/n275 ),
    .Y(\i50/n350 ));
 NAND2xp5_ASAP7_75t_SL \i50/i198  (.A(\i50/n27 ),
    .B(\i50/n209 ),
    .Y(\i50/n348 ));
 NAND2xp5_ASAP7_75t_SL \i50/i199  (.A(\i50/n253 ),
    .B(\i50/n523 ),
    .Y(\i50/n347 ));
 INVx2_ASAP7_75t_SL \i50/i2  (.A(\i50/n9 ),
    .Y(\i50/n2 ));
 NOR2xp67_ASAP7_75t_SL \i50/i20  (.A(\i50/n487 ),
    .B(\i50/n448 ),
    .Y(\i50/n500 ));
 NAND2xp5_ASAP7_75t_SL \i50/i200  (.A(\i50/n196 ),
    .B(\i50/n217 ),
    .Y(\i50/n345 ));
 NOR2x1_ASAP7_75t_SL \i50/i201  (.A(\i50/n255 ),
    .B(\i50/n228 ),
    .Y(\i50/n343 ));
 INVxp67_ASAP7_75t_SL \i50/i202  (.A(\i50/n316 ),
    .Y(\i50/n317 ));
 INVx1_ASAP7_75t_SL \i50/i203  (.A(\i50/n312 ),
    .Y(\i50/n313 ));
 NAND4xp25_ASAP7_75t_SL \i50/i204  (.A(\i50/n121 ),
    .B(\i50/n140 ),
    .C(\i50/n125 ),
    .D(\i50/n124 ),
    .Y(\i50/n305 ));
 AOI31xp33_ASAP7_75t_SL \i50/i205  (.A1(\i50/n141 ),
    .A2(\i50/n541 ),
    .A3(\i50/n51 ),
    .B(\i50/n52 ),
    .Y(\i50/n304 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i50/i206  (.A1(\i50/n92 ),
    .A2(\i50/n56 ),
    .B(\i50/n74 ),
    .C(\i50/n545 ),
    .Y(\i50/n303 ));
 NOR4xp25_ASAP7_75t_SL \i50/i207  (.A(\i50/n119 ),
    .B(\i50/n131 ),
    .C(\i50/n201 ),
    .D(\i50/n97 ),
    .Y(\i50/n302 ));
 AOI211xp5_ASAP7_75t_SL \i50/i208  (.A1(\i50/n142 ),
    .A2(\i50/n85 ),
    .B(\i50/n187 ),
    .C(\i50/n104 ),
    .Y(\i50/n301 ));
 AOI21xp5_ASAP7_75t_R \i50/i209  (.A1(\i50/n171 ),
    .A2(\i50/n92 ),
    .B(\i50/n245 ),
    .Y(\i50/n300 ));
 NAND4xp75_ASAP7_75t_SL \i50/i21  (.A(\i50/n459 ),
    .B(\i50/n471 ),
    .C(\i50/n453 ),
    .D(\i50/n456 ),
    .Y(\i50/n499 ));
 NOR2xp33_ASAP7_75t_L \i50/i210  (.A(\i50/n562 ),
    .B(\i50/n268 ),
    .Y(\i50/n299 ));
 OAI31xp33_ASAP7_75t_SL \i50/i211  (.A1(\i50/n65 ),
    .A2(\i50/n563 ),
    .A3(\i50/n93 ),
    .B(\i50/n551 ),
    .Y(\i50/n298 ));
 OAI22xp5_ASAP7_75t_SL \i50/i212  (.A1(\i50/n82 ),
    .A2(\i50/n173 ),
    .B1(\i50/n72 ),
    .B2(\i50/n103 ),
    .Y(\i50/n297 ));
 NOR2xp33_ASAP7_75t_SL \i50/i213  (.A(\i50/n226 ),
    .B(\i50/n512 ),
    .Y(\i50/n296 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i50/i214  (.A1(\i50/n65 ),
    .A2(\i50/n62 ),
    .B(\i50/n4 ),
    .C(\i50/n183 ),
    .Y(\i50/n295 ));
 NAND2xp33_ASAP7_75t_L \i50/i215  (.A(\i50/n118 ),
    .B(\i50/n218 ),
    .Y(\i50/n294 ));
 NAND2xp33_ASAP7_75t_SL \i50/i216  (.A(\i50/n264 ),
    .B(\i50/n138 ),
    .Y(\i50/n293 ));
 AOI22xp5_ASAP7_75t_SL \i50/i217  (.A1(\i50/n550 ),
    .A2(\i50/n115 ),
    .B1(\i50/n85 ),
    .B2(\i50/n79 ),
    .Y(\i50/n292 ));
 OA21x2_ASAP7_75t_SL \i50/i218  (.A1(\i50/n52 ),
    .A2(\i50/n145 ),
    .B(\i50/n133 ),
    .Y(\i50/n291 ));
 NAND4xp25_ASAP7_75t_SL \i50/i219  (.A(\i50/n135 ),
    .B(\i50/n160 ),
    .C(\i50/n112 ),
    .D(\i50/n109 ),
    .Y(\i50/n290 ));
 OR3x1_ASAP7_75t_SL \i50/i22  (.A(\i50/n479 ),
    .B(\i50/n477 ),
    .C(\i50/n460 ),
    .Y(\i50/n498 ));
 AOI221xp5_ASAP7_75t_SL \i50/i220  (.A1(\i50/n69 ),
    .A2(\i50/n50 ),
    .B1(\i50/n56 ),
    .B2(\i50/n71 ),
    .C(\i50/n561 ),
    .Y(\i50/n289 ));
 OAI221xp5_ASAP7_75t_SL \i50/i221  (.A1(\i50/n94 ),
    .A2(\i50/n87 ),
    .B1(\i50/n75 ),
    .B2(\i50/n16 ),
    .C(\i50/n117 ),
    .Y(\i50/n320 ));
 OAI222xp33_ASAP7_75t_SL \i50/i222  (.A1(\i50/n9 ),
    .A2(\i50/n57 ),
    .B1(\i50/n61 ),
    .B2(\i50/n72 ),
    .C1(\i50/n75 ),
    .C2(\i50/n80 ),
    .Y(\i50/n288 ));
 OAI221xp5_ASAP7_75t_SL \i50/i223  (.A1(\i50/n90 ),
    .A2(\i50/n80 ),
    .B1(\i50/n75 ),
    .B2(\i50/n73 ),
    .C(\i50/n227 ),
    .Y(\i50/n287 ));
 AND3x1_ASAP7_75t_SL \i50/i224  (.A(\i50/n132 ),
    .B(\i50/n140 ),
    .C(\i50/n247 ),
    .Y(\i50/n286 ));
 AOI22xp5_ASAP7_75t_SL \i50/i225  (.A1(\i50/n89 ),
    .A2(\i50/n168 ),
    .B1(\i50/n67 ),
    .B2(\i50/n92 ),
    .Y(\i50/n319 ));
 NAND2xp33_ASAP7_75t_SL \i50/i226  (.A(\i50/n215 ),
    .B(\i50/n248 ),
    .Y(\i50/n285 ));
 OAI221xp5_ASAP7_75t_SL \i50/i227  (.A1(\i50/n90 ),
    .A2(\i50/n84 ),
    .B1(\i50/n535 ),
    .B2(\i50/n17 ),
    .C(\i50/n263 ),
    .Y(\i50/n284 ));
 OAI222xp33_ASAP7_75t_SL \i50/i228  (.A1(\i50/n82 ),
    .A2(\i50/n84 ),
    .B1(\i50/n94 ),
    .B2(\i50/n80 ),
    .C1(\i50/n535 ),
    .C2(\i50/n68 ),
    .Y(\i50/n318 ));
 NAND3x1_ASAP7_75t_SL \i50/i229  (.A(\i50/n219 ),
    .B(\i50/n163 ),
    .C(\i50/n157 ),
    .Y(\i50/n316 ));
 OR3x1_ASAP7_75t_SL \i50/i23  (.A(\i50/n480 ),
    .B(\i50/n446 ),
    .C(\i50/n420 ),
    .Y(\i50/n497 ));
 AOI22xp5_ASAP7_75t_SL \i50/i230  (.A1(\i50/n162 ),
    .A2(\i50/n93 ),
    .B1(\i50/n74 ),
    .B2(\i50/n563 ),
    .Y(\i50/n315 ));
 AOI22xp5_ASAP7_75t_SL \i50/i231  (.A1(\i50/n96 ),
    .A2(\i50/n107 ),
    .B1(\i50/n53 ),
    .B2(\i50/n77 ),
    .Y(\i50/n314 ));
 AOI221x1_ASAP7_75t_SL \i50/i232  (.A1(\i50/n93 ),
    .A2(\i50/n74 ),
    .B1(\i50/n79 ),
    .B2(\i50/n81 ),
    .C(\i50/n250 ),
    .Y(\i50/n312 ));
 AOI211x1_ASAP7_75t_SL \i50/i233  (.A1(\i50/n108 ),
    .A2(\i50/n70 ),
    .B(\i50/n199 ),
    .C(\i50/n201 ),
    .Y(\i50/n311 ));
 OAI21xp5_ASAP7_75t_SL \i50/i234  (.A1(\i50/n51 ),
    .A2(\i50/n87 ),
    .B(\i50/n258 ),
    .Y(\i50/n310 ));
 NOR2x1_ASAP7_75t_SL \i50/i235  (.A(\i50/n134 ),
    .B(\i50/n212 ),
    .Y(\i50/n309 ));
 OAI221xp5_ASAP7_75t_SL \i50/i236  (.A1(\i50/n22 ),
    .A2(\i50/n94 ),
    .B1(\i50/n66 ),
    .B2(\i50/n73 ),
    .C(\i50/n177 ),
    .Y(\i50/n308 ));
 OAI211xp5_ASAP7_75t_SL \i50/i237  (.A1(\i50/n73 ),
    .A2(\i50/n111 ),
    .B(\i50/n120 ),
    .C(\i50/n519 ),
    .Y(\i50/n307 ));
 NOR2xp33_ASAP7_75t_SL \i50/i238  (.A(\i50/n146 ),
    .B(\i50/n277 ),
    .Y(\i50/n283 ));
 AOI222xp33_ASAP7_75t_SL \i50/i239  (.A1(\i50/n79 ),
    .A2(\i50/n69 ),
    .B1(\i50/n4 ),
    .B2(\i50/n50 ),
    .C1(\i50/n77 ),
    .C2(\i50/n67 ),
    .Y(\i50/n306 ));
 NAND3xp33_ASAP7_75t_SL \i50/i24  (.A(\i50/n491 ),
    .B(\i50/n476 ),
    .C(\i50/n459 ),
    .Y(\i50/n496 ));
 INVx1_ASAP7_75t_SL \i50/i240  (.A(\i50/n523 ),
    .Y(\i50/n281 ));
 INVx1_ASAP7_75t_SL \i50/i241  (.A(\i50/n277 ),
    .Y(\i50/n278 ));
 INVxp67_ASAP7_75t_SL \i50/i242  (.A(\i50/n275 ),
    .Y(\i50/n276 ));
 INVxp67_ASAP7_75t_SL \i50/i243  (.A(\i50/n552 ),
    .Y(\i50/n271 ));
 INVx1_ASAP7_75t_SL \i50/i244  (.A(\i50/n268 ),
    .Y(\i50/n269 ));
 OAI21xp33_ASAP7_75t_SL \i50/i245  (.A1(\i50/n78 ),
    .A2(\i50/n540 ),
    .B(\i50/n192 ),
    .Y(\i50/n266 ));
 NAND2xp5_ASAP7_75t_SL \i50/i246  (.A(\i50/n102 ),
    .B(\i50/n139 ),
    .Y(\i50/n265 ));
 OAI21xp5_ASAP7_75t_SL \i50/i247  (.A1(\i50/n563 ),
    .A2(\i50/n60 ),
    .B(\i50/n88 ),
    .Y(\i50/n264 ));
 NOR2xp33_ASAP7_75t_SL \i50/i248  (.A(\i50/n147 ),
    .B(\i50/n186 ),
    .Y(\i50/n263 ));
 AOI21xp5_ASAP7_75t_SL \i50/i249  (.A1(\i50/n542 ),
    .A2(\i50/n57 ),
    .B(\i50/n91 ),
    .Y(\i50/n262 ));
 NOR2x1_ASAP7_75t_SL \i50/i25  (.A(\i50/n401 ),
    .B(\i50/n477 ),
    .Y(\i50/n494 ));
 NAND2xp33_ASAP7_75t_L \i50/i250  (.A(\i50/n182 ),
    .B(\i50/n105 ),
    .Y(\i50/n261 ));
 OAI21xp5_ASAP7_75t_SL \i50/i251  (.A1(\i50/n76 ),
    .A2(\i50/n62 ),
    .B(\i50/n55 ),
    .Y(\i50/n260 ));
 NOR2xp33_ASAP7_75t_SL \i50/i252  (.A(\i50/n19 ),
    .B(\i50/n126 ),
    .Y(\i50/n259 ));
 OAI21xp5_ASAP7_75t_SL \i50/i253  (.A1(\i50/n550 ),
    .A2(\i50/n86 ),
    .B(\i50/n69 ),
    .Y(\i50/n258 ));
 OAI21xp5_ASAP7_75t_SL \i50/i254  (.A1(\i50/n63 ),
    .A2(\i50/n91 ),
    .B(\i50/n184 ),
    .Y(\i50/n257 ));
 AOI22xp5_ASAP7_75t_SL \i50/i255  (.A1(\i50/n88 ),
    .A2(\i50/n62 ),
    .B1(\i50/n81 ),
    .B2(\i50/n77 ),
    .Y(\i50/n256 ));
 OAI21xp5_ASAP7_75t_SL \i50/i256  (.A1(\i50/n17 ),
    .A2(\i50/n75 ),
    .B(\i50/n143 ),
    .Y(\i50/n255 ));
 OAI21xp5_ASAP7_75t_SL \i50/i257  (.A1(\i50/n550 ),
    .A2(\i50/n60 ),
    .B(\i50/n71 ),
    .Y(\i50/n254 ));
 AOI22xp5_ASAP7_75t_SL \i50/i258  (.A1(\i50/n50 ),
    .A2(\i50/n96 ),
    .B1(\i50/n53 ),
    .B2(\i50/n550 ),
    .Y(\i50/n253 ));
 OA21x2_ASAP7_75t_SL \i50/i259  (.A1(\i50/n542 ),
    .A2(\i50/n59 ),
    .B(\i50/n188 ),
    .Y(\i50/n282 ));
 NOR2x1_ASAP7_75t_SL \i50/i26  (.A(\i50/n461 ),
    .B(\i50/n457 ),
    .Y(\i50/n493 ));
 AOI21xp33_ASAP7_75t_SL \i50/i260  (.A1(\i50/n72 ),
    .A2(\i50/n542 ),
    .B(\i50/n51 ),
    .Y(\i50/n252 ));
 OAI21xp5_ASAP7_75t_SL \i50/i261  (.A1(\i50/n81 ),
    .A2(\i50/n96 ),
    .B(\i50/n89 ),
    .Y(\i50/n251 ));
 OA21x2_ASAP7_75t_SL \i50/i262  (.A1(\i50/n4 ),
    .A2(\i50/n96 ),
    .B(\i50/n92 ),
    .Y(\i50/n250 ));
 AOI22xp33_ASAP7_75t_SL \i50/i263  (.A1(\i50/n96 ),
    .A2(\i50/n563 ),
    .B1(\i50/n70 ),
    .B2(\i50/n2 ),
    .Y(\i50/n249 ));
 OAI21xp5_ASAP7_75t_SL \i50/i264  (.A1(\i50/n71 ),
    .A2(\i50/n53 ),
    .B(\i50/n89 ),
    .Y(\i50/n248 ));
 OAI21xp5_ASAP7_75t_SL \i50/i265  (.A1(\i50/n550 ),
    .A2(\i50/n76 ),
    .B(\i50/n96 ),
    .Y(\i50/n247 ));
 AOI21xp33_ASAP7_75t_SL \i50/i266  (.A1(\i50/n68 ),
    .A2(\i50/n87 ),
    .B(\i50/n51 ),
    .Y(\i50/n246 ));
 OAI21xp5_ASAP7_75t_SL \i50/i267  (.A1(\i50/n63 ),
    .A2(\i50/n75 ),
    .B(\i50/n25 ),
    .Y(\i50/n245 ));
 AOI22xp5_ASAP7_75t_SL \i50/i268  (.A1(\i50/n67 ),
    .A2(\i50/n65 ),
    .B1(\i50/n81 ),
    .B2(\i50/n62 ),
    .Y(\i50/n244 ));
 AOI21xp33_ASAP7_75t_SL \i50/i269  (.A1(\i50/n539 ),
    .A2(\i50/n51 ),
    .B(\i50/n73 ),
    .Y(\i50/n243 ));
 NAND3xp33_ASAP7_75t_SL \i50/i27  (.A(\i50/n442 ),
    .B(\i50/n575 ),
    .C(\i50/n440 ),
    .Y(\i50/n492 ));
 OAI21xp5_ASAP7_75t_SL \i50/i270  (.A1(\i50/n92 ),
    .A2(\i50/n550 ),
    .B(\i50/n55 ),
    .Y(\i50/n242 ));
 OAI21xp5_ASAP7_75t_SL \i50/i271  (.A1(\i50/n76 ),
    .A2(\i50/n65 ),
    .B(\i50/n81 ),
    .Y(\i50/n241 ));
 NAND2xp5_ASAP7_75t_SL \i50/i272  (.A(\i50/n89 ),
    .B(\i50/n171 ),
    .Y(\i50/n27 ));
 NAND2xp5_ASAP7_75t_L \i50/i273  (.A(\i50/n202 ),
    .B(\i50/n203 ),
    .Y(\i50/n240 ));
 OAI22xp5_ASAP7_75t_SL \i50/i274  (.A1(\i50/n540 ),
    .A2(\i50/n90 ),
    .B1(\i50/n521 ),
    .B2(\i50/n59 ),
    .Y(\i50/n280 ));
 OAI22xp5_ASAP7_75t_SL \i50/i275  (.A1(\i50/n521 ),
    .A2(\i50/n75 ),
    .B1(\i50/n535 ),
    .B2(\i50/n72 ),
    .Y(\i50/n279 ));
 OAI22xp5_ASAP7_75t_SL \i50/i276  (.A1(\i50/n95 ),
    .A2(\i50/n61 ),
    .B1(\i50/n63 ),
    .B2(\i50/n82 ),
    .Y(\i50/n277 ));
 AOI22xp5_ASAP7_75t_SL \i50/i277  (.A1(\i50/n70 ),
    .A2(\i50/n93 ),
    .B1(\i50/n4 ),
    .B2(\i50/n86 ),
    .Y(\i50/n275 ));
 OAI22xp5_ASAP7_75t_SL \i50/i278  (.A1(\i50/n73 ),
    .A2(\i50/n82 ),
    .B1(\i50/n75 ),
    .B2(\i50/n54 ),
    .Y(\i50/n274 ));
 OAI22xp33_ASAP7_75t_SL \i50/i279  (.A1(\i50/n521 ),
    .A2(\i50/n94 ),
    .B1(\i50/n52 ),
    .B2(\i50/n9 ),
    .Y(\i50/n273 ));
 NOR2x1_ASAP7_75t_SL \i50/i28  (.A(\i50/n466 ),
    .B(\i50/n429 ),
    .Y(\i50/n491 ));
 NAND2xp5_ASAP7_75t_L \i50/i280  (.A(\i50/n18 ),
    .B(\i50/n167 ),
    .Y(\i50/n272 ));
 OAI21xp5_ASAP7_75t_SL \i50/i281  (.A1(\i50/n550 ),
    .A2(\i50/n56 ),
    .B(\i50/n88 ),
    .Y(\i50/n270 ));
 NOR2xp33_ASAP7_75t_L \i50/i282  (.A(\i50/n59 ),
    .B(\i50/n22 ),
    .Y(\i50/n268 ));
 NAND2xp33_ASAP7_75t_L \i50/i283  (.A(\i50/n120 ),
    .B(\i50/n519 ),
    .Y(\i50/n239 ));
 OAI21xp5_ASAP7_75t_SL \i50/i284  (.A1(\i50/n73 ),
    .A2(\i50/n61 ),
    .B(\i50/n532 ),
    .Y(\i50/n267 ));
 INVxp67_ASAP7_75t_SL \i50/i285  (.A(\i50/n237 ),
    .Y(\i50/n238 ));
 INVxp67_ASAP7_75t_SL \i50/i286  (.A(\i50/n235 ),
    .Y(\i50/n236 ));
 INVx1_ASAP7_75t_SL \i50/i287  (.A(\i50/n233 ),
    .Y(\i50/n234 ));
 INVx1_ASAP7_75t_SL \i50/i288  (.A(\i50/n231 ),
    .Y(\i50/n232 ));
 INVxp67_ASAP7_75t_SL \i50/i289  (.A(\i50/n229 ),
    .Y(\i50/n230 ));
 NOR5xp2_ASAP7_75t_SL \i50/i29  (.A(\i50/n431 ),
    .B(\i50/n379 ),
    .C(\i50/n422 ),
    .D(\i50/n347 ),
    .E(\i50/n351 ),
    .Y(\i50/n490 ));
 INVxp67_ASAP7_75t_R \i50/i290  (.A(\i50/n226 ),
    .Y(\i50/n227 ));
 INVxp67_ASAP7_75t_SL \i50/i291  (.A(\i50/n514 ),
    .Y(\i50/n225 ));
 OAI21xp5_ASAP7_75t_SL \i50/i292  (.A1(\i50/n62 ),
    .A2(\i50/n83 ),
    .B(\i50/n81 ),
    .Y(\i50/n221 ));
 OAI21xp5_ASAP7_75t_SL \i50/i293  (.A1(\i50/n16 ),
    .A2(\i50/n9 ),
    .B(\i50/n129 ),
    .Y(\i50/n220 ));
 OAI21xp5_ASAP7_75t_SL \i50/i294  (.A1(\i50/n64 ),
    .A2(\i50/n74 ),
    .B(\i50/n76 ),
    .Y(\i50/n219 ));
 OAI21xp5_ASAP7_75t_SL \i50/i295  (.A1(\i50/n563 ),
    .A2(\i50/n56 ),
    .B(\i50/n64 ),
    .Y(\i50/n218 ));
 AOI22xp5_ASAP7_75t_SL \i50/i296  (.A1(\i50/n85 ),
    .A2(\i50/n65 ),
    .B1(\i50/n55 ),
    .B2(\i50/n2 ),
    .Y(\i50/n217 ));
 AOI21xp33_ASAP7_75t_SL \i50/i297  (.A1(\i50/n75 ),
    .A2(\i50/n82 ),
    .B(\i50/n84 ),
    .Y(\i50/n216 ));
 OAI21xp5_ASAP7_75t_SL \i50/i298  (.A1(\i50/n50 ),
    .A2(\i50/n56 ),
    .B(\i50/n55 ),
    .Y(\i50/n215 ));
 OAI21xp5_ASAP7_75t_SL \i50/i299  (.A1(\i50/n85 ),
    .A2(\i50/n64 ),
    .B(\i50/n563 ),
    .Y(\i50/n214 ));
 INVx1_ASAP7_75t_SL \i50/i3  (.A(\i50/n557 ),
    .Y(\i50/n3 ));
 NOR3xp33_ASAP7_75t_SL \i50/i30  (.A(\i50/n427 ),
    .B(\i50/n444 ),
    .C(\i50/n475 ),
    .Y(\i50/n489 ));
 OAI22xp33_ASAP7_75t_SL \i50/i300  (.A1(\i50/n540 ),
    .A2(\i50/n51 ),
    .B1(\i50/n90 ),
    .B2(\i50/n68 ),
    .Y(\i50/n213 ));
 OAI22xp33_ASAP7_75t_SL \i50/i301  (.A1(\i50/n535 ),
    .A2(\i50/n540 ),
    .B1(\i50/n82 ),
    .B2(\i50/n87 ),
    .Y(\i50/n212 ));
 OAI22xp5_ASAP7_75t_SL \i50/i302  (.A1(\i50/n95 ),
    .A2(\i50/n9 ),
    .B1(\i50/n16 ),
    .B2(\i50/n90 ),
    .Y(\i50/n211 ));
 OAI22xp5_ASAP7_75t_SL \i50/i303  (.A1(\i50/n68 ),
    .A2(\i50/n9 ),
    .B1(\i50/n87 ),
    .B2(\i50/n539 ),
    .Y(\i50/n210 ));
 AOI22xp5_ASAP7_75t_SL \i50/i304  (.A1(\i50/n69 ),
    .A2(\i50/n83 ),
    .B1(\i50/n53 ),
    .B2(\i50/n86 ),
    .Y(\i50/n209 ));
 OAI22xp5_ASAP7_75t_SL \i50/i305  (.A1(\i50/n540 ),
    .A2(\i50/n94 ),
    .B1(\i50/n72 ),
    .B2(\i50/n59 ),
    .Y(\i50/n208 ));
 OAI21xp5_ASAP7_75t_SL \i50/i306  (.A1(\i50/n52 ),
    .A2(\i50/n61 ),
    .B(\i50/n127 ),
    .Y(\i50/n237 ));
 AOI22xp5_ASAP7_75t_SL \i50/i307  (.A1(\i50/n50 ),
    .A2(\i50/n71 ),
    .B1(\i50/n53 ),
    .B2(\i50/n60 ),
    .Y(\i50/n235 ));
 AOI22xp5_ASAP7_75t_SL \i50/i308  (.A1(\i50/n55 ),
    .A2(\i50/n56 ),
    .B1(\i50/n65 ),
    .B2(\i50/n69 ),
    .Y(\i50/n233 ));
 OAI22xp5_ASAP7_75t_SL \i50/i309  (.A1(\i50/n51 ),
    .A2(\i50/n16 ),
    .B1(\i50/n540 ),
    .B2(\i50/n541 ),
    .Y(\i50/n207 ));
 NOR2x1_ASAP7_75t_SL \i50/i31  (.A(\i50/n472 ),
    .B(\i50/n432 ),
    .Y(\i50/n488 ));
 NAND2xp33_ASAP7_75t_SL \i50/i310  (.A(\i50/n204 ),
    .B(\i50/n205 ),
    .Y(\i50/n206 ));
 OAI22x1_ASAP7_75t_SL \i50/i311  (.A1(\i50/n17 ),
    .A2(\i50/n94 ),
    .B1(\i50/n54 ),
    .B2(\i50/n78 ),
    .Y(\i50/n231 ));
 AOI22xp5_ASAP7_75t_SL \i50/i312  (.A1(\i50/n55 ),
    .A2(\i50/n65 ),
    .B1(\i50/n53 ),
    .B2(\i50/n92 ),
    .Y(\i50/n229 ));
 AO22x2_ASAP7_75t_SL \i50/i313  (.A1(\i50/n96 ),
    .A2(\i50/n93 ),
    .B1(\i50/n58 ),
    .B2(\i50/n86 ),
    .Y(\i50/n228 ));
 OAI22xp33_ASAP7_75t_SL \i50/i314  (.A1(\i50/n84 ),
    .A2(\i50/n51 ),
    .B1(\i50/n82 ),
    .B2(\i50/n52 ),
    .Y(\i50/n226 ));
 AOI22xp5_ASAP7_75t_SL \i50/i315  (.A1(\i50/n50 ),
    .A2(\i50/n55 ),
    .B1(\i50/n74 ),
    .B2(\i50/n86 ),
    .Y(\i50/n224 ));
 OAI22xp33_ASAP7_75t_SL \i50/i316  (.A1(\i50/n57 ),
    .A2(\i50/n66 ),
    .B1(\i50/n72 ),
    .B2(\i50/n78 ),
    .Y(\i50/n223 ));
 OAI22xp5_ASAP7_75t_SL \i50/i317  (.A1(\i50/n542 ),
    .A2(\i50/n82 ),
    .B1(\i50/n73 ),
    .B2(\i50/n90 ),
    .Y(\i50/n26 ));
 AOI22xp5_ASAP7_75t_SL \i50/i318  (.A1(\i50/n64 ),
    .A2(\i50/n86 ),
    .B1(\i50/n53 ),
    .B2(\i50/n65 ),
    .Y(\i50/n222 ));
 INVxp67_ASAP7_75t_SL \i50/i319  (.A(\i50/n199 ),
    .Y(\i50/n200 ));
 NAND2xp5_ASAP7_75t_SL \i50/i32  (.A(\i50/n430 ),
    .B(\i50/n449 ),
    .Y(\i50/n487 ));
 INVx1_ASAP7_75t_SL \i50/i320  (.A(\i50/n527 ),
    .Y(\i50/n198 ));
 INVxp67_ASAP7_75t_SL \i50/i321  (.A(\i50/n196 ),
    .Y(\i50/n197 ));
 INVxp67_ASAP7_75t_SL \i50/i322  (.A(\i50/n194 ),
    .Y(\i50/n195 ));
 INVxp67_ASAP7_75t_SL \i50/i323  (.A(\i50/n192 ),
    .Y(\i50/n193 ));
 INVxp67_ASAP7_75t_SL \i50/i324  (.A(\i50/n568 ),
    .Y(\i50/n190 ));
 INVxp67_ASAP7_75t_SL \i50/i325  (.A(\i50/n184 ),
    .Y(\i50/n185 ));
 INVxp67_ASAP7_75t_SL \i50/i326  (.A(\i50/n182 ),
    .Y(\i50/n183 ));
 INVxp67_ASAP7_75t_SL \i50/i327  (.A(\i50/n179 ),
    .Y(\i50/n180 ));
 INVxp67_ASAP7_75t_SL \i50/i328  (.A(\i50/n177 ),
    .Y(\i50/n178 ));
 INVxp67_ASAP7_75t_SL \i50/i329  (.A(\i50/n175 ),
    .Y(\i50/n176 ));
 NOR3x1_ASAP7_75t_SL \i50/i33  (.A(\i50/n29 ),
    .B(\i50/n570 ),
    .C(\i50/n548 ),
    .Y(\i50/n495 ));
 INVxp67_ASAP7_75t_SL \i50/i330  (.A(\i50/n173 ),
    .Y(\i50/n174 ));
 INVxp67_ASAP7_75t_SL \i50/i331  (.A(\i50/n22 ),
    .Y(\i50/n172 ));
 INVx1_ASAP7_75t_SL \i50/i332  (.A(\i50/n171 ),
    .Y(\i50/n170 ));
 NAND2xp5_ASAP7_75t_SL \i50/i333  (.A(\i50/n71 ),
    .B(\i50/n89 ),
    .Y(\i50/n205 ));
 NAND2xp5_ASAP7_75t_SL \i50/i334  (.A(\i50/n88 ),
    .B(\i50/n86 ),
    .Y(\i50/n169 ));
 NAND2xp5_ASAP7_75t_SL \i50/i335  (.A(\i50/n87 ),
    .B(\i50/n84 ),
    .Y(\i50/n168 ));
 NAND2xp5_ASAP7_75t_SL \i50/i336  (.A(\i50/n53 ),
    .B(\i50/n93 ),
    .Y(\i50/n167 ));
 NAND2xp33_ASAP7_75t_SL \i50/i337  (.A(\i50/n68 ),
    .B(\i50/n63 ),
    .Y(\i50/n166 ));
 NAND2xp5_ASAP7_75t_SL \i50/i338  (.A(\i50/n62 ),
    .B(\i50/n67 ),
    .Y(\i50/n165 ));
 NAND2xp5_ASAP7_75t_SL \i50/i339  (.A(\i50/n62 ),
    .B(\i50/n69 ),
    .Y(\i50/n204 ));
 NOR3xp33_ASAP7_75t_SL \i50/i34  (.A(\i50/n469 ),
    .B(\i50/n29 ),
    .C(\i50/n389 ),
    .Y(\i50/n485 ));
 NAND2xp5_ASAP7_75t_SL \i50/i340  (.A(\i50/n67 ),
    .B(\i50/n76 ),
    .Y(\i50/n203 ));
 NAND2xp5_ASAP7_75t_SL \i50/i341  (.A(\i50/n69 ),
    .B(\i50/n89 ),
    .Y(\i50/n164 ));
 NAND2xp5_ASAP7_75t_SL \i50/i342  (.A(\i50/n2 ),
    .B(\i50/n67 ),
    .Y(\i50/n163 ));
 NAND2xp5_ASAP7_75t_SL \i50/i343  (.A(\i50/n72 ),
    .B(\i50/n16 ),
    .Y(\i50/n162 ));
 NAND2xp5_ASAP7_75t_SL \i50/i344  (.A(\i50/n92 ),
    .B(\i50/n88 ),
    .Y(\i50/n161 ));
 NAND2xp5_ASAP7_75t_SL \i50/i345  (.A(\i50/n71 ),
    .B(\i50/n2 ),
    .Y(\i50/n160 ));
 NAND2xp5_ASAP7_75t_SL \i50/i346  (.A(\i50/n77 ),
    .B(\i50/n74 ),
    .Y(\i50/n159 ));
 NAND2xp5_ASAP7_75t_SL \i50/i347  (.A(\i50/n69 ),
    .B(\i50/n77 ),
    .Y(\i50/n158 ));
 NAND2xp5_ASAP7_75t_SL \i50/i348  (.A(\i50/n50 ),
    .B(\i50/n58 ),
    .Y(\i50/n157 ));
 NAND2xp5_ASAP7_75t_SL \i50/i349  (.A(\i50/n58 ),
    .B(\i50/n76 ),
    .Y(\i50/n156 ));
 NOR2xp67_ASAP7_75t_SL \i50/i35  (.A(\i50/n450 ),
    .B(\i50/n29 ),
    .Y(\i50/n484 ));
 NAND2xp5_ASAP7_75t_SL \i50/i350  (.A(\i50/n71 ),
    .B(\i50/n92 ),
    .Y(\i50/n155 ));
 NAND2xp5_ASAP7_75t_SL \i50/i351  (.A(\i50/n50 ),
    .B(\i50/n81 ),
    .Y(\i50/n202 ));
 AND2x2_ASAP7_75t_SL \i50/i352  (.A(\i50/n58 ),
    .B(\i50/n550 ),
    .Y(\i50/n201 ));
 AND2x2_ASAP7_75t_SL \i50/i353  (.A(\i50/n88 ),
    .B(\i50/n76 ),
    .Y(\i50/n199 ));
 NAND2xp5_ASAP7_75t_SL \i50/i354  (.A(\i50/n77 ),
    .B(\i50/n4 ),
    .Y(\i50/n25 ));
 NAND2xp5_ASAP7_75t_SL \i50/i355  (.A(\i50/n81 ),
    .B(\i50/n92 ),
    .Y(\i50/n196 ));
 NAND2xp5_ASAP7_75t_SL \i50/i356  (.A(\i50/n96 ),
    .B(\i50/n56 ),
    .Y(\i50/n194 ));
 NAND2xp5_ASAP7_75t_SL \i50/i357  (.A(\i50/n551 ),
    .B(\i50/n76 ),
    .Y(\i50/n192 ));
 AND2x2_ASAP7_75t_SL \i50/i358  (.A(\i50/n71 ),
    .B(\i50/n65 ),
    .Y(\i50/n191 ));
 NOR2xp67_ASAP7_75t_SL \i50/i359  (.A(\i50/n542 ),
    .B(\i50/n75 ),
    .Y(\i50/n24 ));
 NOR3xp33_ASAP7_75t_SL \i50/i36  (.A(\i50/n428 ),
    .B(\i50/n423 ),
    .C(\i50/n8 ),
    .Y(\i50/n483 ));
 NAND2xp5_ASAP7_75t_SL \i50/i360  (.A(\i50/n70 ),
    .B(\i50/n2 ),
    .Y(\i50/n154 ));
 NAND2xp5_ASAP7_75t_SL \i50/i361  (.A(\i50/n79 ),
    .B(\i50/n70 ),
    .Y(\i50/n189 ));
 NOR2xp33_ASAP7_75t_R \i50/i362  (.A(\i50/n73 ),
    .B(\i50/n82 ),
    .Y(\i50/n153 ));
 NAND2xp5_ASAP7_75t_SL \i50/i363  (.A(\i50/n551 ),
    .B(\i50/n62 ),
    .Y(\i50/n188 ));
 NAND2xp5_ASAP7_75t_SL \i50/i364  (.A(\i50/n65 ),
    .B(\i50/n67 ),
    .Y(\i50/n152 ));
 NOR2xp33_ASAP7_75t_SL \i50/i365  (.A(\i50/n540 ),
    .B(\i50/n82 ),
    .Y(\i50/n187 ));
 AND2x2_ASAP7_75t_SL \i50/i366  (.A(\i50/n69 ),
    .B(\i50/n2 ),
    .Y(\i50/n186 ));
 NOR2xp33_ASAP7_75t_SL \i50/i367  (.A(\i50/n17 ),
    .B(\i50/n59 ),
    .Y(\i50/n151 ));
 NAND2xp5_ASAP7_75t_SL \i50/i368  (.A(\i50/n70 ),
    .B(\i50/n56 ),
    .Y(\i50/n184 ));
 NOR2xp33_ASAP7_75t_SL \i50/i369  (.A(\i50/n551 ),
    .B(\i50/n88 ),
    .Y(\i50/n150 ));
 NAND4xp25_ASAP7_75t_SL \i50/i37  (.A(\i50/n411 ),
    .B(\i50/n405 ),
    .C(\i50/n404 ),
    .D(\i50/n437 ),
    .Y(\i50/n482 ));
 NOR2xp33_ASAP7_75t_SL \i50/i370  (.A(\i50/n540 ),
    .B(\i50/n91 ),
    .Y(\i50/n149 ));
 NAND2xp5_ASAP7_75t_SL \i50/i371  (.A(\i50/n88 ),
    .B(\i50/n2 ),
    .Y(\i50/n182 ));
 NOR2xp33_ASAP7_75t_L \i50/i372  (.A(\i50/n96 ),
    .B(\i50/n55 ),
    .Y(\i50/n181 ));
 NAND2xp5_ASAP7_75t_SL \i50/i373  (.A(\i50/n551 ),
    .B(\i50/n83 ),
    .Y(\i50/n23 ));
 NAND2xp5_ASAP7_75t_SL \i50/i374  (.A(\i50/n96 ),
    .B(\i50/n60 ),
    .Y(\i50/n179 ));
 NAND2xp5_ASAP7_75t_SL \i50/i375  (.A(\i50/n92 ),
    .B(\i50/n69 ),
    .Y(\i50/n177 ));
 NAND2xp5_ASAP7_75t_SL \i50/i376  (.A(\i50/n96 ),
    .B(\i50/n77 ),
    .Y(\i50/n175 ));
 NAND2xp5_ASAP7_75t_SL \i50/i377  (.A(\i50/n71 ),
    .B(\i50/n79 ),
    .Y(\i50/n148 ));
 NOR2xp33_ASAP7_75t_SL \i50/i378  (.A(\i50/n88 ),
    .B(\i50/n71 ),
    .Y(\i50/n173 ));
 NOR2xp33_ASAP7_75t_SL \i50/i379  (.A(\i50/n61 ),
    .B(\i50/n87 ),
    .Y(\i50/n147 ));
 NAND3xp33_ASAP7_75t_L \i50/i38  (.A(\i50/n386 ),
    .B(\i50/n405 ),
    .C(\i50/n454 ),
    .Y(\i50/n481 ));
 NOR2x1_ASAP7_75t_SL \i50/i380  (.A(\i50/n551 ),
    .B(\i50/n85 ),
    .Y(\i50/n22 ));
 OR2x2_ASAP7_75t_SL \i50/i381  (.A(\i50/n55 ),
    .B(\i50/n70 ),
    .Y(\i50/n171 ));
 INVxp67_ASAP7_75t_SL \i50/i382  (.A(\i50/n528 ),
    .Y(\i50/n146 ));
 INVxp67_ASAP7_75t_SL \i50/i383  (.A(\i50/n143 ),
    .Y(\i50/n144 ));
 INVx1_ASAP7_75t_SL \i50/i384  (.A(\i50/n141 ),
    .Y(\i50/n142 ));
 INVxp67_ASAP7_75t_SL \i50/i385  (.A(\i50/n135 ),
    .Y(\i50/n136 ));
 INVxp67_ASAP7_75t_SL \i50/i386  (.A(\i50/n133 ),
    .Y(\i50/n134 ));
 INVxp67_ASAP7_75t_SL \i50/i387  (.A(\i50/n131 ),
    .Y(\i50/n132 ));
 INVxp67_ASAP7_75t_SL \i50/i388  (.A(\i50/n129 ),
    .Y(\i50/n130 ));
 INVxp67_ASAP7_75t_SL \i50/i389  (.A(\i50/n529 ),
    .Y(\i50/n128 ));
 NAND3xp33_ASAP7_75t_SL \i50/i39  (.A(\i50/n391 ),
    .B(\i50/n439 ),
    .C(\i50/n424 ),
    .Y(\i50/n480 ));
 INVxp67_ASAP7_75t_SL \i50/i390  (.A(\i50/n126 ),
    .Y(\i50/n127 ));
 INVxp67_ASAP7_75t_SL \i50/i391  (.A(\i50/n121 ),
    .Y(\i50/n122 ));
 INVx1_ASAP7_75t_SL \i50/i392  (.A(\i50/n118 ),
    .Y(\i50/n119 ));
 INVx1_ASAP7_75t_SL \i50/i393  (.A(\i50/n18 ),
    .Y(\i50/n19 ));
 NAND2xp5_ASAP7_75t_SL \i50/i394  (.A(\i50/n85 ),
    .B(\i50/n550 ),
    .Y(\i50/n117 ));
 NAND2xp5_ASAP7_75t_SL \i50/i395  (.A(\i50/n55 ),
    .B(\i50/n79 ),
    .Y(\i50/n116 ));
 NAND2xp5_ASAP7_75t_SL \i50/i396  (.A(\i50/n64 ),
    .B(\i50/n550 ),
    .Y(\i50/n21 ));
 NAND2xp5_ASAP7_75t_SL \i50/i397  (.A(\i50/n80 ),
    .B(\i50/n73 ),
    .Y(\i50/n115 ));
 NAND2xp5_ASAP7_75t_SL \i50/i398  (.A(\i50/n64 ),
    .B(\i50/n79 ),
    .Y(\i50/n114 ));
 NAND2xp5_ASAP7_75t_SL \i50/i399  (.A(\i50/n79 ),
    .B(\i50/n53 ),
    .Y(\i50/n113 ));
 INVx2_ASAP7_75t_SL \i50/i4  (.A(\i50/n16 ),
    .Y(\i50/n4 ));
 NAND2xp5_ASAP7_75t_L \i50/i40  (.A(\i50/n438 ),
    .B(\i50/n470 ),
    .Y(\i50/n479 ));
 NAND2xp5_ASAP7_75t_SL \i50/i400  (.A(\i50/n81 ),
    .B(\i50/n65 ),
    .Y(\i50/n112 ));
 NOR2xp33_ASAP7_75t_SL \i50/i401  (.A(\i50/n92 ),
    .B(\i50/n2 ),
    .Y(\i50/n111 ));
 NAND2xp5_ASAP7_75t_SL \i50/i402  (.A(\i50/n74 ),
    .B(\i50/n60 ),
    .Y(\i50/n110 ));
 NAND2xp5_ASAP7_75t_SL \i50/i403  (.A(\i50/n53 ),
    .B(\i50/n76 ),
    .Y(\i50/n109 ));
 NAND2xp5_ASAP7_75t_L \i50/i404  (.A(\i50/n535 ),
    .B(\i50/n51 ),
    .Y(\i50/n108 ));
 NAND2xp33_ASAP7_75t_SL \i50/i405  (.A(\i50/n66 ),
    .B(\i50/n9 ),
    .Y(\i50/n107 ));
 NAND2xp5_ASAP7_75t_SL \i50/i406  (.A(\i50/n4 ),
    .B(\i50/n62 ),
    .Y(\i50/n106 ));
 NAND2xp5_ASAP7_75t_SL \i50/i407  (.A(\i50/n85 ),
    .B(\i50/n62 ),
    .Y(\i50/n105 ));
 NOR2xp33_ASAP7_75t_SL \i50/i408  (.A(\i50/n61 ),
    .B(\i50/n63 ),
    .Y(\i50/n104 ));
 NOR2xp33_ASAP7_75t_SL \i50/i409  (.A(\i50/n92 ),
    .B(\i50/n83 ),
    .Y(\i50/n145 ));
 NAND2xp5_ASAP7_75t_SL \i50/i41  (.A(\i50/n435 ),
    .B(\i50/n452 ),
    .Y(\i50/n478 ));
 NAND2xp5_ASAP7_75t_SL \i50/i410  (.A(\i50/n88 ),
    .B(\i50/n65 ),
    .Y(\i50/n143 ));
 NOR2x1_ASAP7_75t_SL \i50/i411  (.A(\i50/n76 ),
    .B(\i50/n86 ),
    .Y(\i50/n141 ));
 NAND2xp5_ASAP7_75t_SL \i50/i412  (.A(\i50/n4 ),
    .B(\i50/n83 ),
    .Y(\i50/n140 ));
 NAND2xp5_ASAP7_75t_SL \i50/i413  (.A(\i50/n81 ),
    .B(\i50/n60 ),
    .Y(\i50/n139 ));
 NAND2xp5_ASAP7_75t_SL \i50/i414  (.A(\i50/n58 ),
    .B(\i50/n62 ),
    .Y(\i50/n138 ));
 AND2x2_ASAP7_75t_SL \i50/i415  (.A(\i50/n4 ),
    .B(\i50/n56 ),
    .Y(\i50/n137 ));
 NOR2xp33_ASAP7_75t_SL \i50/i416  (.A(\i50/n76 ),
    .B(\i50/n62 ),
    .Y(\i50/n103 ));
 NAND2xp5_ASAP7_75t_SL \i50/i417  (.A(\i50/n85 ),
    .B(\i50/n92 ),
    .Y(\i50/n135 ));
 NAND2xp5_ASAP7_75t_SL \i50/i418  (.A(\i50/n85 ),
    .B(\i50/n56 ),
    .Y(\i50/n133 ));
 NOR2xp67_ASAP7_75t_SL \i50/i419  (.A(\i50/n57 ),
    .B(\i50/n90 ),
    .Y(\i50/n131 ));
 NOR2x1_ASAP7_75t_SL \i50/i42  (.A(\i50/n460 ),
    .B(\i50/n451 ),
    .Y(\i50/n486 ));
 NAND2xp5_ASAP7_75t_SL \i50/i420  (.A(\i50/n53 ),
    .B(\i50/n56 ),
    .Y(\i50/n129 ));
 NOR2xp33_ASAP7_75t_SL \i50/i421  (.A(\i50/n51 ),
    .B(\i50/n63 ),
    .Y(\i50/n126 ));
 NAND2xp5_ASAP7_75t_SL \i50/i422  (.A(\i50/n55 ),
    .B(\i50/n83 ),
    .Y(\i50/n20 ));
 NAND2xp5_ASAP7_75t_SL \i50/i423  (.A(\i50/n55 ),
    .B(\i50/n86 ),
    .Y(\i50/n125 ));
 NAND2xp5_ASAP7_75t_SL \i50/i424  (.A(\i50/n2 ),
    .B(\i50/n64 ),
    .Y(\i50/n124 ));
 NAND2xp33_ASAP7_75t_L \i50/i425  (.A(\i50/n2 ),
    .B(\i50/n81 ),
    .Y(\i50/n102 ));
 NOR2xp33_ASAP7_75t_SL \i50/i426  (.A(\i50/n66 ),
    .B(\i50/n52 ),
    .Y(\i50/n101 ));
 NOR2xp67_ASAP7_75t_SL \i50/i427  (.A(\i50/n563 ),
    .B(\i50/n550 ),
    .Y(\i50/n123 ));
 NAND2xp5_ASAP7_75t_SL \i50/i428  (.A(\i50/n4 ),
    .B(\i50/n86 ),
    .Y(\i50/n100 ));
 NAND2xp5_ASAP7_75t_SL \i50/i429  (.A(\i50/n64 ),
    .B(\i50/n60 ),
    .Y(\i50/n121 ));
 NAND2xp33_ASAP7_75t_L \i50/i43  (.A(\i50/n441 ),
    .B(\i50/n413 ),
    .Y(\i50/n475 ));
 NAND2xp5_ASAP7_75t_SL \i50/i430  (.A(\i50/n81 ),
    .B(\i50/n86 ),
    .Y(\i50/n120 ));
 NAND2xp5_ASAP7_75t_SL \i50/i431  (.A(\i50/n64 ),
    .B(\i50/n83 ),
    .Y(\i50/n99 ));
 NOR2xp33_ASAP7_75t_SL \i50/i432  (.A(\i50/n521 ),
    .B(\i50/n59 ),
    .Y(\i50/n98 ));
 NOR2xp33_ASAP7_75t_SL \i50/i433  (.A(\i50/n521 ),
    .B(\i50/n61 ),
    .Y(\i50/n97 ));
 NAND2xp5_ASAP7_75t_SL \i50/i434  (.A(\i50/n64 ),
    .B(\i50/n89 ),
    .Y(\i50/n118 ));
 NAND2xp5_ASAP7_75t_SL \i50/i435  (.A(\i50/n4 ),
    .B(\i50/n60 ),
    .Y(\i50/n18 ));
 INVx1_ASAP7_75t_SL \i50/i436  (.A(\i50/n96 ),
    .Y(\i50/n95 ));
 INVx3_ASAP7_75t_SL \i50/i437  (.A(\i50/n94 ),
    .Y(\i50/n93 ));
 INVx4_ASAP7_75t_SL \i50/i438  (.A(\i50/n92 ),
    .Y(\i50/n91 ));
 INVx3_ASAP7_75t_SL \i50/i439  (.A(\i50/n90 ),
    .Y(\i50/n89 ));
 NAND2xp33_ASAP7_75t_SL \i50/i44  (.A(\i50/n438 ),
    .B(\i50/n418 ),
    .Y(\i50/n474 ));
 INVx2_ASAP7_75t_SL \i50/i440  (.A(\i50/n88 ),
    .Y(\i50/n87 ));
 INVx2_ASAP7_75t_SL \i50/i441  (.A(\i50/n85 ),
    .Y(\i50/n84 ));
 INVx4_ASAP7_75t_SL \i50/i442  (.A(\i50/n83 ),
    .Y(\i50/n82 ));
 INVx2_ASAP7_75t_SL \i50/i443  (.A(\i50/n81 ),
    .Y(\i50/n80 ));
 INVx2_ASAP7_75t_SL \i50/i444  (.A(\i50/n550 ),
    .Y(\i50/n78 ));
 INVx3_ASAP7_75t_SL \i50/i445  (.A(\i50/n76 ),
    .Y(\i50/n75 ));
 INVx3_ASAP7_75t_SL \i50/i446  (.A(\i50/n74 ),
    .Y(\i50/n73 ));
 INVx3_ASAP7_75t_SL \i50/i447  (.A(\i50/n72 ),
    .Y(\i50/n71 ));
 AND2x4_ASAP7_75t_SL \i50/i448  (.A(\i50/n44 ),
    .B(\i50/n517 ),
    .Y(\i50/n96 ));
 OR2x2_ASAP7_75t_SL \i50/i449  (.A(\i50/n35 ),
    .B(\i50/n6 ),
    .Y(\i50/n94 ));
 NOR2xp33_ASAP7_75t_SL \i50/i45  (.A(\i50/n417 ),
    .B(\i50/n443 ),
    .Y(\i50/n473 ));
 AND2x4_ASAP7_75t_SL \i50/i450  (.A(\i50/n40 ),
    .B(\i50/n3 ),
    .Y(\i50/n92 ));
 OR2x6_ASAP7_75t_SL \i50/i451  (.A(\i50/n38 ),
    .B(\i50/n49 ),
    .Y(\i50/n90 ));
 AND2x4_ASAP7_75t_SL \i50/i452  (.A(\i50/n34 ),
    .B(\i50/n47 ),
    .Y(\i50/n88 ));
 AND2x4_ASAP7_75t_SL \i50/i453  (.A(\i50/n37 ),
    .B(\i50/n508 ),
    .Y(\i50/n86 ));
 AND2x4_ASAP7_75t_SL \i50/i454  (.A(\i50/n34 ),
    .B(\i50/n44 ),
    .Y(\i50/n85 ));
 AND2x4_ASAP7_75t_SL \i50/i455  (.A(\i50/n48 ),
    .B(\i50/n36 ),
    .Y(\i50/n83 ));
 AND2x4_ASAP7_75t_SL \i50/i456  (.A(\i50/n34 ),
    .B(\i50/n43 ),
    .Y(\i50/n81 ));
 AND2x4_ASAP7_75t_SL \i50/i457  (.A(\i50/n37 ),
    .B(\i50/n39 ),
    .Y(\i50/n79 ));
 AND2x4_ASAP7_75t_SL \i50/i458  (.A(\i50/n40 ),
    .B(\i50/n37 ),
    .Y(\i50/n77 ));
 AND2x4_ASAP7_75t_SL \i50/i459  (.A(\i50/n37 ),
    .B(\i50/n36 ),
    .Y(\i50/n76 ));
 NAND3xp33_ASAP7_75t_SL \i50/i46  (.A(\i50/n408 ),
    .B(\i50/n415 ),
    .C(\i50/n381 ),
    .Y(\i50/n472 ));
 AND2x4_ASAP7_75t_SL \i50/i460  (.A(\i50/n44 ),
    .B(\i50/n42 ),
    .Y(\i50/n74 ));
 OR2x6_ASAP7_75t_SL \i50/i461  (.A(\i50/n45 ),
    .B(\i50/n33 ),
    .Y(\i50/n72 ));
 INVx3_ASAP7_75t_SL \i50/i462  (.A(\i50/n69 ),
    .Y(\i50/n17 ));
 INVx3_ASAP7_75t_SL \i50/i463  (.A(\i50/n551 ),
    .Y(\i50/n68 ));
 INVx4_ASAP7_75t_SL \i50/i464  (.A(\i50/n66 ),
    .Y(\i50/n65 ));
 INVx4_ASAP7_75t_SL \i50/i465  (.A(\i50/n64 ),
    .Y(\i50/n63 ));
 INVx2_ASAP7_75t_SL \i50/i466  (.A(\i50/n62 ),
    .Y(\i50/n61 ));
 INVx4_ASAP7_75t_SL \i50/i467  (.A(\i50/n58 ),
    .Y(\i50/n57 ));
 INVx3_ASAP7_75t_SL \i50/i468  (.A(\i50/n55 ),
    .Y(\i50/n54 ));
 INVx3_ASAP7_75t_SL \i50/i469  (.A(\i50/n53 ),
    .Y(\i50/n52 ));
 NOR2x1_ASAP7_75t_SL \i50/i47  (.A(\i50/n365 ),
    .B(\i50/n426 ),
    .Y(\i50/n471 ));
 INVx3_ASAP7_75t_SL \i50/i470  (.A(\i50/n51 ),
    .Y(\i50/n50 ));
 AND2x4_ASAP7_75t_SL \i50/i471  (.A(\i50/n44 ),
    .B(\i50/n11 ),
    .Y(\i50/n70 ));
 AND2x4_ASAP7_75t_SL \i50/i472  (.A(\i50/n517 ),
    .B(\i50/n47 ),
    .Y(\i50/n69 ));
 OR2x2_ASAP7_75t_SL \i50/i473  (.A(\i50/n10 ),
    .B(\i50/n46 ),
    .Y(\i50/n16 ));
 AND2x4_ASAP7_75t_SL \i50/i474  (.A(\i50/n43 ),
    .B(\i50/n517 ),
    .Y(\i50/n67 ));
 NAND2x1p5_ASAP7_75t_SL \i50/i475  (.A(\i50/n40 ),
    .B(\i50/n48 ),
    .Y(\i50/n66 ));
 NAND2x1p5_ASAP7_75t_SL \i50/i476  (.A(\i50/n3 ),
    .B(\i50/n39 ),
    .Y(\i50/n9 ));
 AND2x4_ASAP7_75t_SL \i50/i477  (.A(\i50/n43 ),
    .B(\i50/n11 ),
    .Y(\i50/n64 ));
 AND2x4_ASAP7_75t_SL \i50/i478  (.A(\i50/n39 ),
    .B(\i50/n15 ),
    .Y(\i50/n62 ));
 AND2x4_ASAP7_75t_SL \i50/i479  (.A(\i50/n36 ),
    .B(\i50/n15 ),
    .Y(\i50/n60 ));
 NOR2xp33_ASAP7_75t_SL \i50/i48  (.A(\i50/n433 ),
    .B(\i50/n347 ),
    .Y(\i50/n470 ));
 AND2x4_ASAP7_75t_SL \i50/i480  (.A(\i50/n5 ),
    .B(\i50/n11 ),
    .Y(\i50/n58 ));
 AND2x4_ASAP7_75t_SL \i50/i481  (.A(\i50/n3 ),
    .B(\i50/n508 ),
    .Y(\i50/n56 ));
 AND2x4_ASAP7_75t_SL \i50/i482  (.A(\i50/n43 ),
    .B(\i50/n42 ),
    .Y(\i50/n55 ));
 AND2x4_ASAP7_75t_SL \i50/i483  (.A(\i50/n47 ),
    .B(\i50/n42 ),
    .Y(\i50/n53 ));
 OR2x6_ASAP7_75t_SL \i50/i484  (.A(\i50/n32 ),
    .B(\i50/n41 ),
    .Y(\i50/n51 ));
 INVx2_ASAP7_75t_SL \i50/i485  (.A(\i50/n48 ),
    .Y(\i50/n49 ));
 INVx2_ASAP7_75t_SL \i50/i486  (.A(\i50/n46 ),
    .Y(\i50/n47 ));
 NAND2xp5_ASAP7_75t_SL \i50/i487  (.A(\i50/n12 ),
    .B(\i50/n0 ),
    .Y(\i50/n41 ));
 AND2x2_ASAP7_75t_SL \i50/i488  (.A(\i50/n12 ),
    .B(\i50/n0 ),
    .Y(\i50/n48 ));
 NAND2x1_ASAP7_75t_L \i50/i489  (.A(\i50/n507 ),
    .B(n21[5]),
    .Y(\i50/n46 ));
 NAND2xp5_ASAP7_75t_SL \i50/i49  (.A(\i50/n441 ),
    .B(\i50/n436 ),
    .Y(\i50/n469 ));
 NAND2x1p5_ASAP7_75t_SL \i50/i490  (.A(n21[4]),
    .B(n21[5]),
    .Y(\i50/n45 ));
 AND2x2_ASAP7_75t_SL \i50/i491  (.A(\i50/n30 ),
    .B(\i50/n507 ),
    .Y(\i50/n44 ));
 AND2x2_ASAP7_75t_SL \i50/i492  (.A(n21[4]),
    .B(\i50/n30 ),
    .Y(\i50/n43 ));
 AND2x4_ASAP7_75t_SL \i50/i493  (.A(n21[7]),
    .B(\i50/n14 ),
    .Y(\i50/n42 ));
 INVx1_ASAP7_75t_SL \i50/i494  (.A(\i50/n39 ),
    .Y(\i50/n38 ));
 INVx2_ASAP7_75t_SL \i50/i495  (.A(\i50/n558 ),
    .Y(\i50/n36 ));
 INVx2_ASAP7_75t_SL \i50/i496  (.A(\i50/n34 ),
    .Y(\i50/n33 ));
 NAND2xp5_ASAP7_75t_SL \i50/i497  (.A(\i50/n31 ),
    .B(\i50/n1 ),
    .Y(\i50/n32 ));
 AND2x2_ASAP7_75t_SL \i50/i498  (.A(n21[0]),
    .B(n21[1]),
    .Y(\i50/n40 ));
 AND2x4_ASAP7_75t_SL \i50/i499  (.A(n21[0]),
    .B(\i50/n31 ),
    .Y(\i50/n39 ));
 INVx2_ASAP7_75t_SL \i50/i5  (.A(\i50/n45 ),
    .Y(\i50/n5 ));
 NOR2x1_ASAP7_75t_SL \i50/i50  (.A(\i50/n351 ),
    .B(\i50/n443 ),
    .Y(\i50/n468 ));
 AND2x4_ASAP7_75t_SL \i50/i500  (.A(n21[3]),
    .B(n21[2]),
    .Y(\i50/n37 ));
 NAND2x1_ASAP7_75t_SL \i50/i501  (.A(n21[3]),
    .B(\i50/n0 ),
    .Y(\i50/n35 ));
 AND2x2_ASAP7_75t_SL \i50/i502  (.A(n21[7]),
    .B(n21[6]),
    .Y(\i50/n34 ));
 INVx1_ASAP7_75t_SL \i50/i503  (.A(n21[1]),
    .Y(\i50/n31 ));
 INVx3_ASAP7_75t_SL \i50/i504  (.A(n21[5]),
    .Y(\i50/n30 ));
 INVx2_ASAP7_75t_SL \i50/i505  (.A(\i50/n35 ),
    .Y(\i50/n15 ));
 INVx2_ASAP7_75t_SL \i50/i506  (.A(n21[6]),
    .Y(\i50/n14 ));
 INVx2_ASAP7_75t_SL \i50/i507  (.A(n21[7]),
    .Y(\i50/n13 ));
 INVx2_ASAP7_75t_SL \i50/i508  (.A(n21[3]),
    .Y(\i50/n12 ));
 INVx1_ASAP7_75t_SL \i50/i509  (.A(\i50/n439 ),
    .Y(\i50/n8 ));
 NOR2x1_ASAP7_75t_SL \i50/i51  (.A(\i50/n416 ),
    .B(\i50/n427 ),
    .Y(\i50/n467 ));
 AND2x2_ASAP7_75t_SL \i50/i510  (.A(\i50/n13 ),
    .B(n21[6]),
    .Y(\i50/n11 ));
 NAND2xp5_ASAP7_75t_SL \i50/i511  (.A(\i50/n13 ),
    .B(n21[6]),
    .Y(\i50/n10 ));
 OR2x2_ASAP7_75t_SL \i50/i512  (.A(\i50/n137 ),
    .B(\i50/n567 ),
    .Y(\i50/n7 ));
 OR2x2_ASAP7_75t_SL \i50/i513  (.A(n21[0]),
    .B(n21[1]),
    .Y(\i50/n6 ));
 INVx2_ASAP7_75t_SL \i50/i514  (.A(n21[4]),
    .Y(\i50/n507 ));
 INVx2_ASAP7_75t_SL \i50/i515  (.A(\i50/n6 ),
    .Y(\i50/n508 ));
 NAND2x1_ASAP7_75t_SL \i50/i516  (.A(\i50/n3 ),
    .B(\i50/n508 ),
    .Y(\i50/n509 ));
 OAI21xp5_ASAP7_75t_SL \i50/i517  (.A1(\i50/n80 ),
    .A2(\i50/n509 ),
    .B(\i50/n114 ),
    .Y(\i50/n510 ));
 OAI222xp33_ASAP7_75t_SL \i50/i518  (.A1(\i50/n90 ),
    .A2(\i50/n52 ),
    .B1(\i50/n509 ),
    .B2(\i50/n17 ),
    .C1(\i50/n541 ),
    .C2(\i50/n72 ),
    .Y(\i50/n511 ));
 OAI22xp33_ASAP7_75t_SL \i50/i519  (.A1(\i50/n509 ),
    .A2(\i50/n540 ),
    .B1(\i50/n59 ),
    .B2(\i50/n57 ),
    .Y(\i50/n512 ));
 NAND2xp5_ASAP7_75t_SL \i50/i52  (.A(\i50/n538 ),
    .B(\i50/n421 ),
    .Y(\i50/n466 ));
 A2O1A1Ixp33_ASAP7_75t_R \i50/i520  (.A1(\i50/n539 ),
    .A2(\i50/n509 ),
    .B(\i50/n87 ),
    .C(\i50/n241 ),
    .Y(\i50/n513 ));
 OAI22xp5_ASAP7_75t_SL \i50/i521  (.A1(\i50/n68 ),
    .A2(\i50/n509 ),
    .B1(\i50/n72 ),
    .B2(\i50/n82 ),
    .Y(\i50/n514 ));
 NAND2xp33_ASAP7_75t_L \i50/i522  (.A(\i50/n509 ),
    .B(\i50/n78 ),
    .Y(\i50/n515 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i50/i523  (.A1(\i50/n90 ),
    .A2(\i50/n509 ),
    .B(\i50/n73 ),
    .C(\i50/n125 ),
    .Y(\i50/n516 ));
 AND2x2_ASAP7_75t_SL \i50/i524  (.A(\i50/n13 ),
    .B(\i50/n14 ),
    .Y(\i50/n517 ));
 NAND2xp5_ASAP7_75t_SL \i50/i525  (.A(\i50/n2 ),
    .B(\i50/n518 ),
    .Y(\i50/n519 ));
 AND2x4_ASAP7_75t_SL \i50/i526  (.A(\i50/n517 ),
    .B(\i50/n5 ),
    .Y(\i50/n518 ));
 AOI22xp5_ASAP7_75t_SL \i50/i527  (.A1(\i50/n92 ),
    .A2(\i50/n518 ),
    .B1(\i50/n85 ),
    .B2(\i50/n77 ),
    .Y(\i50/n520 ));
 INVx2_ASAP7_75t_SL \i50/i528  (.A(\i50/n518 ),
    .Y(\i50/n521 ));
 AOI22xp33_ASAP7_75t_SL \i50/i529  (.A1(\i50/n70 ),
    .A2(\i50/n65 ),
    .B1(\i50/n518 ),
    .B2(\i50/n62 ),
    .Y(\i50/n522 ));
 NOR5xp2_ASAP7_75t_SL \i50/i53  (.A(\i50/n307 ),
    .B(\i50/n564 ),
    .C(\i50/n320 ),
    .D(\i50/n28 ),
    .E(\i50/n287 ),
    .Y(\i50/n465 ));
 AOI22xp5_ASAP7_75t_SL \i50/i530  (.A1(\i50/n518 ),
    .A2(\i50/n83 ),
    .B1(\i50/n81 ),
    .B2(\i50/n2 ),
    .Y(\i50/n523 ));
 AOI22xp5_ASAP7_75t_R \i50/i531  (.A1(\i50/n518 ),
    .A2(\i50/n89 ),
    .B1(\i50/n88 ),
    .B2(\i50/n60 ),
    .Y(\i50/n524 ));
 AOI22xp33_ASAP7_75t_SL \i50/i532  (.A1(\i50/n50 ),
    .A2(\i50/n53 ),
    .B1(\i50/n518 ),
    .B2(\i50/n550 ),
    .Y(\i50/n525 ));
 AOI22xp5_ASAP7_75t_SL \i50/i533  (.A1(\i50/n518 ),
    .A2(\i50/n56 ),
    .B1(\i50/n551 ),
    .B2(\i50/n77 ),
    .Y(\i50/n526 ));
 AND2x2_ASAP7_75t_SL \i50/i534  (.A(\i50/n518 ),
    .B(\i50/n77 ),
    .Y(\i50/n527 ));
 NAND2xp5_ASAP7_75t_SL \i50/i535  (.A(\i50/n518 ),
    .B(\i50/n563 ),
    .Y(\i50/n528 ));
 NAND2xp5_ASAP7_75t_SL \i50/i536  (.A(\i50/n50 ),
    .B(\i50/n518 ),
    .Y(\i50/n529 ));
 AND2x2_ASAP7_75t_SL \i50/i537  (.A(\i50/n518 ),
    .B(\i50/n86 ),
    .Y(\i50/n530 ));
 AND2x2_ASAP7_75t_SL \i50/i538  (.A(\i50/n518 ),
    .B(\i50/n65 ),
    .Y(\i50/n531 ));
 NAND2xp5_ASAP7_75t_SL \i50/i539  (.A(\i50/n518 ),
    .B(\i50/n79 ),
    .Y(\i50/n532 ));
 NOR2x1_ASAP7_75t_SL \i50/i54  (.A(\i50/n8 ),
    .B(\i50/n428 ),
    .Y(\i50/n464 ));
 INVx1_ASAP7_75t_SL \i50/i540  (.A(\i50/n309 ),
    .Y(\i50/n533 ));
 OA21x2_ASAP7_75t_SL \i50/i541  (.A1(\i50/n57 ),
    .A2(\i50/n559 ),
    .B(\i50/n21 ),
    .Y(\i50/n534 ));
 INVx2_ASAP7_75t_SL \i50/i542  (.A(\i50/n60 ),
    .Y(\i50/n59 ));
 NAND2x1_ASAP7_75t_SL \i50/i543  (.A(\i50/n37 ),
    .B(\i50/n508 ),
    .Y(\i50/n535 ));
 OAI21xp33_ASAP7_75t_L \i50/i544  (.A1(\i50/n536 ),
    .A2(\i50/n550 ),
    .B(\i50/n85 ),
    .Y(\i50/n537 ));
 NAND2xp5_ASAP7_75t_SL \i50/i545  (.A(\i50/n59 ),
    .B(\i50/n535 ),
    .Y(\i50/n536 ));
 AOI211xp5_ASAP7_75t_SL \i50/i546  (.A1(\i50/n536 ),
    .A2(\i50/n58 ),
    .B(\i50/n328 ),
    .C(\i50/n265 ),
    .Y(\i50/n538 ));
 INVx3_ASAP7_75t_SL \i50/i547  (.A(\i50/n79 ),
    .Y(\i50/n539 ));
 INVx3_ASAP7_75t_SL \i50/i548  (.A(\i50/n67 ),
    .Y(\i50/n540 ));
 INVx2_ASAP7_75t_SL \i50/i549  (.A(\i50/n77 ),
    .Y(\i50/n541 ));
 NAND2x1_ASAP7_75t_SL \i50/i55  (.A(\i50/n425 ),
    .B(\i50/n406 ),
    .Y(\i50/n477 ));
 INVx3_ASAP7_75t_SL \i50/i550  (.A(\i50/n70 ),
    .Y(\i50/n542 ));
 AO21x2_ASAP7_75t_SL \i50/i551  (.A1(\i50/n85 ),
    .A2(\i50/n2 ),
    .B(\i50/n543 ),
    .Y(\i50/n544 ));
 OAI22xp5_ASAP7_75t_SL \i50/i552  (.A1(\i50/n539 ),
    .A2(\i50/n540 ),
    .B1(\i50/n541 ),
    .B2(\i50/n542 ),
    .Y(\i50/n543 ));
 AND2x2_ASAP7_75t_SL \i50/i553  (.A(\i50/n4 ),
    .B(\i50/n79 ),
    .Y(\i50/n545 ));
 NAND2xp5_ASAP7_75t_SL \i50/i554  (.A(\i50/n292 ),
    .B(\i50/n547 ),
    .Y(\i50/n548 ));
 NOR2xp67_ASAP7_75t_SL \i50/i555  (.A(\i50/n545 ),
    .B(\i50/n546 ),
    .Y(\i50/n547 ));
 OAI22xp5_ASAP7_75t_SL \i50/i556  (.A1(\i50/n94 ),
    .A2(\i50/n57 ),
    .B1(\i50/n54 ),
    .B2(\i50/n59 ),
    .Y(\i50/n546 ));
 NAND5xp2_ASAP7_75t_SL \i50/i557  (.A(\i50/n547 ),
    .B(\i50/n565 ),
    .C(\i50/n526 ),
    .D(\i50/n99 ),
    .E(\i50/n200 ),
    .Y(\i50/n549 ));
 AND2x4_ASAP7_75t_SL \i50/i558  (.A(\i50/n40 ),
    .B(\i50/n15 ),
    .Y(\i50/n550 ));
 AND2x4_ASAP7_75t_SL \i50/i559  (.A(\i50/n5 ),
    .B(\i50/n42 ),
    .Y(\i50/n551 ));
 NOR2x1_ASAP7_75t_SL \i50/i56  (.A(\i50/n444 ),
    .B(\i50/n427 ),
    .Y(\i50/n463 ));
 OAI22xp5_ASAP7_75t_SL \i50/i560  (.A1(\i50/n63 ),
    .A2(\i50/n94 ),
    .B1(\i50/n72 ),
    .B2(\i50/n91 ),
    .Y(\i50/n552 ));
 NAND2xp5_ASAP7_75t_SL \i50/i561  (.A(\i50/n296 ),
    .B(\i50/n553 ),
    .Y(\i50/n554 ));
 AOI21xp33_ASAP7_75t_SL \i50/i562  (.A1(\i50/n550 ),
    .A2(\i50/n551 ),
    .B(\i50/n552 ),
    .Y(\i50/n553 ));
 INVxp67_ASAP7_75t_SL \i50/i563  (.A(\i50/n553 ),
    .Y(\i50/n555 ));
 AOI31xp33_ASAP7_75t_SL \i50/i564  (.A1(\i50/n57 ),
    .A2(\i50/n84 ),
    .A3(\i50/n73 ),
    .B(\i50/n559 ),
    .Y(\i50/n556 ));
 OR2x2_ASAP7_75t_SL \i50/i565  (.A(\i50/n0 ),
    .B(n21[3]),
    .Y(\i50/n557 ));
 NAND2xp5_ASAP7_75t_SL \i50/i566  (.A(\i50/n1 ),
    .B(n21[1]),
    .Y(\i50/n558 ));
 OAI221xp5_ASAP7_75t_SL \i50/i567  (.A1(\i50/n63 ),
    .A2(\i50/n509 ),
    .B1(\i50/n52 ),
    .B2(\i50/n559 ),
    .C(\i50/n529 ),
    .Y(\i50/n560 ));
 OR2x2_ASAP7_75t_SL \i50/i568  (.A(\i50/n557 ),
    .B(\i50/n558 ),
    .Y(\i50/n559 ));
 OAI22xp5_ASAP7_75t_SL \i50/i569  (.A1(\i50/n57 ),
    .A2(\i50/n509 ),
    .B1(\i50/n559 ),
    .B2(\i50/n54 ),
    .Y(\i50/n561 ));
 NOR2x1_ASAP7_75t_SL \i50/i57  (.A(\i50/n364 ),
    .B(\i50/n426 ),
    .Y(\i50/n476 ));
 OAI21xp5_ASAP7_75t_SL \i50/i570  (.A1(\i50/n80 ),
    .A2(\i50/n559 ),
    .B(\i50/n138 ),
    .Y(\i50/n562 ));
 INVx3_ASAP7_75t_SL \i50/i571  (.A(\i50/n559 ),
    .Y(\i50/n563 ));
 OAI221xp5_ASAP7_75t_SL \i50/i572  (.A1(\i50/n61 ),
    .A2(\i50/n542 ),
    .B1(\i50/n57 ),
    .B2(\i50/n559 ),
    .C(\i50/n21 ),
    .Y(\i50/n564 ));
 AO21x1_ASAP7_75t_SL \i50/i573  (.A1(\i50/n559 ),
    .A2(\i50/n169 ),
    .B(\i50/n150 ),
    .Y(\i50/n565 ));
 OAI22xp33_ASAP7_75t_SL \i50/i574  (.A1(\i50/n54 ),
    .A2(\i50/n94 ),
    .B1(\i50/n559 ),
    .B2(\i50/n540 ),
    .Y(\i50/n566 ));
 OAI22xp5_ASAP7_75t_SL \i50/i575  (.A1(\i50/n57 ),
    .A2(\i50/n82 ),
    .B1(\i50/n72 ),
    .B2(\i50/n559 ),
    .Y(\i50/n567 ));
 NOR2xp33_ASAP7_75t_SL \i50/i576  (.A(\i50/n559 ),
    .B(\i50/n542 ),
    .Y(\i50/n568 ));
 NOR2xp33_ASAP7_75t_SL \i50/i577  (.A(\i50/n559 ),
    .B(\i50/n54 ),
    .Y(\i50/n569 ));
 INVx1_ASAP7_75t_SL \i50/i578  (.A(\i50/n445 ),
    .Y(\i50/n570 ));
 AND4x1_ASAP7_75t_SL \i50/i579  (.A(\i50/n306 ),
    .B(\i50/n349 ),
    .C(\i50/n576 ),
    .D(\i50/n282 ),
    .Y(\i50/n571 ));
 INVxp67_ASAP7_75t_SL \i50/i58  (.A(\i50/n461 ),
    .Y(\i50/n462 ));
 OR4x1_ASAP7_75t_SL \i50/i580  (.A(\i50/n262 ),
    .B(\i50/n276 ),
    .C(\i50/n272 ),
    .D(\i50/n267 ),
    .Y(\i50/n572 ));
 AO221x1_ASAP7_75t_SL \i50/i581  (.A1(\i50/n70 ),
    .A2(\i50/n550 ),
    .B1(\i50/n4 ),
    .B2(\i50/n563 ),
    .C(\i50/n279 ),
    .Y(\i50/n573 ));
 NOR3xp33_ASAP7_75t_SL \i50/i582  (.A(\i50/n574 ),
    .B(\i50/n339 ),
    .C(\i50/n543 ),
    .Y(\i50/n575 ));
 OAI21xp5_ASAP7_75t_SL \i50/i583  (.A1(\i50/n72 ),
    .A2(\i50/n535 ),
    .B(\i50/n124 ),
    .Y(\i50/n574 ));
 AOI21xp5_ASAP7_75t_SL \i50/i584  (.A1(\i50/n58 ),
    .A2(\i50/n77 ),
    .B(\i50/n561 ),
    .Y(\i50/n576 ));
 AND2x2_ASAP7_75t_SL \i50/i585  (.A(\i50/n577 ),
    .B(\i50/n440 ),
    .Y(\i50/n578 ));
 AOI21xp33_ASAP7_75t_SL \i50/i586  (.A1(\i50/n50 ),
    .A2(\i50/n74 ),
    .B(\i50/n530 ),
    .Y(\i50/n577 ));
 NAND2xp33_ASAP7_75t_SL \i50/i587  (.A(\i50/n579 ),
    .B(\i50/n309 ),
    .Y(\i50/n580 ));
 OAI21xp5_ASAP7_75t_SL \i50/i588  (.A1(\i50/n2 ),
    .A2(\i50/n550 ),
    .B(\i50/n53 ),
    .Y(\i50/n579 ));
 INVxp67_ASAP7_75t_SL \i50/i59  (.A(\i50/n457 ),
    .Y(\i50/n458 ));
 NOR2x1p5_ASAP7_75t_SL \i50/i6  (.A(\i50/n502 ),
    .B(\i50/n501 ),
    .Y(n20[4]));
 AND5x1_ASAP7_75t_SL \i50/i60  (.A(\i50/n376 ),
    .B(\i50/n576 ),
    .C(\i50/n369 ),
    .D(\i50/n295 ),
    .E(\i50/n270 ),
    .Y(\i50/n456 ));
 NOR3xp33_ASAP7_75t_SL \i50/i61  (.A(\i50/n388 ),
    .B(\i50/n368 ),
    .C(\i50/n555 ),
    .Y(\i50/n455 ));
 NOR3xp33_ASAP7_75t_SL \i50/i62  (.A(\i50/n414 ),
    .B(\i50/n352 ),
    .C(\i50/n305 ),
    .Y(\i50/n454 ));
 AND5x1_ASAP7_75t_SL \i50/i63  (.A(\i50/n343 ),
    .B(\i50/n355 ),
    .C(\i50/n337 ),
    .D(\i50/n346 ),
    .E(\i50/n278 ),
    .Y(\i50/n453 ));
 NOR2xp33_ASAP7_75t_SL \i50/i64  (.A(\i50/n549 ),
    .B(\i50/n419 ),
    .Y(\i50/n452 ));
 NAND4xp25_ASAP7_75t_SL \i50/i65  (.A(\i50/n397 ),
    .B(\i50/n405 ),
    .C(\i50/n410 ),
    .D(\i50/n393 ),
    .Y(\i50/n451 ));
 NAND5xp2_ASAP7_75t_SL \i50/i66  (.A(\i50/n375 ),
    .B(\i50/n335 ),
    .C(\i50/n238 ),
    .D(\i50/n225 ),
    .E(\i50/n315 ),
    .Y(\i50/n450 ));
 NOR4xp25_ASAP7_75t_SL \i50/i67  (.A(\i50/n366 ),
    .B(\i50/n564 ),
    .C(\i50/n321 ),
    .D(\i50/n513 ),
    .Y(\i50/n449 ));
 NAND4xp25_ASAP7_75t_SL \i50/i68  (.A(\i50/n384 ),
    .B(\i50/n399 ),
    .C(\i50/n402 ),
    .D(\i50/n404 ),
    .Y(\i50/n448 ));
 NAND4xp25_ASAP7_75t_SL \i50/i69  (.A(\i50/n412 ),
    .B(\i50/n410 ),
    .C(\i50/n534 ),
    .D(\i50/n269 ),
    .Y(\i50/n447 ));
 NOR2x1p5_ASAP7_75t_SL \i50/i7  (.A(\i50/n497 ),
    .B(\i50/n503 ),
    .Y(n20[3]));
 NAND3xp33_ASAP7_75t_SL \i50/i70  (.A(\i50/n404 ),
    .B(\i50/n374 ),
    .C(\i50/n20 ),
    .Y(\i50/n461 ));
 NAND4xp75_ASAP7_75t_SL \i50/i71  (.A(\i50/n311 ),
    .B(\i50/n286 ),
    .C(\i50/n363 ),
    .D(\i50/n25 ),
    .Y(\i50/n460 ));
 NAND2xp33_ASAP7_75t_L \i50/i72  (.A(\i50/n383 ),
    .B(\i50/n445 ),
    .Y(\i50/n446 ));
 AND2x2_ASAP7_75t_SL \i50/i73  (.A(\i50/n386 ),
    .B(\i50/n434 ),
    .Y(\i50/n459 ));
 NAND2x1p5_ASAP7_75t_SL \i50/i74  (.A(\i50/n442 ),
    .B(\i50/n398 ),
    .Y(\i50/n457 ));
 NOR5xp2_ASAP7_75t_SL \i50/i75  (.A(\i50/n330 ),
    .B(\i50/n304 ),
    .C(\i50/n231 ),
    .D(\i50/n527 ),
    .E(\i50/n569 ),
    .Y(\i50/n437 ));
 NOR3xp33_ASAP7_75t_SL \i50/i76  (.A(\i50/n409 ),
    .B(\i50/n325 ),
    .C(\i50/n318 ),
    .Y(\i50/n436 ));
 NOR2xp33_ASAP7_75t_SL \i50/i77  (.A(\i50/n580 ),
    .B(\i50/n385 ),
    .Y(\i50/n435 ));
 NOR2xp33_ASAP7_75t_SL \i50/i78  (.A(\i50/n407 ),
    .B(\i50/n357 ),
    .Y(\i50/n434 ));
 NOR2x1_ASAP7_75t_SL \i50/i79  (.A(\i50/n370 ),
    .B(\i50/n344 ),
    .Y(\i50/n445 ));
 AND5x2_ASAP7_75t_SL \i50/i8  (.A(\i50/n495 ),
    .B(\i50/n486 ),
    .C(\i50/n488 ),
    .D(\i50/n473 ),
    .E(\i50/n465 ),
    .Y(n20[6]));
 NAND3xp33_ASAP7_75t_SL \i50/i80  (.A(\i50/n314 ),
    .B(\i50/n342 ),
    .C(\i50/n520 ),
    .Y(\i50/n433 ));
 NAND2xp5_ASAP7_75t_L \i50/i81  (.A(\i50/n406 ),
    .B(\i50/n373 ),
    .Y(\i50/n432 ));
 NAND2xp5_ASAP7_75t_SL \i50/i82  (.A(\i50/n356 ),
    .B(\i50/n396 ),
    .Y(\i50/n431 ));
 NAND3xp33_ASAP7_75t_SL \i50/i83  (.A(\i50/n576 ),
    .B(\i50/n299 ),
    .C(\i50/n282 ),
    .Y(\i50/n444 ));
 NOR3xp33_ASAP7_75t_SL \i50/i84  (.A(\i50/n377 ),
    .B(\i50/n7 ),
    .C(\i50/n284 ),
    .Y(\i50/n430 ));
 NAND2xp5_ASAP7_75t_SL \i50/i85  (.A(\i50/n23 ),
    .B(\i50/n384 ),
    .Y(\i50/n443 ));
 OR3x1_ASAP7_75t_SL \i50/i86  (.A(\i50/n307 ),
    .B(\i50/n320 ),
    .C(\i50/n28 ),
    .Y(\i50/n429 ));
 NOR2x1_ASAP7_75t_SL \i50/i87  (.A(\i50/n318 ),
    .B(\i50/n409 ),
    .Y(\i50/n442 ));
 NOR2xp33_ASAP7_75t_L \i50/i88  (.A(\i50/n367 ),
    .B(\i50/n354 ),
    .Y(\i50/n441 ));
 NOR2xp67_ASAP7_75t_SL \i50/i89  (.A(\i50/n308 ),
    .B(\i50/n395 ),
    .Y(\i50/n440 ));
 AND3x4_ASAP7_75t_SL \i50/i9  (.A(\i50/n495 ),
    .B(\i50/n504 ),
    .C(\i50/n483 ),
    .Y(n20[1]));
 NOR3x1_ASAP7_75t_SL \i50/i90  (.A(\i50/n313 ),
    .B(\i50/n210 ),
    .C(\i50/n360 ),
    .Y(\i50/n439 ));
 NOR2xp67_ASAP7_75t_SL \i50/i91  (.A(\i50/n554 ),
    .B(\i50/n387 ),
    .Y(\i50/n438 ));
 NOR3xp33_ASAP7_75t_SL \i50/i92  (.A(\i50/n322 ),
    .B(\i50/n237 ),
    .C(\i50/n310 ),
    .Y(\i50/n425 ));
 NOR2xp33_ASAP7_75t_SL \i50/i93  (.A(\i50/n572 ),
    .B(\i50/n380 ),
    .Y(\i50/n424 ));
 NAND3xp33_ASAP7_75t_SL \i50/i94  (.A(\i50/n306 ),
    .B(\i50/n371 ),
    .C(\i50/n319 ),
    .Y(\i50/n423 ));
 NAND4xp25_ASAP7_75t_SL \i50/i95  (.A(\i50/n291 ),
    .B(\i50/n303 ),
    .C(\i50/n331 ),
    .D(\i50/n298 ),
    .Y(\i50/n422 ));
 NAND2x1_ASAP7_75t_SL \i50/i96  (.A(\i50/n394 ),
    .B(\i50/n408 ),
    .Y(\i50/n428 ));
 NOR5xp2_ASAP7_75t_SL \i50/i97  (.A(\i50/n403 ),
    .B(\i50/n516 ),
    .C(\i50/n136 ),
    .D(\i50/n252 ),
    .E(\i50/n178 ),
    .Y(\i50/n421 ));
 NAND3xp33_ASAP7_75t_SL \i50/i98  (.A(\i50/n359 ),
    .B(\i50/n378 ),
    .C(\i50/n524 ),
    .Y(\i50/n420 ));
 NAND2xp33_ASAP7_75t_SL \i50/i99  (.A(\i50/n300 ),
    .B(\i50/n400 ),
    .Y(\i50/n419 ));
 AOI22xp5_ASAP7_75t_SL i500 (.A1(n542),
    .A2(n510),
    .B1(n541),
    .B2(n511),
    .Y(n972));
 OAI22xp5_ASAP7_75t_SL i501 (.A1(n515),
    .A2(n124),
    .B1(n516),
    .B2(n474),
    .Y(n971));
 XNOR2xp5_ASAP7_75t_SL i502 (.A(n305),
    .B(n315),
    .Y(n970));
 AOI22xp5_ASAP7_75t_SL i503 (.A1(n517),
    .A2(n497),
    .B1(n518),
    .B2(n498),
    .Y(n969));
 XNOR2xp5_ASAP7_75t_SL i504 (.A(n296),
    .B(n345),
    .Y(n968));
 XOR2xp5_ASAP7_75t_SL i505 (.A(n297),
    .B(n299),
    .Y(n967));
 XOR2xp5_ASAP7_75t_SL i506 (.A(n768),
    .B(n298),
    .Y(n966));
 XOR2xp5_ASAP7_75t_SL i507 (.A(n300),
    .B(n301),
    .Y(n965));
 OAI22xp5_ASAP7_75t_SL i508 (.A1(n528),
    .A2(n498),
    .B1(n527),
    .B2(n497),
    .Y(n964));
 XOR2xp5_ASAP7_75t_SL i509 (.A(n307),
    .B(n306),
    .Y(n963));
 INVx2_ASAP7_75t_SL \i51/i0  (.A(n19[5]),
    .Y(\i51/n0 ));
 INVxp67_ASAP7_75t_SL \i51/i1  (.A(n19[4]),
    .Y(\i51/n1 ));
 NOR2x2_ASAP7_75t_SL \i51/i10  (.A(\i51/n438 ),
    .B(\i51/n444 ),
    .Y(n18[3]));
 NAND3xp33_ASAP7_75t_SL \i51/i100  (.A(\i51/n304 ),
    .B(\i51/n323 ),
    .C(\i51/n538 ),
    .Y(\i51/n362 ));
 NAND2xp33_ASAP7_75t_SL \i51/i101  (.A(\i51/n251 ),
    .B(\i51/n343 ),
    .Y(\i51/n361 ));
 NOR5xp2_ASAP7_75t_SL \i51/i102  (.A(\i51/n290 ),
    .B(\i51/n527 ),
    .C(\i51/n277 ),
    .D(\i51/n230 ),
    .E(\i51/n187 ),
    .Y(\i51/n360 ));
 NAND5xp2_ASAP7_75t_SL \i51/i103  (.A(\i51/n238 ),
    .B(\i51/n303 ),
    .C(\i51/n531 ),
    .D(\i51/n275 ),
    .E(\i51/n532 ),
    .Y(\i51/n359 ));
 NAND3xp33_ASAP7_75t_SL \i51/i104  (.A(\i51/n234 ),
    .B(\i51/n262 ),
    .C(\i51/n327 ),
    .Y(\i51/n358 ));
 NOR5xp2_ASAP7_75t_SL \i51/i105  (.A(\i51/n232 ),
    .B(\i51/n244 ),
    .C(\i51/n525 ),
    .D(\i51/n95 ),
    .E(\i51/n493 ),
    .Y(\i51/n357 ));
 NAND5xp2_ASAP7_75t_SL \i51/i106  (.A(\i51/n27 ),
    .B(\i51/n554 ),
    .C(\i51/n531 ),
    .D(\i51/n73 ),
    .E(\i51/n163 ),
    .Y(\i51/n356 ));
 NAND4xp25_ASAP7_75t_SL \i51/i107  (.A(\i51/n182 ),
    .B(\i51/n193 ),
    .C(\i51/n280 ),
    .D(\i51/n20 ),
    .Y(\i51/n355 ));
 NOR5xp2_ASAP7_75t_SL \i51/i108  (.A(\i51/n197 ),
    .B(\i51/n555 ),
    .C(\i51/n186 ),
    .D(\i51/n159 ),
    .E(\i51/n157 ),
    .Y(\i51/n354 ));
 NOR2xp33_ASAP7_75t_SL \i51/i109  (.A(\i51/n318 ),
    .B(\i51/n348 ),
    .Y(\i51/n353 ));
 AND5x2_ASAP7_75t_SL \i51/i11  (.A(\i51/n436 ),
    .B(\i51/n427 ),
    .C(\i51/n429 ),
    .D(\i51/n416 ),
    .E(\i51/n408 ),
    .Y(n18[6]));
 NOR2xp33_ASAP7_75t_SL \i51/i110  (.A(\i51/n565 ),
    .B(\i51/n335 ),
    .Y(\i51/n352 ));
 NAND3x1_ASAP7_75t_SL \i51/i111  (.A(\i51/n539 ),
    .B(\i51/n303 ),
    .C(\i51/n334 ),
    .Y(\i51/n369 ));
 NAND3x1_ASAP7_75t_SL \i51/i112  (.A(\i51/n299 ),
    .B(\i51/n281 ),
    .C(\i51/n252 ),
    .Y(\i51/n368 ));
 AOI21xp5_ASAP7_75t_L \i51/i113  (.A1(\i51/n467 ),
    .A2(\i51/n199 ),
    .B(\i51/n139 ),
    .Y(\i51/n345 ));
 NAND2xp5_ASAP7_75t_SL \i51/i114  (.A(\i51/n279 ),
    .B(\i51/n306 ),
    .Y(\i51/n344 ));
 NOR2xp33_ASAP7_75t_SL \i51/i115  (.A(\i51/n305 ),
    .B(\i51/n28 ),
    .Y(\i51/n343 ));
 NOR2xp33_ASAP7_75t_SL \i51/i116  (.A(\i51/n285 ),
    .B(\i51/n295 ),
    .Y(\i51/n342 ));
 NOR2xp67_ASAP7_75t_SL \i51/i117  (.A(\i51/n148 ),
    .B(\i51/n292 ),
    .Y(\i51/n341 ));
 NOR2xp33_ASAP7_75t_SL \i51/i118  (.A(\i51/n290 ),
    .B(\i51/n24 ),
    .Y(\i51/n340 ));
 NOR4xp25_ASAP7_75t_SL \i51/i119  (.A(\i51/n266 ),
    .B(\i51/n470 ),
    .C(\i51/n24 ),
    .D(\i51/n559 ),
    .Y(\i51/n339 ));
 AND3x4_ASAP7_75t_SL \i51/i12  (.A(\i51/n436 ),
    .B(\i51/n445 ),
    .C(\i51/n424 ),
    .Y(n18[1]));
 NAND2xp5_ASAP7_75t_SL \i51/i120  (.A(\i51/n223 ),
    .B(\i51/n272 ),
    .Y(\i51/n338 ));
 NOR4xp25_ASAP7_75t_SL \i51/i121  (.A(\i51/n92 ),
    .B(\i51/n214 ),
    .C(\i51/n189 ),
    .D(\i51/n200 ),
    .Y(\i51/n337 ));
 NOR3xp33_ASAP7_75t_SL \i51/i122  (.A(\i51/n220 ),
    .B(\i51/n491 ),
    .C(\i51/n219 ),
    .Y(\i51/n336 ));
 NAND2xp33_ASAP7_75t_SL \i51/i123  (.A(\i51/n480 ),
    .B(\i51/n25 ),
    .Y(\i51/n335 ));
 NOR2x1p5_ASAP7_75t_SL \i51/i124  (.A(\i51/n239 ),
    .B(\i51/n469 ),
    .Y(\i51/n334 ));
 NAND2xp33_ASAP7_75t_SL \i51/i125  (.A(\i51/n304 ),
    .B(\i51/n288 ),
    .Y(\i51/n333 ));
 NAND3xp33_ASAP7_75t_SL \i51/i126  (.A(\i51/n26 ),
    .B(\i51/n181 ),
    .C(\i51/n479 ),
    .Y(\i51/n332 ));
 NOR3xp33_ASAP7_75t_SL \i51/i127  (.A(\i51/n570 ),
    .B(\i51/n194 ),
    .C(\i51/n522 ),
    .Y(\i51/n351 ));
 NAND2xp5_ASAP7_75t_SL \i51/i128  (.A(\i51/n265 ),
    .B(\i51/n182 ),
    .Y(\i51/n350 ));
 NOR2x1_ASAP7_75t_SL \i51/i129  (.A(\i51/n237 ),
    .B(\i51/n260 ),
    .Y(\i51/n349 ));
 NOR2x1p5_ASAP7_75t_SL \i51/i13  (.A(\i51/n446 ),
    .B(\i51/n437 ),
    .Y(n18[5]));
 NAND2xp5_ASAP7_75t_SL \i51/i130  (.A(\i51/n531 ),
    .B(\i51/n267 ),
    .Y(\i51/n348 ));
 NOR2x1_ASAP7_75t_SL \i51/i131  (.A(\i51/n240 ),
    .B(\i51/n293 ),
    .Y(\i51/n347 ));
 NOR3x1_ASAP7_75t_SL \i51/i132  (.A(\i51/n186 ),
    .B(\i51/n179 ),
    .C(\i51/n156 ),
    .Y(\i51/n346 ));
 INVx1_ASAP7_75t_SL \i51/i133  (.A(\i51/n329 ),
    .Y(\i51/n330 ));
 INVx1_ASAP7_75t_SL \i51/i134  (.A(\i51/n29 ),
    .Y(\i51/n328 ));
 NOR4xp25_ASAP7_75t_SL \i51/i135  (.A(\i51/n458 ),
    .B(\i51/n568 ),
    .C(\i51/n192 ),
    .D(\i51/n168 ),
    .Y(\i51/n327 ));
 AOI211xp5_ASAP7_75t_SL \i51/i136  (.A1(\i51/n97 ),
    .A2(\i51/n46 ),
    .B(\i51/n276 ),
    .C(\i51/n218 ),
    .Y(\i51/n326 ));
 NAND2xp33_ASAP7_75t_L \i51/i137  (.A(\i51/n253 ),
    .B(\i51/n274 ),
    .Y(\i51/n325 ));
 NAND5xp2_ASAP7_75t_SL \i51/i138  (.A(\i51/n201 ),
    .B(\i51/n213 ),
    .C(\i51/n224 ),
    .D(\i51/n514 ),
    .E(\i51/n544 ),
    .Y(\i51/n324 ));
 NOR4xp25_ASAP7_75t_SL \i51/i139  (.A(\i51/n566 ),
    .B(\i51/n123 ),
    .C(\i51/n125 ),
    .D(\i51/n144 ),
    .Y(\i51/n323 ));
 AND2x4_ASAP7_75t_SL \i51/i14  (.A(\i51/n447 ),
    .B(\i51/n430 ),
    .Y(n18[0]));
 NOR2xp33_ASAP7_75t_SL \i51/i140  (.A(\i51/n245 ),
    .B(\i51/n248 ),
    .Y(\i51/n322 ));
 AOI211xp5_ASAP7_75t_SL \i51/i141  (.A1(\i51/n142 ),
    .A2(\i51/n57 ),
    .B(\i51/n457 ),
    .C(\i51/n161 ),
    .Y(\i51/n321 ));
 OA21x2_ASAP7_75t_SL \i51/i142  (.A1(\i51/n460 ),
    .A2(\i51/n467 ),
    .B(\i51/n554 ),
    .Y(\i51/n320 ));
 NOR4xp25_ASAP7_75t_SL \i51/i143  (.A(\i51/n226 ),
    .B(\i51/n152 ),
    .C(\i51/n176 ),
    .D(\i51/n156 ),
    .Y(\i51/n319 ));
 NAND5xp2_ASAP7_75t_SL \i51/i144  (.A(\i51/n124 ),
    .B(\i51/n81 ),
    .C(\i51/n134 ),
    .D(\i51/n126 ),
    .E(\i51/n75 ),
    .Y(\i51/n318 ));
 NOR3xp33_ASAP7_75t_SL \i51/i145  (.A(\i51/n261 ),
    .B(\i51/n154 ),
    .C(\i51/n72 ),
    .Y(\i51/n317 ));
 NAND2xp5_ASAP7_75t_SL \i51/i146  (.A(\i51/n243 ),
    .B(\i51/n27 ),
    .Y(\i51/n316 ));
 NAND5xp2_ASAP7_75t_SL \i51/i147  (.A(\i51/n180 ),
    .B(\i51/n86 ),
    .C(\i51/n173 ),
    .D(\i51/n167 ),
    .E(\i51/n166 ),
    .Y(\i51/n315 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i51/i148  (.A1(\i51/n60 ),
    .A2(\i51/n77 ),
    .B(\i51/n577 ),
    .C(\i51/n235 ),
    .Y(\i51/n314 ));
 NAND4xp25_ASAP7_75t_SL \i51/i149  (.A(\i51/n271 ),
    .B(\i51/n498 ),
    .C(\i51/n93 ),
    .D(\i51/n484 ),
    .Y(\i51/n313 ));
 NOR3xp33_ASAP7_75t_SL \i51/i15  (.A(\i51/n421 ),
    .B(\i51/n417 ),
    .C(\i51/n473 ),
    .Y(\i51/n447 ));
 NAND5xp2_ASAP7_75t_SL \i51/i150  (.A(\i51/n143 ),
    .B(\i51/n483 ),
    .C(\i51/n205 ),
    .D(\i51/n89 ),
    .E(\i51/n83 ),
    .Y(\i51/n312 ));
 NAND2xp5_ASAP7_75t_SL \i51/i151  (.A(\i51/n242 ),
    .B(\i51/n264 ),
    .Y(\i51/n311 ));
 NAND3xp33_ASAP7_75t_SL \i51/i152  (.A(\i51/n259 ),
    .B(\i51/n74 ),
    .C(\i51/n78 ),
    .Y(\i51/n310 ));
 NAND2xp5_ASAP7_75t_SL \i51/i153  (.A(\i51/n539 ),
    .B(\i51/n303 ),
    .Y(\i51/n309 ));
 NOR2xp33_ASAP7_75t_L \i51/i154  (.A(\i51/n283 ),
    .B(\i51/n295 ),
    .Y(\i51/n331 ));
 NAND2xp5_ASAP7_75t_SL \i51/i155  (.A(\i51/n538 ),
    .B(\i51/n304 ),
    .Y(\i51/n308 ));
 NOR2x1p5_ASAP7_75t_SL \i51/i156  (.A(\i51/n454 ),
    .B(\i51/n286 ),
    .Y(\i51/n329 ));
 NAND3x1_ASAP7_75t_SL \i51/i157  (.A(\i51/n229 ),
    .B(\i51/n541 ),
    .C(\i51/n128 ),
    .Y(\i51/n29 ));
 INVxp67_ASAP7_75t_SL \i51/i158  (.A(\i51/n565 ),
    .Y(\i51/n307 ));
 INVxp67_ASAP7_75t_SL \i51/i159  (.A(\i51/n9 ),
    .Y(\i51/n306 ));
 NOR2x2_ASAP7_75t_SL \i51/i16  (.A(\i51/n439 ),
    .B(\i51/n440 ),
    .Y(n18[2]));
 INVxp67_ASAP7_75t_SL \i51/i160  (.A(\i51/n301 ),
    .Y(\i51/n302 ));
 INVxp67_ASAP7_75t_SL \i51/i161  (.A(\i51/n567 ),
    .Y(\i51/n300 ));
 INVx2_ASAP7_75t_SL \i51/i162  (.A(\i51/n298 ),
    .Y(\i51/n299 ));
 INVxp67_ASAP7_75t_SL \i51/i163  (.A(\i51/n513 ),
    .Y(\i51/n297 ));
 INVxp67_ASAP7_75t_SL \i51/i164  (.A(\i51/n293 ),
    .Y(\i51/n294 ));
 INVxp67_ASAP7_75t_SL \i51/i165  (.A(\i51/n553 ),
    .Y(\i51/n291 ));
 INVx1_ASAP7_75t_SL \i51/i166  (.A(\i51/n288 ),
    .Y(\i51/n289 ));
 OAI31xp33_ASAP7_75t_SL \i51/i167  (.A1(\i51/n57 ),
    .A2(\i51/n5 ),
    .A3(\i51/n47 ),
    .B(\i51/n43 ),
    .Y(\i51/n287 ));
 NAND2x1_ASAP7_75t_SL \i51/i168  (.A(\i51/n191 ),
    .B(\i51/n190 ),
    .Y(\i51/n286 ));
 NAND2xp33_ASAP7_75t_SL \i51/i169  (.A(\i51/n181 ),
    .B(\i51/n531 ),
    .Y(\i51/n285 ));
 NAND4xp75_ASAP7_75t_SL \i51/i17  (.A(\i51/n407 ),
    .B(\i51/n425 ),
    .C(\i51/n405 ),
    .D(\i51/n578 ),
    .Y(\i51/n446 ));
 OAI21xp5_ASAP7_75t_SL \i51/i170  (.A1(\i51/n45 ),
    .A2(\i51/n117 ),
    .B(\i51/n165 ),
    .Y(\i51/n284 ));
 NAND2xp5_ASAP7_75t_SL \i51/i171  (.A(\i51/n155 ),
    .B(\i51/n181 ),
    .Y(\i51/n283 ));
 NOR3xp33_ASAP7_75t_SL \i51/i172  (.A(\i51/n491 ),
    .B(\i51/n116 ),
    .C(\i51/n102 ),
    .Y(\i51/n282 ));
 NOR3xp33_ASAP7_75t_SL \i51/i173  (.A(\i51/n543 ),
    .B(\i51/n110 ),
    .C(\i51/n225 ),
    .Y(\i51/n281 ));
 OAI31xp33_ASAP7_75t_SL \i51/i174  (.A1(\i51/n41 ),
    .A2(\i51/n43 ),
    .A3(\i51/n56 ),
    .B(\i51/n526 ),
    .Y(\i51/n280 ));
 AOI221xp5_ASAP7_75t_SL \i51/i175  (.A1(\i51/n60 ),
    .A2(\i51/n70 ),
    .B1(\i51/n552 ),
    .B2(\i51/n52 ),
    .C(\i51/n169 ),
    .Y(\i51/n279 ));
 OAI31xp33_ASAP7_75t_R \i51/i176  (.A1(\i51/n57 ),
    .A2(\i51/n59 ),
    .A3(\i51/n60 ),
    .B(\i51/n56 ),
    .Y(\i51/n278 ));
 OAI221xp5_ASAP7_75t_SL \i51/i177  (.A1(\i51/n19 ),
    .A2(\i51/n69 ),
    .B1(\i51/n42 ),
    .B2(\i51/n48 ),
    .C(\i51/n188 ),
    .Y(\i51/n277 ));
 AOI21xp33_ASAP7_75t_SL \i51/i178  (.A1(\i51/n149 ),
    .A2(\i51/n462 ),
    .B(\i51/n465 ),
    .Y(\i51/n276 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i51/i179  (.A1(\i51/n574 ),
    .A2(\i51/n7 ),
    .B(\i51/n68 ),
    .C(\i51/n21 ),
    .Y(\i51/n275 ));
 NOR3xp33_ASAP7_75t_SL \i51/i18  (.A(\i51/n472 ),
    .B(\i51/n391 ),
    .C(\i51/n433 ),
    .Y(\i51/n445 ));
 NOR3xp33_ASAP7_75t_SL \i51/i180  (.A(\i51/n198 ),
    .B(\i51/n543 ),
    .C(\i51/n122 ),
    .Y(\i51/n274 ));
 NAND3xp33_ASAP7_75t_SL \i51/i181  (.A(\i51/n22 ),
    .B(\i51/n516 ),
    .C(\i51/n147 ),
    .Y(\i51/n273 ));
 AOI22xp5_ASAP7_75t_SL \i51/i182  (.A1(\i51/n490 ),
    .A2(\i51/n571 ),
    .B1(\i51/n52 ),
    .B2(\i51/n47 ),
    .Y(\i51/n272 ));
 OAI21xp5_ASAP7_75t_SL \i51/i183  (.A1(\i51/n51 ),
    .A2(\i51/n140 ),
    .B(\i51/n57 ),
    .Y(\i51/n271 ));
 NAND4xp25_ASAP7_75t_SL \i51/i184  (.A(\i51/n158 ),
    .B(\i51/n484 ),
    .C(\i51/n504 ),
    .D(\i51/n129 ),
    .Y(\i51/n270 ));
 NAND2xp33_ASAP7_75t_SL \i51/i185  (.A(\i51/n208 ),
    .B(\i51/n121 ),
    .Y(\i51/n269 ));
 OAI211xp5_ASAP7_75t_SL \i51/i186  (.A1(\i51/n465 ),
    .A2(\i51/n54 ),
    .B(\i51/n131 ),
    .C(\i51/n135 ),
    .Y(\i51/n305 ));
 NOR2xp67_ASAP7_75t_SL \i51/i187  (.A(\i51/n548 ),
    .B(\i51/n525 ),
    .Y(\i51/n304 ));
 AOI21xp5_ASAP7_75t_SL \i51/i188  (.A1(\i51/n47 ),
    .A2(\i51/n51 ),
    .B(\i51/n457 ),
    .Y(\i51/n303 ));
 NAND2xp5_ASAP7_75t_SL \i51/i189  (.A(\i51/n210 ),
    .B(\i51/n535 ),
    .Y(\i51/n28 ));
 NAND4xp75_ASAP7_75t_SL \i51/i19  (.A(\i51/n406 ),
    .B(\i51/n435 ),
    .C(\i51/n411 ),
    .D(\i51/n401 ),
    .Y(\i51/n444 ));
 NOR2xp33_ASAP7_75t_SL \i51/i190  (.A(\i51/n211 ),
    .B(\i51/n226 ),
    .Y(\i51/n301 ));
 OR2x2_ASAP7_75t_SL \i51/i191  (.A(\i51/n563 ),
    .B(\i51/n557 ),
    .Y(\i51/n298 ));
 OAI211xp5_ASAP7_75t_SL \i51/i192  (.A1(\i51/n69 ),
    .A2(\i51/n62 ),
    .B(\i51/n162 ),
    .C(\i51/n112 ),
    .Y(\i51/n296 ));
 NAND2xp5_ASAP7_75t_SL \i51/i193  (.A(\i51/n532 ),
    .B(\i51/n481 ),
    .Y(\i51/n295 ));
 NAND2xp5_ASAP7_75t_SL \i51/i194  (.A(\i51/n26 ),
    .B(\i51/n170 ),
    .Y(\i51/n293 ));
 NAND2xp5_ASAP7_75t_SL \i51/i195  (.A(\i51/n537 ),
    .B(\i51/n207 ),
    .Y(\i51/n292 ));
 NAND2xp5_ASAP7_75t_SL \i51/i196  (.A(\i51/n160 ),
    .B(\i51/n177 ),
    .Y(\i51/n290 ));
 NOR2x1_ASAP7_75t_SL \i51/i197  (.A(\i51/n209 ),
    .B(\i51/n187 ),
    .Y(\i51/n288 ));
 INVxp67_ASAP7_75t_SL \i51/i198  (.A(\i51/n266 ),
    .Y(\i51/n267 ));
 INVx1_ASAP7_75t_SL \i51/i199  (.A(\i51/n262 ),
    .Y(\i51/n263 ));
 INVx2_ASAP7_75t_SL \i51/i2  (.A(n19[2]),
    .Y(\i51/n2 ));
 AND3x4_ASAP7_75t_SL \i51/i20  (.A(\i51/n426 ),
    .B(\i51/n441 ),
    .C(\i51/n431 ),
    .Y(n18[7]));
 INVx2_ASAP7_75t_SL \i51/i200  (.A(\i51/n259 ),
    .Y(\i51/n260 ));
 NAND4xp25_ASAP7_75t_SL \i51/i201  (.A(\i51/n94 ),
    .B(\i51/n113 ),
    .C(\i51/n99 ),
    .D(\i51/n98 ),
    .Y(\i51/n256 ));
 AOI31xp33_ASAP7_75t_SL \i51/i202  (.A1(\i51/n507 ),
    .A2(\i51/n467 ),
    .A3(\i51/n40 ),
    .B(\i51/n462 ),
    .Y(\i51/n255 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i51/i203  (.A1(\i51/n68 ),
    .A2(\i51/n44 ),
    .B(\i51/n56 ),
    .C(\i51/n118 ),
    .Y(\i51/n254 ));
 NOR4xp25_ASAP7_75t_SL \i51/i204  (.A(\i51/n92 ),
    .B(\i51/n459 ),
    .C(\i51/n164 ),
    .D(\i51/n71 ),
    .Y(\i51/n253 ));
 AOI211xp5_ASAP7_75t_SL \i51/i205  (.A1(\i51/n114 ),
    .A2(\i51/n576 ),
    .B(\i51/n154 ),
    .C(\i51/n79 ),
    .Y(\i51/n252 ));
 AOI21xp5_ASAP7_75t_SL \i51/i206  (.A1(\i51/n486 ),
    .A2(\i51/n68 ),
    .B(\i51/n202 ),
    .Y(\i51/n251 ));
 NOR2xp33_ASAP7_75t_L \i51/i207  (.A(\i51/n551 ),
    .B(\i51/n221 ),
    .Y(\i51/n250 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i51/i208  (.A1(\i51/n465 ),
    .A2(\i51/n461 ),
    .B(\i51/n66 ),
    .C(\i51/n497 ),
    .Y(\i51/n249 ));
 OAI22xp5_ASAP7_75t_SL \i51/i209  (.A1(\i51/n62 ),
    .A2(\i51/n141 ),
    .B1(\i51/n54 ),
    .B2(\i51/n508 ),
    .Y(\i51/n248 ));
 NAND4xp75_ASAP7_75t_SL \i51/i21  (.A(\i51/n390 ),
    .B(\i51/n410 ),
    .C(\i51/n419 ),
    .D(\i51/n434 ),
    .Y(\i51/n443 ));
 NOR2xp33_ASAP7_75t_SL \i51/i210  (.A(\i51/n184 ),
    .B(\i51/n171 ),
    .Y(\i51/n247 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i51/i211  (.A1(\i51/n490 ),
    .A2(\i51/n49 ),
    .B(\i51/n7 ),
    .C(\i51/n151 ),
    .Y(\i51/n246 ));
 NAND2xp33_ASAP7_75t_L \i51/i212  (.A(\i51/n91 ),
    .B(\i51/n178 ),
    .Y(\i51/n245 ));
 NAND2xp33_ASAP7_75t_SL \i51/i213  (.A(\i51/n217 ),
    .B(\i51/n111 ),
    .Y(\i51/n244 ));
 AOI22xp5_ASAP7_75t_SL \i51/i214  (.A1(\i51/n59 ),
    .A2(\i51/n88 ),
    .B1(\i51/n576 ),
    .B2(\i51/n60 ),
    .Y(\i51/n243 ));
 OAI21xp33_ASAP7_75t_SL \i51/i215  (.A1(\i51/n97 ),
    .A2(\i51/n59 ),
    .B(\i51/n576 ),
    .Y(\i51/n242 ));
 OA21x2_ASAP7_75t_SL \i51/i216  (.A1(\i51/n462 ),
    .A2(\i51/n117 ),
    .B(\i51/n106 ),
    .Y(\i51/n241 ));
 NAND2xp5_ASAP7_75t_SL \i51/i217  (.A(\i51/n482 ),
    .B(\i51/n231 ),
    .Y(\i51/n240 ));
 NAND4xp25_ASAP7_75t_SL \i51/i218  (.A(\i51/n108 ),
    .B(\i51/n130 ),
    .C(\i51/n85 ),
    .D(\i51/n506 ),
    .Y(\i51/n239 ));
 AOI221xp5_ASAP7_75t_SL \i51/i219  (.A1(\i51/n52 ),
    .A2(\i51/n39 ),
    .B1(\i51/n44 ),
    .B2(\i51/n53 ),
    .C(\i51/n558 ),
    .Y(\i51/n238 ));
 NAND2x1_ASAP7_75t_SL \i51/i22  (.A(\i51/n427 ),
    .B(\i51/n398 ),
    .Y(\i51/n442 ));
 OAI222xp33_ASAP7_75t_SL \i51/i220  (.A1(\i51/n10 ),
    .A2(\i51/n45 ),
    .B1(\i51/n48 ),
    .B2(\i51/n54 ),
    .C1(\i51/n499 ),
    .C2(\i51/n61 ),
    .Y(\i51/n237 ));
 AND3x1_ASAP7_75t_SL \i51/i221  (.A(\i51/n105 ),
    .B(\i51/n113 ),
    .C(\i51/n501 ),
    .Y(\i51/n236 ));
 AOI22xp5_ASAP7_75t_SL \i51/i222  (.A1(\i51/n452 ),
    .A2(\i51/n137 ),
    .B1(\i51/n51 ),
    .B2(\i51/n68 ),
    .Y(\i51/n268 ));
 NAND2xp33_ASAP7_75t_SL \i51/i223  (.A(\i51/n174 ),
    .B(\i51/n203 ),
    .Y(\i51/n235 ));
 NAND3x1_ASAP7_75t_SL \i51/i224  (.A(\i51/n502 ),
    .B(\i51/n133 ),
    .C(\i51/n127 ),
    .Y(\i51/n266 ));
 AOI22xp5_ASAP7_75t_SL \i51/i225  (.A1(\i51/n132 ),
    .A2(\i51/n526 ),
    .B1(\i51/n552 ),
    .B2(\i51/n56 ),
    .Y(\i51/n265 ));
 AOI22xp5_ASAP7_75t_SL \i51/i226  (.A1(\i51/n70 ),
    .A2(\i51/n492 ),
    .B1(\i51/n41 ),
    .B2(\i51/n57 ),
    .Y(\i51/n264 ));
 AOI221x1_ASAP7_75t_SL \i51/i227  (.A1(\i51/n526 ),
    .A2(\i51/n56 ),
    .B1(\i51/n60 ),
    .B2(\i51/n577 ),
    .C(\i51/n204 ),
    .Y(\i51/n262 ));
 OAI21xp5_ASAP7_75t_SL \i51/i228  (.A1(\i51/n40 ),
    .A2(\i51/n66 ),
    .B(\i51/n212 ),
    .Y(\i51/n261 ));
 NOR2x1_ASAP7_75t_SL \i51/i229  (.A(\i51/n107 ),
    .B(\i51/n172 ),
    .Y(\i51/n259 ));
 NOR2xp67_ASAP7_75t_SL \i51/i23  (.A(\i51/n392 ),
    .B(\i51/n428 ),
    .Y(\i51/n441 ));
 OAI211xp5_ASAP7_75t_SL \i51/i230  (.A1(\i51/n55 ),
    .A2(\i51/n84 ),
    .B(\i51/n93 ),
    .C(\i51/n534 ),
    .Y(\i51/n258 ));
 NOR2xp33_ASAP7_75t_L \i51/i231  (.A(\i51/n118 ),
    .B(\i51/n523 ),
    .Y(\i51/n27 ));
 NOR2xp33_ASAP7_75t_SL \i51/i232  (.A(\i51/n119 ),
    .B(\i51/n228 ),
    .Y(\i51/n234 ));
 AOI222xp33_ASAP7_75t_SL \i51/i233  (.A1(\i51/n60 ),
    .A2(\i51/n52 ),
    .B1(\i51/n7 ),
    .B2(\i51/n39 ),
    .C1(\i51/n57 ),
    .C2(\i51/n51 ),
    .Y(\i51/n257 ));
 INVx1_ASAP7_75t_SL \i51/i234  (.A(\i51/n537 ),
    .Y(\i51/n232 ));
 INVx1_ASAP7_75t_SL \i51/i235  (.A(\i51/n230 ),
    .Y(\i51/n231 ));
 INVx1_ASAP7_75t_SL \i51/i236  (.A(\i51/n228 ),
    .Y(\i51/n229 ));
 INVxp67_ASAP7_75t_SL \i51/i237  (.A(\i51/n481 ),
    .Y(\i51/n227 ));
 INVxp67_ASAP7_75t_SL \i51/i238  (.A(\i51/n524 ),
    .Y(\i51/n224 ));
 INVx1_ASAP7_75t_SL \i51/i239  (.A(\i51/n221 ),
    .Y(\i51/n222 ));
 NAND4xp75_ASAP7_75t_SL \i51/i24  (.A(\i51/n402 ),
    .B(\i51/n414 ),
    .C(\i51/n396 ),
    .D(\i51/n399 ),
    .Y(\i51/n440 ));
 OAI21xp33_ASAP7_75t_SL \i51/i240  (.A1(\i51/n58 ),
    .A2(\i51/n466 ),
    .B(\i51/n510 ),
    .Y(\i51/n219 ));
 NAND2xp5_ASAP7_75t_SL \i51/i241  (.A(\i51/n76 ),
    .B(\i51/n112 ),
    .Y(\i51/n218 ));
 OAI21xp5_ASAP7_75t_SL \i51/i242  (.A1(\i51/n552 ),
    .A2(\i51/n47 ),
    .B(\i51/n574 ),
    .Y(\i51/n217 ));
 NOR2xp33_ASAP7_75t_SL \i51/i243  (.A(\i51/n120 ),
    .B(\i51/n153 ),
    .Y(\i51/n216 ));
 AOI21xp5_ASAP7_75t_SL \i51/i244  (.A1(\i51/n478 ),
    .A2(\i51/n45 ),
    .B(\i51/n67 ),
    .Y(\i51/n215 ));
 NAND2xp33_ASAP7_75t_L \i51/i245  (.A(\i51/n150 ),
    .B(\i51/n80 ),
    .Y(\i51/n214 ));
 NOR2xp33_ASAP7_75t_SL \i51/i246  (.A(\i51/n21 ),
    .B(\i51/n100 ),
    .Y(\i51/n213 ));
 OAI21xp33_ASAP7_75t_SL \i51/i247  (.A1(\i51/n59 ),
    .A2(\i51/n65 ),
    .B(\i51/n52 ),
    .Y(\i51/n212 ));
 OAI21xp5_ASAP7_75t_SL \i51/i248  (.A1(\i51/n460 ),
    .A2(\i51/n67 ),
    .B(\i51/n485 ),
    .Y(\i51/n211 ));
 AOI22xp33_ASAP7_75t_SL \i51/i249  (.A1(\i51/n574 ),
    .A2(\i51/n49 ),
    .B1(\i51/n577 ),
    .B2(\i51/n57 ),
    .Y(\i51/n210 ));
 OR3x1_ASAP7_75t_SL \i51/i25  (.A(\i51/n422 ),
    .B(\i51/n420 ),
    .C(\i51/n403 ),
    .Y(\i51/n439 ));
 OAI21xp5_ASAP7_75t_SL \i51/i250  (.A1(\i51/n18 ),
    .A2(\i51/n499 ),
    .B(\i51/n115 ),
    .Y(\i51/n209 ));
 OAI21xp5_ASAP7_75t_SL \i51/i251  (.A1(\i51/n59 ),
    .A2(\i51/n47 ),
    .B(\i51/n53 ),
    .Y(\i51/n208 ));
 AOI22xp5_ASAP7_75t_SL \i51/i252  (.A1(\i51/n39 ),
    .A2(\i51/n70 ),
    .B1(\i51/n41 ),
    .B2(\i51/n59 ),
    .Y(\i51/n207 ));
 OA21x2_ASAP7_75t_SL \i51/i253  (.A1(\i51/n478 ),
    .A2(\i51/n16 ),
    .B(\i51/n514 ),
    .Y(\i51/n233 ));
 AOI21xp33_ASAP7_75t_SL \i51/i254  (.A1(\i51/n54 ),
    .A2(\i51/n478 ),
    .B(\i51/n40 ),
    .Y(\i51/n206 ));
 OAI21xp5_ASAP7_75t_SL \i51/i255  (.A1(\i51/n577 ),
    .A2(\i51/n70 ),
    .B(\i51/n452 ),
    .Y(\i51/n205 ));
 OA21x2_ASAP7_75t_SL \i51/i256  (.A1(\i51/n7 ),
    .A2(\i51/n70 ),
    .B(\i51/n68 ),
    .Y(\i51/n204 ));
 OAI21xp5_ASAP7_75t_SL \i51/i257  (.A1(\i51/n53 ),
    .A2(\i51/n41 ),
    .B(\i51/n452 ),
    .Y(\i51/n203 ));
 OAI21xp5_ASAP7_75t_SL \i51/i258  (.A1(\i51/n460 ),
    .A2(\i51/n499 ),
    .B(\i51/n25 ),
    .Y(\i51/n202 ));
 AOI22xp5_ASAP7_75t_SL \i51/i259  (.A1(\i51/n51 ),
    .A2(\i51/n490 ),
    .B1(\i51/n577 ),
    .B2(\i51/n49 ),
    .Y(\i51/n201 ));
 OR3x1_ASAP7_75t_SL \i51/i26  (.A(\i51/n423 ),
    .B(\i51/n389 ),
    .C(\i51/n362 ),
    .Y(\i51/n438 ));
 AOI21xp33_ASAP7_75t_SL \i51/i260  (.A1(\i51/n465 ),
    .A2(\i51/n40 ),
    .B(\i51/n55 ),
    .Y(\i51/n200 ));
 OAI21xp33_ASAP7_75t_SL \i51/i261  (.A1(\i51/n68 ),
    .A2(\i51/n59 ),
    .B(\i51/n43 ),
    .Y(\i51/n199 ));
 NAND2xp5_ASAP7_75t_SL \i51/i262  (.A(\i51/n452 ),
    .B(\i51/n486 ),
    .Y(\i51/n26 ));
 NAND2xp5_ASAP7_75t_L \i51/i263  (.A(\i51/n165 ),
    .B(\i51/n503 ),
    .Y(\i51/n198 ));
 OAI22xp5_ASAP7_75t_SL \i51/i264  (.A1(\i51/n536 ),
    .A2(\i51/n499 ),
    .B1(\i51/n19 ),
    .B2(\i51/n54 ),
    .Y(\i51/n230 ));
 OAI22xp5_ASAP7_75t_SL \i51/i265  (.A1(\i51/n69 ),
    .A2(\i51/n48 ),
    .B1(\i51/n62 ),
    .B2(\i51/n460 ),
    .Y(\i51/n228 ));
 OAI22xp5_ASAP7_75t_SL \i51/i266  (.A1(\i51/n55 ),
    .A2(\i51/n62 ),
    .B1(\i51/n499 ),
    .B2(\i51/n42 ),
    .Y(\i51/n226 ));
 NAND2xp5_ASAP7_75t_L \i51/i267  (.A(\i51/n20 ),
    .B(\i51/n136 ),
    .Y(\i51/n225 ));
 OAI21xp5_ASAP7_75t_SL \i51/i268  (.A1(\i51/n59 ),
    .A2(\i51/n44 ),
    .B(\i51/n574 ),
    .Y(\i51/n223 ));
 NOR2xp33_ASAP7_75t_L \i51/i269  (.A(\i51/n16 ),
    .B(\i51/n517 ),
    .Y(\i51/n221 ));
 NAND3xp33_ASAP7_75t_SL \i51/i27  (.A(\i51/n432 ),
    .B(\i51/n419 ),
    .C(\i51/n402 ),
    .Y(\i51/n437 ));
 NAND2xp33_ASAP7_75t_L \i51/i270  (.A(\i51/n93 ),
    .B(\i51/n534 ),
    .Y(\i51/n197 ));
 OAI21xp5_ASAP7_75t_SL \i51/i271  (.A1(\i51/n55 ),
    .A2(\i51/n48 ),
    .B(\i51/n544 ),
    .Y(\i51/n220 ));
 INVxp67_ASAP7_75t_SL \i51/i272  (.A(\i51/n195 ),
    .Y(\i51/n196 ));
 INVxp67_ASAP7_75t_SL \i51/i273  (.A(\i51/n193 ),
    .Y(\i51/n194 ));
 INVx1_ASAP7_75t_SL \i51/i274  (.A(\i51/n191 ),
    .Y(\i51/n192 ));
 INVx1_ASAP7_75t_SL \i51/i275  (.A(\i51/n521 ),
    .Y(\i51/n190 ));
 INVxp67_ASAP7_75t_SL \i51/i276  (.A(\i51/n188 ),
    .Y(\i51/n189 ));
 INVxp67_ASAP7_75t_SL \i51/i277  (.A(\i51/n184 ),
    .Y(\i51/n185 ));
 INVxp67_ASAP7_75t_SL \i51/i278  (.A(\i51/n570 ),
    .Y(\i51/n183 ));
 OAI21xp5_ASAP7_75t_SL \i51/i279  (.A1(\i51/n49 ),
    .A2(\i51/n63 ),
    .B(\i51/n577 ),
    .Y(\i51/n180 ));
 NOR2x1_ASAP7_75t_SL \i51/i28  (.A(\i51/n344 ),
    .B(\i51/n420 ),
    .Y(\i51/n435 ));
 OAI21xp5_ASAP7_75t_SL \i51/i280  (.A1(\i51/n17 ),
    .A2(\i51/n10 ),
    .B(\i51/n103 ),
    .Y(\i51/n179 ));
 OAI21xp33_ASAP7_75t_SL \i51/i281  (.A1(\i51/n552 ),
    .A2(\i51/n44 ),
    .B(\i51/n50 ),
    .Y(\i51/n178 ));
 AOI22xp5_ASAP7_75t_SL \i51/i282  (.A1(\i51/n576 ),
    .A2(\i51/n490 ),
    .B1(\i51/n43 ),
    .B2(\i51/n5 ),
    .Y(\i51/n177 ));
 AOI21xp33_ASAP7_75t_SL \i51/i283  (.A1(\i51/n499 ),
    .A2(\i51/n62 ),
    .B(\i51/n64 ),
    .Y(\i51/n176 ));
 AO21x1_ASAP7_75t_SL \i51/i284  (.A1(\i51/n39 ),
    .A2(\i51/n56 ),
    .B(\i51/n542 ),
    .Y(\i51/n175 ));
 OAI21xp5_ASAP7_75t_SL \i51/i285  (.A1(\i51/n39 ),
    .A2(\i51/n44 ),
    .B(\i51/n43 ),
    .Y(\i51/n174 ));
 OAI21xp5_ASAP7_75t_SL \i51/i286  (.A1(\i51/n576 ),
    .A2(\i51/n50 ),
    .B(\i51/n552 ),
    .Y(\i51/n173 ));
 OAI22xp33_ASAP7_75t_SL \i51/i287  (.A1(\i51/n19 ),
    .A2(\i51/n466 ),
    .B1(\i51/n62 ),
    .B2(\i51/n66 ),
    .Y(\i51/n172 ));
 OAI22xp33_ASAP7_75t_SL \i51/i288  (.A1(\i51/n461 ),
    .A2(\i51/n466 ),
    .B1(\i51/n16 ),
    .B2(\i51/n45 ),
    .Y(\i51/n171 ));
 AOI22xp5_ASAP7_75t_SL \i51/i289  (.A1(\i51/n52 ),
    .A2(\i51/n63 ),
    .B1(\i51/n41 ),
    .B2(\i51/n65 ),
    .Y(\i51/n170 ));
 NOR2x1_ASAP7_75t_SL \i51/i29  (.A(\i51/n404 ),
    .B(\i51/n400 ),
    .Y(\i51/n434 ));
 OAI21xp5_ASAP7_75t_SL \i51/i290  (.A1(\i51/n462 ),
    .A2(\i51/n48 ),
    .B(\i51/n101 ),
    .Y(\i51/n195 ));
 AOI22xp5_ASAP7_75t_SL \i51/i291  (.A1(\i51/n39 ),
    .A2(\i51/n53 ),
    .B1(\i51/n41 ),
    .B2(\i51/n47 ),
    .Y(\i51/n193 ));
 AOI22xp5_ASAP7_75t_SL \i51/i292  (.A1(\i51/n43 ),
    .A2(\i51/n44 ),
    .B1(\i51/n490 ),
    .B2(\i51/n52 ),
    .Y(\i51/n191 ));
 OAI22xp5_ASAP7_75t_SL \i51/i293  (.A1(\i51/n40 ),
    .A2(\i51/n17 ),
    .B1(\i51/n466 ),
    .B2(\i51/n467 ),
    .Y(\i51/n169 ));
 NAND2xp33_ASAP7_75t_SL \i51/i294  (.A(\i51/n166 ),
    .B(\i51/n167 ),
    .Y(\i51/n168 ));
 AOI22xp5_ASAP7_75t_SL \i51/i295  (.A1(\i51/n43 ),
    .A2(\i51/n490 ),
    .B1(\i51/n41 ),
    .B2(\i51/n68 ),
    .Y(\i51/n188 ));
 AO22x2_ASAP7_75t_SL \i51/i296  (.A1(\i51/n70 ),
    .A2(\i51/n526 ),
    .B1(\i51/n46 ),
    .B2(\i51/n65 ),
    .Y(\i51/n187 ));
 OAI21xp5_ASAP7_75t_SL \i51/i297  (.A1(\i51/n61 ),
    .A2(\i51/n461 ),
    .B(\i51/n87 ),
    .Y(\i51/n186 ));
 OAI22xp5_ASAP7_75t_L \i51/i298  (.A1(\i51/n64 ),
    .A2(\i51/n40 ),
    .B1(\i51/n62 ),
    .B2(\i51/n462 ),
    .Y(\i51/n184 ));
 AOI22xp5_ASAP7_75t_SL \i51/i299  (.A1(\i51/n39 ),
    .A2(\i51/n43 ),
    .B1(\i51/n56 ),
    .B2(\i51/n65 ),
    .Y(\i51/n182 ));
 INVx2_ASAP7_75t_SL \i51/i3  (.A(n19[0]),
    .Y(\i51/n3 ));
 NAND3xp33_ASAP7_75t_SL \i51/i30  (.A(\i51/n384 ),
    .B(\i51/n583 ),
    .C(\i51/n381 ),
    .Y(\i51/n433 ));
 AOI22xp5_ASAP7_75t_SL \i51/i300  (.A1(\i51/n50 ),
    .A2(\i51/n65 ),
    .B1(\i51/n41 ),
    .B2(\i51/n490 ),
    .Y(\i51/n181 ));
 INVxp67_ASAP7_75t_R \i51/i301  (.A(\i51/n505 ),
    .Y(\i51/n163 ));
 INVx1_ASAP7_75t_SL \i51/i302  (.A(\i51/n540 ),
    .Y(\i51/n162 ));
 INVxp67_ASAP7_75t_SL \i51/i303  (.A(\i51/n160 ),
    .Y(\i51/n161 ));
 INVxp67_ASAP7_75t_SL \i51/i304  (.A(\i51/n158 ),
    .Y(\i51/n159 ));
 INVxp67_ASAP7_75t_SL \i51/i305  (.A(\i51/n510 ),
    .Y(\i51/n157 ));
 INVxp67_ASAP7_75t_R \i51/i306  (.A(\i51/n559 ),
    .Y(\i51/n155 ));
 INVxp67_ASAP7_75t_SL \i51/i307  (.A(\i51/n485 ),
    .Y(\i51/n152 ));
 INVxp67_ASAP7_75t_SL \i51/i308  (.A(\i51/n150 ),
    .Y(\i51/n151 ));
 INVxp67_ASAP7_75t_SL \i51/i309  (.A(\i51/n147 ),
    .Y(\i51/n148 ));
 NOR2xp33_ASAP7_75t_SL \i51/i31  (.A(\i51/n409 ),
    .B(\i51/n371 ),
    .Y(\i51/n432 ));
 INVxp67_ASAP7_75t_SL \i51/i310  (.A(\i51/n145 ),
    .Y(\i51/n146 ));
 INVxp67_ASAP7_75t_SL \i51/i311  (.A(\i51/n143 ),
    .Y(\i51/n144 ));
 INVxp67_ASAP7_75t_SL \i51/i312  (.A(\i51/n141 ),
    .Y(\i51/n142 ));
 INVxp67_ASAP7_75t_SL \i51/i313  (.A(\i51/n517 ),
    .Y(\i51/n140 ));
 INVx1_ASAP7_75t_SL \i51/i314  (.A(\i51/n486 ),
    .Y(\i51/n139 ));
 NAND2xp5_ASAP7_75t_SL \i51/i315  (.A(\i51/n53 ),
    .B(\i51/n452 ),
    .Y(\i51/n167 ));
 NAND2xp5_ASAP7_75t_SL \i51/i316  (.A(\i51/n574 ),
    .B(\i51/n65 ),
    .Y(\i51/n138 ));
 NAND2xp5_ASAP7_75t_SL \i51/i317  (.A(\i51/n66 ),
    .B(\i51/n64 ),
    .Y(\i51/n137 ));
 NAND2xp5_ASAP7_75t_SL \i51/i318  (.A(\i51/n41 ),
    .B(\i51/n526 ),
    .Y(\i51/n136 ));
 NAND2xp5_ASAP7_75t_SL \i51/i319  (.A(\i51/n49 ),
    .B(\i51/n51 ),
    .Y(\i51/n135 ));
 NOR5xp2_ASAP7_75t_SL \i51/i32  (.A(\i51/n373 ),
    .B(\i51/n324 ),
    .C(\i51/n364 ),
    .D(\i51/n292 ),
    .E(\i51/n296 ),
    .Y(\i51/n431 ));
 NAND2xp5_ASAP7_75t_SL \i51/i320  (.A(\i51/n49 ),
    .B(\i51/n52 ),
    .Y(\i51/n166 ));
 NAND2xp5_ASAP7_75t_SL \i51/i321  (.A(\i51/n52 ),
    .B(\i51/n452 ),
    .Y(\i51/n134 ));
 NAND2xp5_ASAP7_75t_SL \i51/i322  (.A(\i51/n5 ),
    .B(\i51/n51 ),
    .Y(\i51/n133 ));
 NAND2xp5_ASAP7_75t_SL \i51/i323  (.A(\i51/n54 ),
    .B(\i51/n17 ),
    .Y(\i51/n132 ));
 NAND2xp5_ASAP7_75t_SL \i51/i324  (.A(\i51/n574 ),
    .B(\i51/n68 ),
    .Y(\i51/n131 ));
 NAND2xp5_ASAP7_75t_SL \i51/i325  (.A(\i51/n53 ),
    .B(\i51/n5 ),
    .Y(\i51/n130 ));
 NAND2xp5_ASAP7_75t_SL \i51/i326  (.A(\i51/n57 ),
    .B(\i51/n56 ),
    .Y(\i51/n129 ));
 NAND2xp5_ASAP7_75t_SL \i51/i327  (.A(\i51/n52 ),
    .B(\i51/n57 ),
    .Y(\i51/n128 ));
 NAND2x1_ASAP7_75t_SL \i51/i328  (.A(\i51/n46 ),
    .B(\i51/n39 ),
    .Y(\i51/n127 ));
 NAND2xp5_ASAP7_75t_SL \i51/i329  (.A(\i51/n53 ),
    .B(\i51/n68 ),
    .Y(\i51/n126 ));
 NOR3xp33_ASAP7_75t_SL \i51/i33  (.A(\i51/n369 ),
    .B(\i51/n386 ),
    .C(\i51/n418 ),
    .Y(\i51/n430 ));
 NAND2xp5_ASAP7_75t_SL \i51/i330  (.A(\i51/n39 ),
    .B(\i51/n577 ),
    .Y(\i51/n165 ));
 AND2x2_ASAP7_75t_SL \i51/i331  (.A(\i51/n46 ),
    .B(\i51/n59 ),
    .Y(\i51/n164 ));
 NAND2xp5_ASAP7_75t_SL \i51/i332  (.A(\i51/n57 ),
    .B(\i51/n7 ),
    .Y(\i51/n25 ));
 NAND2xp5_ASAP7_75t_SL \i51/i333  (.A(\i51/n577 ),
    .B(\i51/n68 ),
    .Y(\i51/n160 ));
 NAND2xp5_ASAP7_75t_SL \i51/i334  (.A(\i51/n70 ),
    .B(\i51/n44 ),
    .Y(\i51/n158 ));
 AND2x2_ASAP7_75t_SL \i51/i335  (.A(\i51/n53 ),
    .B(\i51/n490 ),
    .Y(\i51/n156 ));
 NOR2xp67_ASAP7_75t_SL \i51/i336  (.A(\i51/n478 ),
    .B(\i51/n499 ),
    .Y(\i51/n24 ));
 NOR2xp33_ASAP7_75t_SL \i51/i337  (.A(\i51/n55 ),
    .B(\i51/n62 ),
    .Y(\i51/n125 ));
 NAND2xp5_ASAP7_75t_SL \i51/i338  (.A(\i51/n490 ),
    .B(\i51/n51 ),
    .Y(\i51/n124 ));
 NOR2xp33_ASAP7_75t_SL \i51/i339  (.A(\i51/n466 ),
    .B(\i51/n62 ),
    .Y(\i51/n154 ));
 NOR2x1_ASAP7_75t_SL \i51/i34  (.A(\i51/n415 ),
    .B(\i51/n374 ),
    .Y(\i51/n429 ));
 AND2x2_ASAP7_75t_SL \i51/i340  (.A(\i51/n52 ),
    .B(\i51/n5 ),
    .Y(\i51/n153 ));
 NOR2xp33_ASAP7_75t_SL \i51/i341  (.A(\i51/n18 ),
    .B(\i51/n16 ),
    .Y(\i51/n123 ));
 NOR2xp33_ASAP7_75t_SL \i51/i342  (.A(\i51/n466 ),
    .B(\i51/n67 ),
    .Y(\i51/n122 ));
 NAND2xp5_ASAP7_75t_SL \i51/i343  (.A(\i51/n574 ),
    .B(\i51/n5 ),
    .Y(\i51/n150 ));
 NOR2xp33_ASAP7_75t_L \i51/i344  (.A(\i51/n70 ),
    .B(\i51/n43 ),
    .Y(\i51/n149 ));
 NAND2xp5_ASAP7_75t_SL \i51/i345  (.A(\i51/n70 ),
    .B(\i51/n47 ),
    .Y(\i51/n147 ));
 NAND2xp5_ASAP7_75t_SL \i51/i346  (.A(\i51/n68 ),
    .B(\i51/n52 ),
    .Y(\i51/n145 ));
 NAND2xp5_ASAP7_75t_SL \i51/i347  (.A(\i51/n70 ),
    .B(\i51/n57 ),
    .Y(\i51/n143 ));
 NAND2xp5_ASAP7_75t_SL \i51/i348  (.A(\i51/n53 ),
    .B(\i51/n60 ),
    .Y(\i51/n121 ));
 NOR2xp67_ASAP7_75t_SL \i51/i349  (.A(\i51/n574 ),
    .B(\i51/n53 ),
    .Y(\i51/n141 ));
 NAND2xp5_ASAP7_75t_SL \i51/i35  (.A(\i51/n372 ),
    .B(\i51/n393 ),
    .Y(\i51/n428 ));
 NOR2xp33_ASAP7_75t_SL \i51/i350  (.A(\i51/n48 ),
    .B(\i51/n66 ),
    .Y(\i51/n120 ));
 INVxp67_ASAP7_75t_SL \i51/i351  (.A(\i51/n541 ),
    .Y(\i51/n119 ));
 INVxp67_ASAP7_75t_SL \i51/i352  (.A(\i51/n115 ),
    .Y(\i51/n116 ));
 INVx1_ASAP7_75t_SL \i51/i353  (.A(\i51/n507 ),
    .Y(\i51/n114 ));
 INVxp67_ASAP7_75t_SL \i51/i354  (.A(\i51/n108 ),
    .Y(\i51/n109 ));
 INVxp67_ASAP7_75t_SL \i51/i355  (.A(\i51/n106 ),
    .Y(\i51/n107 ));
 INVxp67_ASAP7_75t_SL \i51/i356  (.A(\i51/n459 ),
    .Y(\i51/n105 ));
 INVxp67_ASAP7_75t_SL \i51/i357  (.A(\i51/n103 ),
    .Y(\i51/n104 ));
 INVxp67_ASAP7_75t_R \i51/i358  (.A(\i51/n533 ),
    .Y(\i51/n102 ));
 INVxp67_ASAP7_75t_SL \i51/i359  (.A(\i51/n100 ),
    .Y(\i51/n101 ));
 NOR3x1_ASAP7_75t_SL \i51/i36  (.A(\i51/n29 ),
    .B(\i51/n388 ),
    .C(\i51/n316 ),
    .Y(\i51/n436 ));
 INVxp67_ASAP7_75t_SL \i51/i360  (.A(\i51/n94 ),
    .Y(\i51/n95 ));
 INVx1_ASAP7_75t_SL \i51/i361  (.A(\i51/n91 ),
    .Y(\i51/n92 ));
 INVx2_ASAP7_75t_SL \i51/i362  (.A(\i51/n20 ),
    .Y(\i51/n21 ));
 NAND2xp5_ASAP7_75t_SL \i51/i363  (.A(\i51/n576 ),
    .B(\i51/n59 ),
    .Y(\i51/n90 ));
 NAND2xp5_ASAP7_75t_SL \i51/i364  (.A(\i51/n43 ),
    .B(\i51/n60 ),
    .Y(\i51/n89 ));
 NAND2xp5_ASAP7_75t_SL \i51/i365  (.A(\i51/n50 ),
    .B(\i51/n59 ),
    .Y(\i51/n23 ));
 NAND2xp5_ASAP7_75t_SL \i51/i366  (.A(\i51/n61 ),
    .B(\i51/n55 ),
    .Y(\i51/n88 ));
 NAND2xp5_ASAP7_75t_SL \i51/i367  (.A(\i51/n50 ),
    .B(\i51/n60 ),
    .Y(\i51/n87 ));
 NAND2xp5_ASAP7_75t_SL \i51/i368  (.A(\i51/n60 ),
    .B(\i51/n41 ),
    .Y(\i51/n86 ));
 NAND2xp5_ASAP7_75t_SL \i51/i369  (.A(\i51/n577 ),
    .B(\i51/n490 ),
    .Y(\i51/n85 ));
 NOR3xp33_ASAP7_75t_SL \i51/i37  (.A(\i51/n333 ),
    .B(\i51/n29 ),
    .C(\i51/n412 ),
    .Y(\i51/n426 ));
 NOR2xp33_ASAP7_75t_SL \i51/i370  (.A(\i51/n68 ),
    .B(\i51/n5 ),
    .Y(\i51/n84 ));
 NAND2xp5_ASAP7_75t_SL \i51/i371  (.A(\i51/n56 ),
    .B(\i51/n47 ),
    .Y(\i51/n83 ));
 NAND2xp5_ASAP7_75t_L \i51/i372  (.A(\i51/n19 ),
    .B(\i51/n40 ),
    .Y(\i51/n82 ));
 NAND2xp5_ASAP7_75t_SL \i51/i373  (.A(\i51/n7 ),
    .B(\i51/n49 ),
    .Y(\i51/n81 ));
 NAND2xp5_ASAP7_75t_SL \i51/i374  (.A(\i51/n576 ),
    .B(\i51/n49 ),
    .Y(\i51/n80 ));
 NOR2xp33_ASAP7_75t_SL \i51/i375  (.A(\i51/n48 ),
    .B(\i51/n460 ),
    .Y(\i51/n79 ));
 AND2x2_ASAP7_75t_SL \i51/i376  (.A(\i51/n7 ),
    .B(\i51/n60 ),
    .Y(\i51/n118 ));
 NOR2xp67_ASAP7_75t_L \i51/i377  (.A(\i51/n68 ),
    .B(\i51/n63 ),
    .Y(\i51/n117 ));
 NAND2xp5_ASAP7_75t_SL \i51/i378  (.A(\i51/n574 ),
    .B(\i51/n490 ),
    .Y(\i51/n115 ));
 NAND2xp5_ASAP7_75t_SL \i51/i379  (.A(\i51/n7 ),
    .B(\i51/n63 ),
    .Y(\i51/n113 ));
 NOR2xp33_ASAP7_75t_SL \i51/i38  (.A(\i51/n394 ),
    .B(\i51/n29 ),
    .Y(\i51/n425 ));
 NAND2xp5_ASAP7_75t_SL \i51/i380  (.A(\i51/n577 ),
    .B(\i51/n47 ),
    .Y(\i51/n112 ));
 NAND2xp5_ASAP7_75t_SL \i51/i381  (.A(\i51/n41 ),
    .B(\i51/n59 ),
    .Y(\i51/n78 ));
 NAND2xp5_ASAP7_75t_SL \i51/i382  (.A(\i51/n46 ),
    .B(\i51/n49 ),
    .Y(\i51/n111 ));
 AND2x2_ASAP7_75t_SL \i51/i383  (.A(\i51/n7 ),
    .B(\i51/n44 ),
    .Y(\i51/n110 ));
 NAND2xp5_ASAP7_75t_SL \i51/i384  (.A(\i51/n576 ),
    .B(\i51/n68 ),
    .Y(\i51/n108 ));
 NAND2xp5_ASAP7_75t_SL \i51/i385  (.A(\i51/n576 ),
    .B(\i51/n44 ),
    .Y(\i51/n106 ));
 NAND2xp5_ASAP7_75t_SL \i51/i386  (.A(\i51/n41 ),
    .B(\i51/n44 ),
    .Y(\i51/n103 ));
 NAND2xp33_ASAP7_75t_L \i51/i387  (.A(\i51/n461 ),
    .B(\i51/n58 ),
    .Y(\i51/n77 ));
 NOR2xp67_ASAP7_75t_L \i51/i388  (.A(\i51/n40 ),
    .B(\i51/n460 ),
    .Y(\i51/n100 ));
 NAND2xp5_ASAP7_75t_SL \i51/i389  (.A(\i51/n43 ),
    .B(\i51/n63 ),
    .Y(\i51/n22 ));
 NOR3xp33_ASAP7_75t_SL \i51/i39  (.A(\i51/n370 ),
    .B(\i51/n365 ),
    .C(\i51/n4 ),
    .Y(\i51/n424 ));
 NAND2xp5_ASAP7_75t_SL \i51/i390  (.A(\i51/n43 ),
    .B(\i51/n65 ),
    .Y(\i51/n99 ));
 NAND2xp5_ASAP7_75t_SL \i51/i391  (.A(\i51/n5 ),
    .B(\i51/n50 ),
    .Y(\i51/n98 ));
 NAND2xp5_ASAP7_75t_L \i51/i392  (.A(\i51/n16 ),
    .B(\i51/n19 ),
    .Y(\i51/n97 ));
 NAND2xp33_ASAP7_75t_L \i51/i393  (.A(\i51/n5 ),
    .B(\i51/n577 ),
    .Y(\i51/n76 ));
 NOR2xp33_ASAP7_75t_L \i51/i394  (.A(\i51/n552 ),
    .B(\i51/n59 ),
    .Y(\i51/n96 ));
 NAND2xp5_ASAP7_75t_SL \i51/i395  (.A(\i51/n7 ),
    .B(\i51/n65 ),
    .Y(\i51/n75 ));
 NAND2xp5_ASAP7_75t_SL \i51/i396  (.A(\i51/n50 ),
    .B(\i51/n47 ),
    .Y(\i51/n94 ));
 NAND2xp5_ASAP7_75t_SL \i51/i397  (.A(\i51/n41 ),
    .B(\i51/n5 ),
    .Y(\i51/n74 ));
 NAND2xp5_ASAP7_75t_SL \i51/i398  (.A(\i51/n577 ),
    .B(\i51/n65 ),
    .Y(\i51/n93 ));
 NAND2xp5_ASAP7_75t_SL \i51/i399  (.A(\i51/n50 ),
    .B(\i51/n63 ),
    .Y(\i51/n73 ));
 INVx1_ASAP7_75t_SL \i51/i4  (.A(\i51/n380 ),
    .Y(\i51/n4 ));
 NAND3xp33_ASAP7_75t_SL \i51/i40  (.A(\i51/n464 ),
    .B(\i51/n380 ),
    .C(\i51/n366 ),
    .Y(\i51/n423 ));
 NOR2xp33_ASAP7_75t_SL \i51/i400  (.A(\i51/n536 ),
    .B(\i51/n16 ),
    .Y(\i51/n72 ));
 NOR2xp33_ASAP7_75t_SL \i51/i401  (.A(\i51/n536 ),
    .B(\i51/n48 ),
    .Y(\i51/n71 ));
 NAND2xp5_ASAP7_75t_SL \i51/i402  (.A(\i51/n50 ),
    .B(\i51/n452 ),
    .Y(\i51/n91 ));
 NAND2x1p5_ASAP7_75t_L \i51/i403  (.A(\i51/n7 ),
    .B(\i51/n47 ),
    .Y(\i51/n20 ));
 INVx1_ASAP7_75t_SL \i51/i404  (.A(\i51/n70 ),
    .Y(\i51/n69 ));
 INVx3_ASAP7_75t_SL \i51/i405  (.A(\i51/n68 ),
    .Y(\i51/n67 ));
 INVx3_ASAP7_75t_SL \i51/i406  (.A(\i51/n574 ),
    .Y(\i51/n66 ));
 INVx2_ASAP7_75t_SL \i51/i407  (.A(\i51/n576 ),
    .Y(\i51/n64 ));
 INVx4_ASAP7_75t_SL \i51/i408  (.A(\i51/n63 ),
    .Y(\i51/n62 ));
 INVx2_ASAP7_75t_SL \i51/i409  (.A(\i51/n577 ),
    .Y(\i51/n61 ));
 NAND2xp5_ASAP7_75t_L \i51/i41  (.A(\i51/n579 ),
    .B(\i51/n413 ),
    .Y(\i51/n422 ));
 INVx2_ASAP7_75t_SL \i51/i410  (.A(\i51/n59 ),
    .Y(\i51/n58 ));
 INVx3_ASAP7_75t_SL \i51/i411  (.A(\i51/n56 ),
    .Y(\i51/n55 ));
 INVx3_ASAP7_75t_SL \i51/i412  (.A(\i51/n54 ),
    .Y(\i51/n53 ));
 AND2x4_ASAP7_75t_SL \i51/i413  (.A(\i51/n475 ),
    .B(\i51/n529 ),
    .Y(\i51/n70 ));
 AND2x4_ASAP7_75t_SL \i51/i414  (.A(\i51/n6 ),
    .B(\i51/n487 ),
    .Y(\i51/n68 ));
 AND2x4_ASAP7_75t_SL \i51/i415  (.A(\i51/n494 ),
    .B(\i51/n33 ),
    .Y(\i51/n65 ));
 NAND2x1_ASAP7_75t_SL \i51/i416  (.A(\i51/n494 ),
    .B(\i51/n33 ),
    .Y(\i51/n19 ));
 AND2x4_ASAP7_75t_SL \i51/i417  (.A(\i51/n488 ),
    .B(\i51/n495 ),
    .Y(\i51/n63 ));
 AND2x4_ASAP7_75t_SL \i51/i418  (.A(\i51/n494 ),
    .B(\i51/n32 ),
    .Y(\i51/n60 ));
 AND2x4_ASAP7_75t_SL \i51/i419  (.A(\i51/n487 ),
    .B(\i51/n15 ),
    .Y(\i51/n59 ));
 NAND2xp33_ASAP7_75t_SL \i51/i42  (.A(\i51/n377 ),
    .B(\i51/n395 ),
    .Y(\i51/n421 ));
 AND2x4_ASAP7_75t_SL \i51/i420  (.A(\i51/n487 ),
    .B(\i51/n494 ),
    .Y(\i51/n57 ));
 AND2x4_ASAP7_75t_SL \i51/i421  (.A(\i51/n475 ),
    .B(\i51/n509 ),
    .Y(\i51/n56 ));
 OR2x6_ASAP7_75t_SL \i51/i422  (.A(\i51/n36 ),
    .B(\i51/n573 ),
    .Y(\i51/n54 ));
 INVx3_ASAP7_75t_SL \i51/i423  (.A(\i51/n52 ),
    .Y(\i51/n18 ));
 INVx3_ASAP7_75t_SL \i51/i424  (.A(\i51/n49 ),
    .Y(\i51/n48 ));
 INVx3_ASAP7_75t_SL \i51/i425  (.A(\i51/n47 ),
    .Y(\i51/n16 ));
 INVx4_ASAP7_75t_SL \i51/i426  (.A(\i51/n46 ),
    .Y(\i51/n45 ));
 INVx3_ASAP7_75t_SL \i51/i427  (.A(\i51/n43 ),
    .Y(\i51/n42 ));
 INVx3_ASAP7_75t_SL \i51/i428  (.A(\i51/n40 ),
    .Y(\i51/n39 ));
 AND2x4_ASAP7_75t_SL \i51/i429  (.A(\i51/n529 ),
    .B(\i51/n38 ),
    .Y(\i51/n52 ));
 NOR2x1_ASAP7_75t_SL \i51/i43  (.A(\i51/n474 ),
    .B(\i51/n403 ),
    .Y(\i51/n427 ));
 OR2x2_ASAP7_75t_SL \i51/i430  (.A(\i51/n11 ),
    .B(\i51/n37 ),
    .Y(\i51/n17 ));
 AND2x4_ASAP7_75t_SL \i51/i431  (.A(\i51/n35 ),
    .B(\i51/n529 ),
    .Y(\i51/n51 ));
 NAND2x1p5_ASAP7_75t_SL \i51/i432  (.A(\i51/n6 ),
    .B(\i51/n32 ),
    .Y(\i51/n10 ));
 AND2x4_ASAP7_75t_SL \i51/i433  (.A(\i51/n35 ),
    .B(\i51/n476 ),
    .Y(\i51/n50 ));
 AND2x4_ASAP7_75t_SL \i51/i434  (.A(\i51/n32 ),
    .B(\i51/n15 ),
    .Y(\i51/n49 ));
 AND2x4_ASAP7_75t_SL \i51/i435  (.A(\i51/n495 ),
    .B(\i51/n15 ),
    .Y(\i51/n47 ));
 AND2x4_ASAP7_75t_SL \i51/i436  (.A(\i51/n8 ),
    .B(\i51/n476 ),
    .Y(\i51/n46 ));
 AND2x4_ASAP7_75t_SL \i51/i437  (.A(\i51/n6 ),
    .B(\i51/n33 ),
    .Y(\i51/n44 ));
 AND2x4_ASAP7_75t_SL \i51/i438  (.A(\i51/n509 ),
    .B(\i51/n35 ),
    .Y(\i51/n43 ));
 AND2x4_ASAP7_75t_SL \i51/i439  (.A(\i51/n38 ),
    .B(\i51/n509 ),
    .Y(\i51/n41 ));
 NAND2xp33_ASAP7_75t_L \i51/i44  (.A(\i51/n383 ),
    .B(\i51/n354 ),
    .Y(\i51/n418 ));
 OR2x6_ASAP7_75t_SL \i51/i440  (.A(\i51/n31 ),
    .B(\i51/n34 ),
    .Y(\i51/n40 ));
 INVx2_ASAP7_75t_SL \i51/i441  (.A(\i51/n37 ),
    .Y(\i51/n38 ));
 NAND2xp5_ASAP7_75t_SL \i51/i442  (.A(\i51/n12 ),
    .B(\i51/n2 ),
    .Y(\i51/n34 ));
 NAND2xp5_ASAP7_75t_SL \i51/i443  (.A(\i51/n1 ),
    .B(n19[5]),
    .Y(\i51/n37 ));
 NAND2x1p5_ASAP7_75t_SL \i51/i444  (.A(n19[4]),
    .B(n19[5]),
    .Y(\i51/n36 ));
 AND2x2_ASAP7_75t_SL \i51/i445  (.A(n19[4]),
    .B(\i51/n0 ),
    .Y(\i51/n35 ));
 INVx2_ASAP7_75t_SL \i51/i446  (.A(\i51/n519 ),
    .Y(\i51/n33 ));
 NAND2xp5_ASAP7_75t_SL \i51/i447  (.A(\i51/n30 ),
    .B(\i51/n3 ),
    .Y(\i51/n31 ));
 AND2x4_ASAP7_75t_SL \i51/i448  (.A(n19[0]),
    .B(\i51/n30 ),
    .Y(\i51/n32 ));
 INVx1_ASAP7_75t_SL \i51/i449  (.A(n19[1]),
    .Y(\i51/n30 ));
 NAND2xp33_ASAP7_75t_L \i51/i45  (.A(\i51/n579 ),
    .B(\i51/n360 ),
    .Y(\i51/n417 ));
 INVx2_ASAP7_75t_SL \i51/i450  (.A(\i51/n518 ),
    .Y(\i51/n15 ));
 INVx2_ASAP7_75t_SL \i51/i451  (.A(n19[6]),
    .Y(\i51/n14 ));
 INVx2_ASAP7_75t_SL \i51/i452  (.A(n19[7]),
    .Y(\i51/n13 ));
 INVx2_ASAP7_75t_SL \i51/i453  (.A(n19[3]),
    .Y(\i51/n12 ));
 NAND2xp33_ASAP7_75t_SL \i51/i454  (.A(\i51/n13 ),
    .B(n19[6]),
    .Y(\i51/n11 ));
 OR2x2_ASAP7_75t_SL \i51/i455  (.A(\i51/n110 ),
    .B(\i51/n557 ),
    .Y(\i51/n9 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i51/i456  (.A1(\i51/n69 ),
    .A2(\i51/n17 ),
    .B(\i51/n96 ),
    .C(\i51/n480 ),
    .Y(\i51/n448 ));
 INVx5_ASAP7_75t_SL \i51/i457  (.A(\i51/n451 ),
    .Y(\i51/n452 ));
 OR2x6_ASAP7_75t_SL \i51/i458  (.A(\i51/n449 ),
    .B(\i51/n450 ),
    .Y(\i51/n451 ));
 INVx1_ASAP7_75t_SL \i51/i459  (.A(\i51/n32 ),
    .Y(\i51/n449 ));
 NOR2xp33_ASAP7_75t_SL \i51/i46  (.A(\i51/n359 ),
    .B(\i51/n385 ),
    .Y(\i51/n416 ));
 INVx2_ASAP7_75t_SL \i51/i460  (.A(\i51/n488 ),
    .Y(\i51/n450 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i51/i461  (.A1(\i51/n451 ),
    .A2(\i51/n461 ),
    .B(\i51/n55 ),
    .C(\i51/n99 ),
    .Y(\i51/n453 ));
 OAI222xp33_ASAP7_75t_SL \i51/i462  (.A1(\i51/n451 ),
    .A2(\i51/n462 ),
    .B1(\i51/n461 ),
    .B2(\i51/n18 ),
    .C1(\i51/n467 ),
    .C2(\i51/n54 ),
    .Y(\i51/n454 ));
 OAI221xp5_ASAP7_75t_SL \i51/i463  (.A1(\i51/n451 ),
    .A2(\i51/n61 ),
    .B1(\i51/n499 ),
    .B2(\i51/n55 ),
    .C(\i51/n185 ),
    .Y(\i51/n455 ));
 OAI221xp5_ASAP7_75t_SL \i51/i464  (.A1(\i51/n451 ),
    .A2(\i51/n64 ),
    .B1(\i51/n19 ),
    .B2(\i51/n18 ),
    .C(\i51/n216 ),
    .Y(\i51/n456 ));
 OAI22xp5_ASAP7_75t_SL \i51/i465  (.A1(\i51/n466 ),
    .A2(\i51/n451 ),
    .B1(\i51/n536 ),
    .B2(\i51/n16 ),
    .Y(\i51/n457 ));
 OAI22xp5_ASAP7_75t_SL \i51/i466  (.A1(\i51/n69 ),
    .A2(\i51/n10 ),
    .B1(\i51/n17 ),
    .B2(\i51/n451 ),
    .Y(\i51/n458 ));
 NOR2xp67_ASAP7_75t_SL \i51/i467  (.A(\i51/n45 ),
    .B(\i51/n451 ),
    .Y(\i51/n459 ));
 INVx4_ASAP7_75t_SL \i51/i468  (.A(\i51/n50 ),
    .Y(\i51/n460 ));
 NAND2x1_ASAP7_75t_SL \i51/i469  (.A(\i51/n6 ),
    .B(\i51/n33 ),
    .Y(\i51/n461 ));
 NAND3xp33_ASAP7_75t_SL \i51/i47  (.A(\i51/n349 ),
    .B(\i51/n357 ),
    .C(\i51/n500 ),
    .Y(\i51/n415 ));
 INVx3_ASAP7_75t_SL \i51/i470  (.A(\i51/n41 ),
    .Y(\i51/n462 ));
 NOR2xp33_ASAP7_75t_SL \i51/i471  (.A(\i51/n290 ),
    .B(\i51/n549 ),
    .Y(\i51/n463 ));
 NOR2xp33_ASAP7_75t_SL \i51/i472  (.A(\i51/n550 ),
    .B(\i51/n258 ),
    .Y(\i51/n464 ));
 INVx3_ASAP7_75t_SL \i51/i473  (.A(\i51/n60 ),
    .Y(\i51/n465 ));
 INVx3_ASAP7_75t_SL \i51/i474  (.A(\i51/n51 ),
    .Y(\i51/n466 ));
 INVx3_ASAP7_75t_SL \i51/i475  (.A(\i51/n57 ),
    .Y(\i51/n467 ));
 AO21x2_ASAP7_75t_SL \i51/i476  (.A1(\i51/n576 ),
    .A2(\i51/n5 ),
    .B(\i51/n468 ),
    .Y(\i51/n469 ));
 OAI22xp5_ASAP7_75t_SL \i51/i477  (.A1(\i51/n465 ),
    .A2(\i51/n466 ),
    .B1(\i51/n467 ),
    .B2(\i51/n478 ),
    .Y(\i51/n468 ));
 OAI22x1_ASAP7_75t_SL \i51/i478  (.A1(\i51/n478 ),
    .A2(\i51/n62 ),
    .B1(\i51/n55 ),
    .B2(\i51/n451 ),
    .Y(\i51/n470 ));
 NAND4xp25_ASAP7_75t_SL \i51/i479  (.A(\i51/n352 ),
    .B(\i51/n471 ),
    .C(\i51/n346 ),
    .D(\i51/n379 ),
    .Y(\i51/n472 ));
 NOR2x1_ASAP7_75t_SL \i51/i48  (.A(\i51/n309 ),
    .B(\i51/n368 ),
    .Y(\i51/n414 ));
 NOR2x1_ASAP7_75t_SL \i51/i480  (.A(\i51/n470 ),
    .B(\i51/n549 ),
    .Y(\i51/n471 ));
 NAND3xp33_ASAP7_75t_L \i51/i481  (.A(\i51/n331 ),
    .B(\i51/n471 ),
    .C(\i51/n397 ),
    .Y(\i51/n473 ));
 NAND4xp25_ASAP7_75t_SL \i51/i482  (.A(\i51/n471 ),
    .B(\i51/n340 ),
    .C(\i51/n351 ),
    .D(\i51/n336 ),
    .Y(\i51/n474 ));
 AND2x4_ASAP7_75t_SL \i51/i483  (.A(\i51/n0 ),
    .B(\i51/n1 ),
    .Y(\i51/n475 ));
 AND2x2_ASAP7_75t_L \i51/i484  (.A(\i51/n13 ),
    .B(n19[6]),
    .Y(\i51/n476 ));
 INVx3_ASAP7_75t_SL \i51/i485  (.A(\i51/n477 ),
    .Y(\i51/n478 ));
 AND2x4_ASAP7_75t_SL \i51/i486  (.A(\i51/n475 ),
    .B(\i51/n476 ),
    .Y(\i51/n477 ));
 AOI22xp33_ASAP7_75t_SL \i51/i487  (.A1(\i51/n70 ),
    .A2(\i51/n552 ),
    .B1(\i51/n477 ),
    .B2(\i51/n5 ),
    .Y(\i51/n479 ));
 AOI211x1_ASAP7_75t_SL \i51/i488  (.A1(\i51/n82 ),
    .A2(\i51/n477 ),
    .B(\i51/n505 ),
    .C(\i51/n164 ),
    .Y(\i51/n480 ));
 AOI22xp5_ASAP7_75t_SL \i51/i489  (.A1(\i51/n477 ),
    .A2(\i51/n526 ),
    .B1(\i51/n7 ),
    .B2(\i51/n65 ),
    .Y(\i51/n481 ));
 NOR2xp33_ASAP7_75t_SL \i51/i49  (.A(\i51/n375 ),
    .B(\i51/n292 ),
    .Y(\i51/n413 ));
 AOI22xp33_ASAP7_75t_SL \i51/i490  (.A1(\i51/n477 ),
    .A2(\i51/n59 ),
    .B1(\i51/n7 ),
    .B2(\i51/n552 ),
    .Y(\i51/n482 ));
 NAND2xp5_ASAP7_75t_SL \i51/i491  (.A(\i51/n477 ),
    .B(\i51/n5 ),
    .Y(\i51/n483 ));
 NAND2xp5_ASAP7_75t_SL \i51/i492  (.A(\i51/n60 ),
    .B(\i51/n477 ),
    .Y(\i51/n484 ));
 NAND2xp5_ASAP7_75t_SL \i51/i493  (.A(\i51/n477 ),
    .B(\i51/n44 ),
    .Y(\i51/n485 ));
 OR2x2_ASAP7_75t_SL \i51/i494  (.A(\i51/n43 ),
    .B(\i51/n477 ),
    .Y(\i51/n486 ));
 AND2x2_ASAP7_75t_SL \i51/i495  (.A(n19[0]),
    .B(n19[1]),
    .Y(\i51/n487 ));
 AND2x2_ASAP7_75t_SL \i51/i496  (.A(\i51/n12 ),
    .B(\i51/n2 ),
    .Y(\i51/n488 ));
 INVx4_ASAP7_75t_SL \i51/i497  (.A(\i51/n489 ),
    .Y(\i51/n490 ));
 NAND2x1p5_ASAP7_75t_SL \i51/i498  (.A(\i51/n487 ),
    .B(\i51/n488 ),
    .Y(\i51/n489 ));
 OAI22xp5_ASAP7_75t_SL \i51/i499  (.A1(\i51/n45 ),
    .A2(\i51/n489 ),
    .B1(\i51/n54 ),
    .B2(\i51/n58 ),
    .Y(\i51/n491 ));
 INVx2_ASAP7_75t_SL \i51/i5  (.A(\i51/n10 ),
    .Y(\i51/n5 ));
 NAND2xp5_ASAP7_75t_SL \i51/i50  (.A(\i51/n383 ),
    .B(\i51/n378 ),
    .Y(\i51/n412 ));
 NAND2xp33_ASAP7_75t_SL \i51/i500  (.A(\i51/n489 ),
    .B(\i51/n10 ),
    .Y(\i51/n492 ));
 NOR2xp33_ASAP7_75t_SL \i51/i501  (.A(\i51/n489 ),
    .B(\i51/n462 ),
    .Y(\i51/n493 ));
 AND2x4_ASAP7_75t_SL \i51/i502  (.A(n19[2]),
    .B(n19[3]),
    .Y(\i51/n494 ));
 INVx2_ASAP7_75t_SL \i51/i503  (.A(\i51/n546 ),
    .Y(\i51/n495 ));
 OAI21xp5_ASAP7_75t_SL \i51/i504  (.A1(\i51/n496 ),
    .A2(\i51/n490 ),
    .B(\i51/n577 ),
    .Y(\i51/n497 ));
 AND2x4_ASAP7_75t_SL \i51/i505  (.A(\i51/n494 ),
    .B(\i51/n495 ),
    .Y(\i51/n496 ));
 OAI21xp5_ASAP7_75t_SL \i51/i506  (.A1(\i51/n496 ),
    .A2(\i51/n49 ),
    .B(\i51/n43 ),
    .Y(\i51/n498 ));
 INVx4_ASAP7_75t_SL \i51/i507  (.A(\i51/n496 ),
    .Y(\i51/n499 ));
 AOI211xp5_ASAP7_75t_SL \i51/i508  (.A1(\i51/n496 ),
    .A2(\i51/n53 ),
    .B(\i51/n469 ),
    .C(\i51/n153 ),
    .Y(\i51/n500 ));
 OAI21xp5_ASAP7_75t_SL \i51/i509  (.A1(\i51/n59 ),
    .A2(\i51/n496 ),
    .B(\i51/n70 ),
    .Y(\i51/n501 ));
 NOR2x1_ASAP7_75t_SL \i51/i51  (.A(\i51/n296 ),
    .B(\i51/n385 ),
    .Y(\i51/n411 ));
 OAI21xp5_ASAP7_75t_SL \i51/i510  (.A1(\i51/n50 ),
    .A2(\i51/n56 ),
    .B(\i51/n496 ),
    .Y(\i51/n502 ));
 NAND2xp5_ASAP7_75t_SL \i51/i511  (.A(\i51/n51 ),
    .B(\i51/n496 ),
    .Y(\i51/n503 ));
 NAND2xp5_ASAP7_75t_SL \i51/i512  (.A(\i51/n46 ),
    .B(\i51/n496 ),
    .Y(\i51/n504 ));
 AND2x2_ASAP7_75t_SL \i51/i513  (.A(\i51/n574 ),
    .B(\i51/n496 ),
    .Y(\i51/n505 ));
 NAND2xp5_ASAP7_75t_SL \i51/i514  (.A(\i51/n41 ),
    .B(\i51/n496 ),
    .Y(\i51/n506 ));
 NOR2x1_ASAP7_75t_SL \i51/i515  (.A(\i51/n496 ),
    .B(\i51/n65 ),
    .Y(\i51/n507 ));
 NOR2xp33_ASAP7_75t_SL \i51/i516  (.A(\i51/n496 ),
    .B(\i51/n49 ),
    .Y(\i51/n508 ));
 AND2x2_ASAP7_75t_SL \i51/i517  (.A(n19[7]),
    .B(\i51/n14 ),
    .Y(\i51/n509 ));
 NAND2xp5_ASAP7_75t_SL \i51/i518  (.A(\i51/n512 ),
    .B(\i51/n496 ),
    .Y(\i51/n510 ));
 OAI31xp33_ASAP7_75t_SL \i51/i519  (.A1(\i51/n490 ),
    .A2(\i51/n552 ),
    .A3(\i51/n526 ),
    .B(\i51/n512 ),
    .Y(\i51/n511 ));
 NOR2x1_ASAP7_75t_SL \i51/i52  (.A(\i51/n358 ),
    .B(\i51/n369 ),
    .Y(\i51/n410 ));
 AOI21xp5_ASAP7_75t_SL \i51/i520  (.A1(\i51/n59 ),
    .A2(\i51/n512 ),
    .B(\i51/n524 ),
    .Y(\i51/n513 ));
 NAND2xp5_ASAP7_75t_SL \i51/i521  (.A(\i51/n512 ),
    .B(\i51/n49 ),
    .Y(\i51/n514 ));
 NOR2xp33_ASAP7_75t_SL \i51/i522  (.A(\i51/n512 ),
    .B(\i51/n574 ),
    .Y(\i51/n515 ));
 NAND2xp5_ASAP7_75t_SL \i51/i523  (.A(\i51/n512 ),
    .B(\i51/n63 ),
    .Y(\i51/n516 ));
 NOR2x1_ASAP7_75t_SL \i51/i524  (.A(\i51/n512 ),
    .B(\i51/n576 ),
    .Y(\i51/n517 ));
 NAND2x1_ASAP7_75t_SL \i51/i525  (.A(n19[3]),
    .B(\i51/n2 ),
    .Y(\i51/n518 ));
 OR2x2_ASAP7_75t_SL \i51/i526  (.A(n19[0]),
    .B(n19[1]),
    .Y(\i51/n519 ));
 OAI22x1_ASAP7_75t_SL \i51/i527  (.A1(\i51/n18 ),
    .A2(\i51/n520 ),
    .B1(\i51/n58 ),
    .B2(\i51/n42 ),
    .Y(\i51/n521 ));
 OR2x2_ASAP7_75t_SL \i51/i528  (.A(\i51/n518 ),
    .B(\i51/n519 ),
    .Y(\i51/n520 ));
 OAI22xp5_ASAP7_75t_SL \i51/i529  (.A1(\i51/n466 ),
    .A2(\i51/n520 ),
    .B1(\i51/n54 ),
    .B2(\i51/n16 ),
    .Y(\i51/n522 ));
 NAND2xp5_ASAP7_75t_SL \i51/i53  (.A(\i51/n326 ),
    .B(\i51/n363 ),
    .Y(\i51/n409 ));
 OAI22xp5_ASAP7_75t_SL \i51/i530  (.A1(\i51/n520 ),
    .A2(\i51/n45 ),
    .B1(\i51/n42 ),
    .B2(\i51/n16 ),
    .Y(\i51/n523 ));
 OAI22xp5_ASAP7_75t_SL \i51/i531  (.A1(\i51/n460 ),
    .A2(\i51/n520 ),
    .B1(\i51/n54 ),
    .B2(\i51/n67 ),
    .Y(\i51/n524 ));
 OAI22xp5_ASAP7_75t_SL \i51/i532  (.A1(\i51/n536 ),
    .A2(\i51/n520 ),
    .B1(\i51/n462 ),
    .B2(\i51/n10 ),
    .Y(\i51/n525 ));
 INVx3_ASAP7_75t_SL \i51/i533  (.A(\i51/n520 ),
    .Y(\i51/n526 ));
 OAI221xp5_ASAP7_75t_SL \i51/i534  (.A1(\i51/n517 ),
    .A2(\i51/n520 ),
    .B1(\i51/n489 ),
    .B2(\i51/n55 ),
    .C(\i51/n145 ),
    .Y(\i51/n527 ));
 OAI221xp5_ASAP7_75t_SL \i51/i535  (.A1(\i51/n520 ),
    .A2(\i51/n66 ),
    .B1(\i51/n499 ),
    .B2(\i51/n17 ),
    .C(\i51/n90 ),
    .Y(\i51/n528 ));
 AND2x2_ASAP7_75t_SL \i51/i536  (.A(\i51/n13 ),
    .B(\i51/n14 ),
    .Y(\i51/n529 ));
 AOI22xp5_ASAP7_75t_SL \i51/i537  (.A1(\i51/n530 ),
    .A2(\i51/n44 ),
    .B1(\i51/n512 ),
    .B2(\i51/n57 ),
    .Y(\i51/n531 ));
 AND2x4_ASAP7_75t_SL \i51/i538  (.A(\i51/n529 ),
    .B(\i51/n8 ),
    .Y(\i51/n530 ));
 AOI22xp33_ASAP7_75t_SL \i51/i539  (.A1(\i51/n477 ),
    .A2(\i51/n490 ),
    .B1(\i51/n530 ),
    .B2(\i51/n49 ),
    .Y(\i51/n532 ));
 NOR5xp2_ASAP7_75t_SL \i51/i54  (.A(\i51/n258 ),
    .B(\i51/n553 ),
    .C(\i51/n528 ),
    .D(\i51/n28 ),
    .E(\i51/n455 ),
    .Y(\i51/n408 ));
 NAND2xp5_ASAP7_75t_SL \i51/i540  (.A(\i51/n39 ),
    .B(\i51/n530 ),
    .Y(\i51/n533 ));
 NAND2xp5_ASAP7_75t_SL \i51/i541  (.A(\i51/n530 ),
    .B(\i51/n5 ),
    .Y(\i51/n534 ));
 AOI22xp5_ASAP7_75t_SL \i51/i542  (.A1(\i51/n68 ),
    .A2(\i51/n530 ),
    .B1(\i51/n576 ),
    .B2(\i51/n57 ),
    .Y(\i51/n535 ));
 INVx2_ASAP7_75t_SL \i51/i543  (.A(\i51/n530 ),
    .Y(\i51/n536 ));
 AOI22xp5_ASAP7_75t_SL \i51/i544  (.A1(\i51/n530 ),
    .A2(\i51/n63 ),
    .B1(\i51/n577 ),
    .B2(\i51/n5 ),
    .Y(\i51/n537 ));
 AOI22xp5_ASAP7_75t_SL \i51/i545  (.A1(\i51/n530 ),
    .A2(\i51/n452 ),
    .B1(\i51/n574 ),
    .B2(\i51/n47 ),
    .Y(\i51/n538 ));
 AOI22xp33_ASAP7_75t_SL \i51/i546  (.A1(\i51/n39 ),
    .A2(\i51/n41 ),
    .B1(\i51/n530 ),
    .B2(\i51/n59 ),
    .Y(\i51/n539 ));
 AND2x2_ASAP7_75t_SL \i51/i547  (.A(\i51/n530 ),
    .B(\i51/n57 ),
    .Y(\i51/n540 ));
 NAND2xp5_ASAP7_75t_SL \i51/i548  (.A(\i51/n530 ),
    .B(\i51/n552 ),
    .Y(\i51/n541 ));
 AND2x2_ASAP7_75t_SL \i51/i549  (.A(\i51/n530 ),
    .B(\i51/n65 ),
    .Y(\i51/n542 ));
 NOR2x1_ASAP7_75t_SL \i51/i55  (.A(\i51/n4 ),
    .B(\i51/n370 ),
    .Y(\i51/n407 ));
 AND2x2_ASAP7_75t_SL \i51/i550  (.A(\i51/n530 ),
    .B(\i51/n490 ),
    .Y(\i51/n543 ));
 NAND2xp5_ASAP7_75t_SL \i51/i551  (.A(\i51/n530 ),
    .B(\i51/n60 ),
    .Y(\i51/n544 ));
 OR2x2_ASAP7_75t_SL \i51/i552  (.A(\i51/n2 ),
    .B(n19[3]),
    .Y(\i51/n545 ));
 NAND2xp5_ASAP7_75t_SL \i51/i553  (.A(\i51/n3 ),
    .B(n19[1]),
    .Y(\i51/n546 ));
 OAI22xp33_ASAP7_75t_SL \i51/i554  (.A1(\i51/n42 ),
    .A2(\i51/n520 ),
    .B1(\i51/n547 ),
    .B2(\i51/n466 ),
    .Y(\i51/n548 ));
 OR2x4_ASAP7_75t_SL \i51/i555  (.A(\i51/n545 ),
    .B(\i51/n546 ),
    .Y(\i51/n547 ));
 OAI221xp5_ASAP7_75t_SL \i51/i556  (.A1(\i51/n460 ),
    .A2(\i51/n461 ),
    .B1(\i51/n547 ),
    .B2(\i51/n462 ),
    .C(\i51/n533 ),
    .Y(\i51/n549 ));
 OAI221xp5_ASAP7_75t_L \i51/i557  (.A1(\i51/n460 ),
    .A2(\i51/n461 ),
    .B1(\i51/n547 ),
    .B2(\i51/n462 ),
    .C(\i51/n533 ),
    .Y(\i51/n550 ));
 OAI21xp5_ASAP7_75t_SL \i51/i558  (.A1(\i51/n61 ),
    .A2(\i51/n547 ),
    .B(\i51/n111 ),
    .Y(\i51/n551 ));
 INVx4_ASAP7_75t_SL \i51/i559  (.A(\i51/n547 ),
    .Y(\i51/n552 ));
 NAND2xp5_ASAP7_75t_SL \i51/i56  (.A(\i51/n367 ),
    .B(\i51/n347 ),
    .Y(\i51/n420 ));
 OAI221xp5_ASAP7_75t_SL \i51/i560  (.A1(\i51/n48 ),
    .A2(\i51/n478 ),
    .B1(\i51/n45 ),
    .B2(\i51/n547 ),
    .C(\i51/n23 ),
    .Y(\i51/n553 ));
 AO21x1_ASAP7_75t_SL \i51/i561  (.A1(\i51/n547 ),
    .A2(\i51/n138 ),
    .B(\i51/n515 ),
    .Y(\i51/n554 ));
 AOI31xp33_ASAP7_75t_SL \i51/i562  (.A1(\i51/n45 ),
    .A2(\i51/n64 ),
    .A3(\i51/n55 ),
    .B(\i51/n547 ),
    .Y(\i51/n555 ));
 OA21x2_ASAP7_75t_SL \i51/i563  (.A1(\i51/n45 ),
    .A2(\i51/n547 ),
    .B(\i51/n23 ),
    .Y(\i51/n556 ));
 OAI22xp5_ASAP7_75t_SL \i51/i564  (.A1(\i51/n45 ),
    .A2(\i51/n62 ),
    .B1(\i51/n54 ),
    .B2(\i51/n547 ),
    .Y(\i51/n557 ));
 OAI22xp5_ASAP7_75t_SL \i51/i565  (.A1(\i51/n45 ),
    .A2(\i51/n461 ),
    .B1(\i51/n547 ),
    .B2(\i51/n42 ),
    .Y(\i51/n558 ));
 NOR2xp33_ASAP7_75t_SL \i51/i566  (.A(\i51/n547 ),
    .B(\i51/n478 ),
    .Y(\i51/n559 ));
 NOR2xp33_ASAP7_75t_SL \i51/i567  (.A(\i51/n547 ),
    .B(\i51/n42 ),
    .Y(\i51/n560 ));
 AND2x4_ASAP7_75t_SL \i51/i568  (.A(\i51/n8 ),
    .B(\i51/n509 ),
    .Y(\i51/n512 ));
 OAI222xp33_ASAP7_75t_SL \i51/i569  (.A1(\i51/n62 ),
    .A2(\i51/n64 ),
    .B1(\i51/n520 ),
    .B2(\i51/n61 ),
    .C1(\i51/n19 ),
    .C2(\i51/n561 ),
    .Y(\i51/n562 ));
 NOR2x1_ASAP7_75t_SL \i51/i57  (.A(\i51/n386 ),
    .B(\i51/n369 ),
    .Y(\i51/n406 ));
 INVx4_ASAP7_75t_SL \i51/i570  (.A(\i51/n512 ),
    .Y(\i51/n561 ));
 OAI22xp33_ASAP7_75t_SL \i51/i571  (.A1(\i51/n466 ),
    .A2(\i51/n40 ),
    .B1(\i51/n451 ),
    .B2(\i51/n561 ),
    .Y(\i51/n563 ));
 AOI21xp5_ASAP7_75t_L \i51/i572  (.A1(\i51/n561 ),
    .A2(\i51/n149 ),
    .B(\i51/n451 ),
    .Y(\i51/n564 ));
 AOI21xp5_ASAP7_75t_SL \i51/i573  (.A1(\i51/n139 ),
    .A2(\i51/n561 ),
    .B(\i51/n67 ),
    .Y(\i51/n565 ));
 AOI31xp33_ASAP7_75t_SL \i51/i574  (.A1(\i51/n45 ),
    .A2(\i51/n18 ),
    .A3(\i51/n561 ),
    .B(\i51/n40 ),
    .Y(\i51/n566 ));
 OAI211xp5_ASAP7_75t_SL \i51/i575  (.A1(\i51/n561 ),
    .A2(\i51/n465 ),
    .B(\i51/n165 ),
    .C(\i51/n503 ),
    .Y(\i51/n567 ));
 AOI21xp33_ASAP7_75t_SL \i51/i576  (.A1(\i51/n561 ),
    .A2(\i51/n66 ),
    .B(\i51/n40 ),
    .Y(\i51/n568 ));
 OAI22xp5_ASAP7_75t_SL \i51/i577  (.A1(\i51/n561 ),
    .A2(\i51/n10 ),
    .B1(\i51/n66 ),
    .B2(\i51/n465 ),
    .Y(\i51/n569 ));
 OAI22xp5_ASAP7_75t_SL \i51/i578  (.A1(\i51/n561 ),
    .A2(\i51/n461 ),
    .B1(\i51/n54 ),
    .B2(\i51/n62 ),
    .Y(\i51/n570 ));
 NAND2xp33_ASAP7_75t_SL \i51/i579  (.A(\i51/n561 ),
    .B(\i51/n460 ),
    .Y(\i51/n571 ));
 NOR2x1_ASAP7_75t_SL \i51/i58  (.A(\i51/n308 ),
    .B(\i51/n368 ),
    .Y(\i51/n419 ));
 INVx2_ASAP7_75t_SL \i51/i580  (.A(\i51/n572 ),
    .Y(\i51/n573 ));
 AND2x2_ASAP7_75t_SL \i51/i581  (.A(n19[7]),
    .B(n19[6]),
    .Y(\i51/n572 ));
 AND2x4_ASAP7_75t_SL \i51/i582  (.A(\i51/n572 ),
    .B(\i51/n38 ),
    .Y(\i51/n574 ));
 AOI211xp5_ASAP7_75t_SL \i51/i583  (.A1(\i51/n526 ),
    .A2(\i51/n572 ),
    .B(\i51/n542 ),
    .C(\i51/n104 ),
    .Y(\i51/n575 ));
 AND2x4_ASAP7_75t_SL \i51/i584  (.A(\i51/n572 ),
    .B(\i51/n475 ),
    .Y(\i51/n576 ));
 AND2x4_ASAP7_75t_SL \i51/i585  (.A(\i51/n572 ),
    .B(\i51/n35 ),
    .Y(\i51/n577 ));
 AND4x1_ASAP7_75t_SL \i51/i586  (.A(\i51/n257 ),
    .B(\i51/n294 ),
    .C(\i51/n581 ),
    .D(\i51/n233 ),
    .Y(\i51/n578 ));
 AND4x1_ASAP7_75t_SL \i51/i587  (.A(\i51/n247 ),
    .B(\i51/n513 ),
    .C(\i51/n268 ),
    .D(\i51/n257 ),
    .Y(\i51/n579 ));
 OR4x1_ASAP7_75t_SL \i51/i588  (.A(\i51/n215 ),
    .B(\i51/n227 ),
    .C(\i51/n225 ),
    .D(\i51/n220 ),
    .Y(\i51/n580 ));
 AOI21xp5_ASAP7_75t_SL \i51/i589  (.A1(\i51/n46 ),
    .A2(\i51/n57 ),
    .B(\i51/n558 ),
    .Y(\i51/n581 ));
 INVxp67_ASAP7_75t_SL \i51/i59  (.A(\i51/n404 ),
    .Y(\i51/n405 ));
 NOR3xp33_ASAP7_75t_SL \i51/i590  (.A(\i51/n582 ),
    .B(\i51/n284 ),
    .C(\i51/n468 ),
    .Y(\i51/n583 ));
 OAI21xp5_ASAP7_75t_SL \i51/i591  (.A1(\i51/n54 ),
    .A2(\i51/n19 ),
    .B(\i51/n98 ),
    .Y(\i51/n582 ));
 INVx2_ASAP7_75t_SL \i51/i6  (.A(\i51/n545 ),
    .Y(\i51/n6 ));
 INVx1_ASAP7_75t_L \i51/i60  (.A(\i51/n400 ),
    .Y(\i51/n401 ));
 AND5x1_ASAP7_75t_SL \i51/i61  (.A(\i51/n322 ),
    .B(\i51/n581 ),
    .C(\i51/n314 ),
    .D(\i51/n246 ),
    .E(\i51/n223 ),
    .Y(\i51/n399 ));
 NOR3xp33_ASAP7_75t_SL \i51/i62  (.A(\i51/n332 ),
    .B(\i51/n313 ),
    .C(\i51/n297 ),
    .Y(\i51/n398 ));
 NOR3xp33_ASAP7_75t_SL \i51/i63  (.A(\i51/n355 ),
    .B(\i51/n298 ),
    .C(\i51/n256 ),
    .Y(\i51/n397 ));
 AND5x1_ASAP7_75t_SL \i51/i64  (.A(\i51/n288 ),
    .B(\i51/n300 ),
    .C(\i51/n575 ),
    .D(\i51/n291 ),
    .E(\i51/n229 ),
    .Y(\i51/n396 ));
 NOR2xp33_ASAP7_75t_SL \i51/i65  (.A(\i51/n356 ),
    .B(\i51/n361 ),
    .Y(\i51/n395 ));
 NAND5xp2_ASAP7_75t_SL \i51/i66  (.A(\i51/n321 ),
    .B(\i51/n282 ),
    .C(\i51/n196 ),
    .D(\i51/n183 ),
    .E(\i51/n265 ),
    .Y(\i51/n394 ));
 NOR4xp25_ASAP7_75t_SL \i51/i67  (.A(\i51/n311 ),
    .B(\i51/n553 ),
    .C(\i51/n269 ),
    .D(\i51/n249 ),
    .Y(\i51/n393 ));
 NAND4xp25_ASAP7_75t_SL \i51/i68  (.A(\i51/n329 ),
    .B(\i51/n463 ),
    .C(\i51/n342 ),
    .D(\i51/n346 ),
    .Y(\i51/n392 ));
 NAND4xp25_ASAP7_75t_SL \i51/i69  (.A(\i51/n353 ),
    .B(\i51/n351 ),
    .C(\i51/n556 ),
    .D(\i51/n222 ),
    .Y(\i51/n391 ));
 INVx2_ASAP7_75t_SL \i51/i7  (.A(\i51/n17 ),
    .Y(\i51/n7 ));
 NOR2x1_ASAP7_75t_SL \i51/i70  (.A(\i51/n175 ),
    .B(\i51/n382 ),
    .Y(\i51/n390 ));
 NAND3xp33_ASAP7_75t_SL \i51/i71  (.A(\i51/n346 ),
    .B(\i51/n320 ),
    .C(\i51/n22 ),
    .Y(\i51/n404 ));
 NAND4xp75_ASAP7_75t_SL \i51/i72  (.A(\i51/n480 ),
    .B(\i51/n236 ),
    .C(\i51/n307 ),
    .D(\i51/n25 ),
    .Y(\i51/n403 ));
 NAND2xp33_ASAP7_75t_L \i51/i73  (.A(\i51/n328 ),
    .B(\i51/n387 ),
    .Y(\i51/n389 ));
 AND2x2_ASAP7_75t_SL \i51/i74  (.A(\i51/n331 ),
    .B(\i51/n376 ),
    .Y(\i51/n402 ));
 NAND2x1p5_ASAP7_75t_SL \i51/i75  (.A(\i51/n384 ),
    .B(\i51/n341 ),
    .Y(\i51/n400 ));
 INVxp67_ASAP7_75t_SL \i51/i76  (.A(\i51/n387 ),
    .Y(\i51/n388 ));
 INVxp67_ASAP7_75t_SL \i51/i77  (.A(\i51/n381 ),
    .Y(\i51/n382 ));
 NOR5xp2_ASAP7_75t_SL \i51/i78  (.A(\i51/n564 ),
    .B(\i51/n255 ),
    .C(\i51/n521 ),
    .D(\i51/n540 ),
    .E(\i51/n560 ),
    .Y(\i51/n379 ));
 NOR3xp33_ASAP7_75t_SL \i51/i79  (.A(\i51/n350 ),
    .B(\i51/n273 ),
    .C(\i51/n562 ),
    .Y(\i51/n378 ));
 INVx2_ASAP7_75t_SL \i51/i8  (.A(\i51/n36 ),
    .Y(\i51/n8 ));
 NOR2xp33_ASAP7_75t_SL \i51/i80  (.A(\i51/n310 ),
    .B(\i51/n330 ),
    .Y(\i51/n377 ));
 NOR2xp33_ASAP7_75t_SL \i51/i81  (.A(\i51/n348 ),
    .B(\i51/n302 ),
    .Y(\i51/n376 ));
 NOR2x1_ASAP7_75t_SL \i51/i82  (.A(\i51/n315 ),
    .B(\i51/n289 ),
    .Y(\i51/n387 ));
 NAND3xp33_ASAP7_75t_SL \i51/i83  (.A(\i51/n264 ),
    .B(\i51/n287 ),
    .C(\i51/n535 ),
    .Y(\i51/n375 ));
 NAND2xp5_ASAP7_75t_L \i51/i84  (.A(\i51/n347 ),
    .B(\i51/n319 ),
    .Y(\i51/n374 ));
 NAND2xp5_ASAP7_75t_SL \i51/i85  (.A(\i51/n301 ),
    .B(\i51/n339 ),
    .Y(\i51/n373 ));
 NAND3xp33_ASAP7_75t_SL \i51/i86  (.A(\i51/n581 ),
    .B(\i51/n250 ),
    .C(\i51/n233 ),
    .Y(\i51/n386 ));
 NOR3xp33_ASAP7_75t_SL \i51/i87  (.A(\i51/n456 ),
    .B(\i51/n9 ),
    .C(\i51/n448 ),
    .Y(\i51/n372 ));
 NAND2xp5_ASAP7_75t_SL \i51/i88  (.A(\i51/n516 ),
    .B(\i51/n329 ),
    .Y(\i51/n385 ));
 OR3x1_ASAP7_75t_SL \i51/i89  (.A(\i51/n258 ),
    .B(\i51/n528 ),
    .C(\i51/n28 ),
    .Y(\i51/n371 ));
 NOR2x2_ASAP7_75t_SL \i51/i9  (.A(\i51/n443 ),
    .B(\i51/n442 ),
    .Y(n18[4]));
 NOR2x1_ASAP7_75t_SL \i51/i90  (.A(\i51/n562 ),
    .B(\i51/n350 ),
    .Y(\i51/n384 ));
 NOR2xp33_ASAP7_75t_L \i51/i91  (.A(\i51/n312 ),
    .B(\i51/n567 ),
    .Y(\i51/n383 ));
 NOR2xp33_ASAP7_75t_SL \i51/i92  (.A(\i51/n527 ),
    .B(\i51/n338 ),
    .Y(\i51/n381 ));
 NOR3x1_ASAP7_75t_SL \i51/i93  (.A(\i51/n263 ),
    .B(\i51/n569 ),
    .C(\i51/n305 ),
    .Y(\i51/n380 ));
 NOR3xp33_ASAP7_75t_SL \i51/i94  (.A(\i51/n270 ),
    .B(\i51/n195 ),
    .C(\i51/n261 ),
    .Y(\i51/n367 ));
 NOR2xp33_ASAP7_75t_SL \i51/i95  (.A(\i51/n580 ),
    .B(\i51/n325 ),
    .Y(\i51/n366 ));
 NAND3xp33_ASAP7_75t_SL \i51/i96  (.A(\i51/n257 ),
    .B(\i51/n317 ),
    .C(\i51/n268 ),
    .Y(\i51/n365 ));
 NAND4xp25_ASAP7_75t_SL \i51/i97  (.A(\i51/n241 ),
    .B(\i51/n254 ),
    .C(\i51/n278 ),
    .D(\i51/n511 ),
    .Y(\i51/n364 ));
 NAND2x1_ASAP7_75t_SL \i51/i98  (.A(\i51/n337 ),
    .B(\i51/n349 ),
    .Y(\i51/n370 ));
 NOR5xp2_ASAP7_75t_SL \i51/i99  (.A(\i51/n345 ),
    .B(\i51/n453 ),
    .C(\i51/n109 ),
    .D(\i51/n206 ),
    .E(\i51/n146 ),
    .Y(\i51/n363 ));
 AOI22xp5_ASAP7_75t_SL i510 (.A1(n530),
    .A2(n805),
    .B1(n529),
    .B2(n806),
    .Y(n962));
 XNOR2xp5_ASAP7_75t_SL i511 (.A(n309),
    .B(n308),
    .Y(n961));
 XOR2xp5_ASAP7_75t_SL i512 (.A(n311),
    .B(n310),
    .Y(n960));
 XNOR2xp5_ASAP7_75t_SL i513 (.A(n313),
    .B(n588),
    .Y(n959));
 XOR2xp5_ASAP7_75t_SL i514 (.A(n1168),
    .B(n590),
    .Y(n958));
 AOI22xp5_ASAP7_75t_SL i515 (.A1(n1181),
    .A2(n1210),
    .B1(n502),
    .B2(n534),
    .Y(n957));
 XOR2xp5_ASAP7_75t_SL i516 (.A(n316),
    .B(n606),
    .Y(n956));
 OAI22xp5_ASAP7_75t_SL i517 (.A1(n532),
    .A2(n509),
    .B1(n531),
    .B2(n508),
    .Y(n955));
 XOR2xp5_ASAP7_75t_SL i518 (.A(n318),
    .B(n593),
    .Y(n954));
 AOI22xp5_ASAP7_75t_SL i519 (.A1(n537),
    .A2(n492),
    .B1(n538),
    .B2(n493),
    .Y(n953));
 INVx2_ASAP7_75t_SL \i52/i0  (.A(n17[2]),
    .Y(\i52/n0 ));
 INVx2_ASAP7_75t_SL \i52/i1  (.A(n17[0]),
    .Y(\i52/n1 ));
 NOR2x1p5_ASAP7_75t_SL \i52/i10  (.A(\i52/n405 ),
    .B(\i52/n396 ),
    .Y(n16[5]));
 NOR5xp2_ASAP7_75t_SL \i52/i100  (.A(\i52/n246 ),
    .B(\i52/n456 ),
    .C(\i52/n233 ),
    .D(\i52/n193 ),
    .E(\i52/n156 ),
    .Y(\i52/n318 ));
 NAND5xp2_ASAP7_75t_SL \i52/i101  (.A(\i52/n421 ),
    .B(\i52/n258 ),
    .C(\i52/n512 ),
    .D(\i52/n429 ),
    .E(\i52/n511 ),
    .Y(\i52/n317 ));
 NAND3xp33_ASAP7_75t_L \i52/i102  (.A(\i52/n197 ),
    .B(\i52/n220 ),
    .C(\i52/n282 ),
    .Y(\i52/n316 ));
 NOR5xp2_ASAP7_75t_SL \i52/i103  (.A(\i52/n195 ),
    .B(\i52/n81 ),
    .C(\i52/n190 ),
    .D(\i52/n206 ),
    .E(\i52/n458 ),
    .Y(\i52/n315 ));
 NAND5xp2_ASAP7_75t_SL \i52/i104  (.A(\i52/n23 ),
    .B(\i52/n532 ),
    .C(\i52/n512 ),
    .D(\i52/n410 ),
    .E(\i52/n137 ),
    .Y(\i52/n314 ));
 NAND4xp25_ASAP7_75t_SL \i52/i105  (.A(\i52/n152 ),
    .B(\i52/n161 ),
    .C(\i52/n235 ),
    .D(\i52/n17 ),
    .Y(\i52/n313 ));
 NOR5xp2_ASAP7_75t_SL \i52/i106  (.A(\i52/n165 ),
    .B(\i52/n531 ),
    .C(\i52/n155 ),
    .D(\i52/n134 ),
    .E(\i52/n132 ),
    .Y(\i52/n312 ));
 NOR2xp33_ASAP7_75t_SL \i52/i107  (.A(\i52/n274 ),
    .B(\i52/n306 ),
    .Y(\i52/n311 ));
 NOR2xp33_ASAP7_75t_SL \i52/i108  (.A(\i52/n262 ),
    .B(\i52/n291 ),
    .Y(\i52/n310 ));
 NAND3x2_ASAP7_75t_SL \i52/i109  (.B(\i52/n258 ),
    .C(\i52/n289 ),
    .Y(\i52/n327 ),
    .A(\i52/n517 ));
 AND2x4_ASAP7_75t_SL \i52/i11  (.A(\i52/n406 ),
    .B(\i52/n389 ),
    .Y(n16[0]));
 NAND3x1_ASAP7_75t_SL \i52/i110  (.A(\i52/n254 ),
    .B(\i52/n236 ),
    .C(\i52/n211 ),
    .Y(\i52/n326 ));
 AOI21xp5_ASAP7_75t_L \i52/i111  (.A1(\i52/n447 ),
    .A2(\i52/n433 ),
    .B(\i52/n115 ),
    .Y(\i52/n302 ));
 NOR2xp33_ASAP7_75t_SL \i52/i112  (.A(\i52/n535 ),
    .B(\i52/n246 ),
    .Y(\i52/n301 ));
 NAND2xp5_ASAP7_75t_SL \i52/i113  (.A(\i52/n423 ),
    .B(\i52/n261 ),
    .Y(\i52/n300 ));
 NOR2xp33_ASAP7_75t_SL \i52/i114  (.A(\i52/n260 ),
    .B(\i52/n24 ),
    .Y(\i52/n299 ));
 NOR2xp33_ASAP7_75t_SL \i52/i115  (.A(\i52/n241 ),
    .B(\i52/n251 ),
    .Y(\i52/n298 ));
 NOR2xp67_ASAP7_75t_SL \i52/i116  (.A(\i52/n124 ),
    .B(\i52/n248 ),
    .Y(\i52/n297 ));
 NOR2xp33_ASAP7_75t_SL \i52/i117  (.A(\i52/n20 ),
    .B(\i52/n246 ),
    .Y(\i52/n296 ));
 NOR4xp25_ASAP7_75t_SL \i52/i118  (.A(\i52/n224 ),
    .B(\i52/n538 ),
    .C(\i52/n20 ),
    .D(\i52/n527 ),
    .Y(\i52/n295 ));
 NAND2xp5_ASAP7_75t_SL \i52/i119  (.A(\i52/n186 ),
    .B(\i52/n420 ),
    .Y(\i52/n294 ));
 NOR3xp33_ASAP7_75t_SL \i52/i12  (.A(\i52/n378 ),
    .B(\i52/n374 ),
    .C(\i52/n381 ),
    .Y(\i52/n406 ));
 NOR4xp25_ASAP7_75t_SL \i52/i120  (.A(\i52/n78 ),
    .B(\i52/n178 ),
    .C(\i52/n157 ),
    .D(\i52/n167 ),
    .Y(\i52/n293 ));
 NOR3xp33_ASAP7_75t_SL \i52/i121  (.A(\i52/n183 ),
    .B(\i52/n455 ),
    .C(\i52/n182 ),
    .Y(\i52/n292 ));
 NAND2xp33_ASAP7_75t_SL \i52/i122  (.A(\i52/n219 ),
    .B(\i52/n21 ),
    .Y(\i52/n291 ));
 NOR2xp33_ASAP7_75t_SL \i52/i123  (.A(\i52/n535 ),
    .B(\i52/n215 ),
    .Y(\i52/n290 ));
 NOR2x1p5_ASAP7_75t_SL \i52/i124  (.A(\i52/n201 ),
    .B(\i52/n506 ),
    .Y(\i52/n289 ));
 NAND2xp33_ASAP7_75t_SL \i52/i125  (.A(\i52/n259 ),
    .B(\i52/n244 ),
    .Y(\i52/n288 ));
 NAND3xp33_ASAP7_75t_SL \i52/i126  (.A(\i52/n22 ),
    .B(\i52/n151 ),
    .C(\i52/n450 ),
    .Y(\i52/n287 ));
 NOR3xp33_ASAP7_75t_SL \i52/i127  (.A(\i52/n547 ),
    .B(\i52/n162 ),
    .C(\i52/n143 ),
    .Y(\i52/n309 ));
 NAND2xp5_ASAP7_75t_SL \i52/i128  (.A(\i52/n223 ),
    .B(\i52/n152 ),
    .Y(\i52/n308 ));
 NOR2x1_ASAP7_75t_SL \i52/i129  (.A(\i52/n200 ),
    .B(\i52/n217 ),
    .Y(\i52/n307 ));
 NOR2x2_ASAP7_75t_SL \i52/i13  (.A(\i52/n398 ),
    .B(\i52/n399 ),
    .Y(n16[2]));
 NAND2xp5_ASAP7_75t_SL \i52/i130  (.A(\i52/n512 ),
    .B(\i52/n225 ),
    .Y(\i52/n306 ));
 NOR2x1_ASAP7_75t_SL \i52/i131  (.A(\i52/n202 ),
    .B(\i52/n249 ),
    .Y(\i52/n305 ));
 NOR2x1_ASAP7_75t_SL \i52/i132  (.A(\i52/n538 ),
    .B(\i52/n535 ),
    .Y(\i52/n304 ));
 NOR3x1_ASAP7_75t_SL \i52/i133  (.A(\i52/n155 ),
    .B(\i52/n572 ),
    .C(\i52/n131 ),
    .Y(\i52/n303 ));
 INVx1_ASAP7_75t_SL \i52/i134  (.A(\i52/n284 ),
    .Y(\i52/n285 ));
 INVx1_ASAP7_75t_SL \i52/i135  (.A(\i52/n25 ),
    .Y(\i52/n283 ));
 NOR4xp25_ASAP7_75t_SL \i52/i136  (.A(\i52/n475 ),
    .B(\i52/n169 ),
    .C(\i52/n160 ),
    .D(\i52/n141 ),
    .Y(\i52/n282 ));
 AOI211xp5_ASAP7_75t_SL \i52/i137  (.A1(\i52/n83 ),
    .A2(\i52/n43 ),
    .B(\i52/n232 ),
    .C(\i52/n181 ),
    .Y(\i52/n281 ));
 NAND2xp33_ASAP7_75t_SL \i52/i138  (.A(\i52/n212 ),
    .B(\i52/n231 ),
    .Y(\i52/n280 ));
 NAND5xp2_ASAP7_75t_SL \i52/i139  (.A(\i52/n493 ),
    .B(\i52/n177 ),
    .C(\i52/n188 ),
    .D(\i52/n487 ),
    .E(\i52/n522 ),
    .Y(\i52/n279 ));
 NAND4xp25_ASAP7_75t_SL \i52/i14  (.A(\i52/n364 ),
    .B(\i52/n384 ),
    .C(\i52/n362 ),
    .D(\i52/n573 ),
    .Y(\i52/n405 ));
 NOR4xp25_ASAP7_75t_SL \i52/i140  (.A(\i52/n238 ),
    .B(\i52/n104 ),
    .C(\i52/n548 ),
    .D(\i52/n121 ),
    .Y(\i52/n278 ));
 NOR2xp33_ASAP7_75t_SL \i52/i141  (.A(\i52/n207 ),
    .B(\i52/n540 ),
    .Y(\i52/n277 ));
 AOI211xp5_ASAP7_75t_SL \i52/i142  (.A1(\i52/n119 ),
    .A2(\i52/n52 ),
    .B(\i52/n473 ),
    .C(\i52/n135 ),
    .Y(\i52/n276 ));
 OA21x2_ASAP7_75t_SL \i52/i143  (.A1(\i52/n45 ),
    .A2(\i52/n447 ),
    .B(\i52/n532 ),
    .Y(\i52/n275 ));
 NAND5xp2_ASAP7_75t_SL \i52/i144  (.A(\i52/n105 ),
    .B(\i52/n491 ),
    .C(\i52/n414 ),
    .D(\i52/n436 ),
    .E(\i52/n65 ),
    .Y(\i52/n274 ));
 NOR3xp33_ASAP7_75t_SL \i52/i145  (.A(\i52/n218 ),
    .B(\i52/n549 ),
    .C(\i52/n64 ),
    .Y(\i52/n273 ));
 NAND2xp5_ASAP7_75t_SL \i52/i146  (.A(\i52/n205 ),
    .B(\i52/n23 ),
    .Y(\i52/n272 ));
 NAND5xp2_ASAP7_75t_SL \i52/i147  (.A(\i52/n497 ),
    .B(\i52/n72 ),
    .C(\i52/n147 ),
    .D(\i52/n140 ),
    .E(\i52/n488 ),
    .Y(\i52/n271 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i52/i148  (.A1(\i52/n54 ),
    .A2(\i52/n66 ),
    .B(\i52/n444 ),
    .C(\i52/n198 ),
    .Y(\i52/n270 ));
 NAND4xp25_ASAP7_75t_SL \i52/i149  (.A(\i52/n229 ),
    .B(\i52/n557 ),
    .C(\i52/n79 ),
    .D(\i52/n129 ),
    .Y(\i52/n269 ));
 NOR3xp33_ASAP7_75t_SL \i52/i15  (.A(\i52/n382 ),
    .B(\i52/n347 ),
    .C(\i52/n392 ),
    .Y(\i52/n404 ));
 NAND5xp2_ASAP7_75t_SL \i52/i150  (.A(\i52/n120 ),
    .B(\i52/n106 ),
    .C(\i52/n171 ),
    .D(\i52/n75 ),
    .E(\i52/n70 ),
    .Y(\i52/n268 ));
 NAND2xp5_ASAP7_75t_SL \i52/i151  (.A(\i52/n204 ),
    .B(\i52/n222 ),
    .Y(\i52/n267 ));
 NAND3xp33_ASAP7_75t_SL \i52/i152  (.A(\i52/n216 ),
    .B(\i52/n499 ),
    .C(\i52/n67 ),
    .Y(\i52/n266 ));
 NAND2xp5_ASAP7_75t_SL \i52/i153  (.A(\i52/n517 ),
    .B(\i52/n258 ),
    .Y(\i52/n265 ));
 NOR2xp33_ASAP7_75t_L \i52/i154  (.A(\i52/n239 ),
    .B(\i52/n251 ),
    .Y(\i52/n286 ));
 NAND2xp5_ASAP7_75t_SL \i52/i155  (.A(\i52/n516 ),
    .B(\i52/n259 ),
    .Y(\i52/n264 ));
 NOR2x1p5_ASAP7_75t_SL \i52/i156  (.A(\i52/n470 ),
    .B(\i52/n243 ),
    .Y(\i52/n284 ));
 NAND3x1_ASAP7_75t_SL \i52/i157  (.A(\i52/n192 ),
    .B(\i52/n518 ),
    .C(\i52/n419 ),
    .Y(\i52/n25 ));
 INVxp67_ASAP7_75t_SL \i52/i158  (.A(\i52/n262 ),
    .Y(\i52/n263 ));
 INVxp67_ASAP7_75t_SL \i52/i159  (.A(\i52/n7 ),
    .Y(\i52/n261 ));
 NAND4xp75_ASAP7_75t_SL \i52/i16  (.A(\i52/n363 ),
    .B(\i52/n394 ),
    .C(\i52/n368 ),
    .D(\i52/n358 ),
    .Y(\i52/n403 ));
 INVxp67_ASAP7_75t_SL \i52/i160  (.A(\i52/n461 ),
    .Y(\i52/n257 ));
 INVxp67_ASAP7_75t_SL \i52/i161  (.A(\i52/n255 ),
    .Y(\i52/n256 ));
 INVx1_ASAP7_75t_SL \i52/i162  (.A(\i52/n253 ),
    .Y(\i52/n254 ));
 INVxp67_ASAP7_75t_SL \i52/i163  (.A(\i52/n482 ),
    .Y(\i52/n252 ));
 INVxp67_ASAP7_75t_SL \i52/i164  (.A(\i52/n249 ),
    .Y(\i52/n250 ));
 INVxp67_ASAP7_75t_SL \i52/i165  (.A(\i52/n533 ),
    .Y(\i52/n247 ));
 INVx1_ASAP7_75t_SL \i52/i166  (.A(\i52/n244 ),
    .Y(\i52/n245 ));
 NAND2x1_ASAP7_75t_SL \i52/i167  (.A(\i52/n417 ),
    .B(\i52/n159 ),
    .Y(\i52/n243 ));
 NOR2xp33_ASAP7_75t_SL \i52/i168  (.A(\i52/n189 ),
    .B(\i52/n183 ),
    .Y(\i52/n242 ));
 NAND2xp33_ASAP7_75t_SL \i52/i169  (.A(\i52/n151 ),
    .B(\i52/n512 ),
    .Y(\i52/n241 ));
 AND3x4_ASAP7_75t_SL \i52/i17  (.A(\i52/n385 ),
    .B(\i52/n400 ),
    .C(\i52/n390 ),
    .Y(n16[7]));
 OAI21xp33_ASAP7_75t_SL \i52/i170  (.A1(\i52/n42 ),
    .A2(\i52/n426 ),
    .B(\i52/n139 ),
    .Y(\i52/n240 ));
 NAND2xp5_ASAP7_75t_SL \i52/i171  (.A(\i52/n130 ),
    .B(\i52/n151 ),
    .Y(\i52/n239 ));
 AOI31xp33_ASAP7_75t_SL \i52/i172  (.A1(\i52/n42 ),
    .A2(\i52/n415 ),
    .A3(\i52/n480 ),
    .B(\i52/n36 ),
    .Y(\i52/n238 ));
 NOR3xp33_ASAP7_75t_SL \i52/i173  (.A(\i52/n455 ),
    .B(\i52/n98 ),
    .C(\i52/n87 ),
    .Y(\i52/n237 ));
 NOR3xp33_ASAP7_75t_SL \i52/i174  (.A(\i52/n521 ),
    .B(\i52/n94 ),
    .C(\i52/n189 ),
    .Y(\i52/n236 ));
 OAI31xp33_ASAP7_75t_SL \i52/i175  (.A1(\i52/n38 ),
    .A2(\i52/n39 ),
    .A3(\i52/n51 ),
    .B(\i52/n59 ),
    .Y(\i52/n235 ));
 OAI31xp33_ASAP7_75t_SL \i52/i176  (.A1(\i52/n52 ),
    .A2(\i52/n53 ),
    .A3(\i52/n54 ),
    .B(\i52/n51 ),
    .Y(\i52/n234 ));
 AOI21xp5_ASAP7_75t_SL \i52/i177  (.A1(\i52/n115 ),
    .A2(\i52/n480 ),
    .B(\i52/n427 ),
    .Y(\i52/n262 ));
 OAI221xp5_ASAP7_75t_SL \i52/i178  (.A1(\i52/n16 ),
    .A2(\i52/n61 ),
    .B1(\i52/n460 ),
    .B2(\i52/n496 ),
    .C(\i52/n434 ),
    .Y(\i52/n233 ));
 AOI21xp33_ASAP7_75t_SL \i52/i179  (.A1(\i52/n125 ),
    .A2(\i52/n37 ),
    .B(\i52/n445 ),
    .Y(\i52/n232 ));
 NAND4xp75_ASAP7_75t_SL \i52/i18  (.A(\i52/n576 ),
    .B(\i52/n367 ),
    .C(\i52/n376 ),
    .D(\i52/n393 ),
    .Y(\i52/n402 ));
 NOR3xp33_ASAP7_75t_SL \i52/i180  (.A(\i52/n166 ),
    .B(\i52/n521 ),
    .C(\i52/n103 ),
    .Y(\i52/n231 ));
 NAND3xp33_ASAP7_75t_SL \i52/i181  (.A(\i52/n408 ),
    .B(\i52/n479 ),
    .C(\i52/n123 ),
    .Y(\i52/n230 ));
 OAI21xp5_ASAP7_75t_SL \i52/i182  (.A1(\i52/n47 ),
    .A2(\i52/n117 ),
    .B(\i52/n52 ),
    .Y(\i52/n229 ));
 NAND4xp25_ASAP7_75t_SL \i52/i183  (.A(\i52/n133 ),
    .B(\i52/n129 ),
    .C(\i52/n563 ),
    .D(\i52/n108 ),
    .Y(\i52/n228 ));
 NAND2xp33_ASAP7_75t_SL \i52/i184  (.A(\i52/n174 ),
    .B(\i52/n102 ),
    .Y(\i52/n227 ));
 OAI211xp5_ASAP7_75t_SL \i52/i185  (.A1(\i52/n50 ),
    .A2(\i52/n445 ),
    .B(\i52/n435 ),
    .C(\i52/n492 ),
    .Y(\i52/n260 ));
 NOR2xp67_ASAP7_75t_SL \i52/i186  (.A(\i52/n530 ),
    .B(\i52/n190 ),
    .Y(\i52/n259 ));
 AOI21x1_ASAP7_75t_SL \i52/i187  (.A1(\i52/n44 ),
    .A2(\i52/n47 ),
    .B(\i52/n473 ),
    .Y(\i52/n258 ));
 NAND2xp5_ASAP7_75t_SL \i52/i188  (.A(\i52/n494 ),
    .B(\i52/n513 ),
    .Y(\i52/n24 ));
 OAI211xp5_ASAP7_75t_SL \i52/i189  (.A1(\i52/n480 ),
    .A2(\i52/n445 ),
    .B(\i52/n139 ),
    .C(\i52/n562 ),
    .Y(\i52/n255 ));
 NAND2x1_ASAP7_75t_SL \i52/i19  (.A(\i52/n355 ),
    .B(\i52/n386 ),
    .Y(\i52/n401 ));
 OR2x2_ASAP7_75t_SL \i52/i190  (.A(\i52/n474 ),
    .B(\i52/n537 ),
    .Y(\i52/n253 ));
 NAND2xp5_ASAP7_75t_SL \i52/i191  (.A(\i52/n511 ),
    .B(\i52/n191 ),
    .Y(\i52/n251 ));
 NAND2xp5_ASAP7_75t_SL \i52/i192  (.A(\i52/n22 ),
    .B(\i52/n413 ),
    .Y(\i52/n249 ));
 NAND2xp5_ASAP7_75t_SL \i52/i193  (.A(\i52/n173 ),
    .B(\i52/n509 ),
    .Y(\i52/n248 ));
 NAND2xp5_ASAP7_75t_SL \i52/i194  (.A(\i52/n437 ),
    .B(\i52/n503 ),
    .Y(\i52/n246 ));
 NOR2x1_ASAP7_75t_SL \i52/i195  (.A(\i52/n175 ),
    .B(\i52/n156 ),
    .Y(\i52/n244 ));
 INVxp67_ASAP7_75t_SL \i52/i196  (.A(\i52/n224 ),
    .Y(\i52/n225 ));
 INVx1_ASAP7_75t_SL \i52/i197  (.A(\i52/n220 ),
    .Y(\i52/n221 ));
 INVx1_ASAP7_75t_SL \i52/i198  (.A(\i52/n216 ),
    .Y(\i52/n217 ));
 NAND4xp25_ASAP7_75t_SL \i52/i199  (.A(\i52/n80 ),
    .B(\i52/n407 ),
    .C(\i52/n84 ),
    .D(\i52/n501 ),
    .Y(\i52/n214 ));
 INVx2_ASAP7_75t_SL \i52/i2  (.A(\i52/n523 ),
    .Y(\i52/n2 ));
 NOR2xp67_ASAP7_75t_SL \i52/i20  (.A(\i52/n387 ),
    .B(\i52/n348 ),
    .Y(\i52/n400 ));
 AOI31xp33_ASAP7_75t_SL \i52/i200  (.A1(\i52/n566 ),
    .A2(\i52/n447 ),
    .A3(\i52/n36 ),
    .B(\i52/n37 ),
    .Y(\i52/n213 ));
 NOR4xp25_ASAP7_75t_SL \i52/i201  (.A(\i52/n78 ),
    .B(\i52/n476 ),
    .C(\i52/n138 ),
    .D(\i52/n63 ),
    .Y(\i52/n212 ));
 AOI211xp5_ASAP7_75t_SL \i52/i202  (.A1(\i52/n96 ),
    .A2(\i52/n443 ),
    .B(\i52/n549 ),
    .C(\i52/n68 ),
    .Y(\i52/n211 ));
 NOR2xp33_ASAP7_75t_L \i52/i203  (.A(\i52/n529 ),
    .B(\i52/n184 ),
    .Y(\i52/n210 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i52/i204  (.A1(\i52/n445 ),
    .A2(\i52/n40 ),
    .B(\i52/n58 ),
    .C(\i52/n560 ),
    .Y(\i52/n209 ));
 NOR2xp33_ASAP7_75t_SL \i52/i205  (.A(\i52/n546 ),
    .B(\i52/n144 ),
    .Y(\i52/n208 ));
 NAND2xp33_ASAP7_75t_L \i52/i206  (.A(\i52/n77 ),
    .B(\i52/n150 ),
    .Y(\i52/n207 ));
 NAND2xp33_ASAP7_75t_SL \i52/i207  (.A(\i52/n180 ),
    .B(\i52/n489 ),
    .Y(\i52/n206 ));
 AOI22xp5_ASAP7_75t_SL \i52/i208  (.A1(\i52/n53 ),
    .A2(\i52/n74 ),
    .B1(\i52/n443 ),
    .B2(\i52/n54 ),
    .Y(\i52/n205 ));
 OAI21xp5_ASAP7_75t_SL \i52/i209  (.A1(\i52/n83 ),
    .A2(\i52/n53 ),
    .B(\i52/n443 ),
    .Y(\i52/n204 ));
 NAND4xp75_ASAP7_75t_SL \i52/i21  (.A(\i52/n359 ),
    .B(\i52/n371 ),
    .C(\i52/n353 ),
    .D(\i52/n356 ),
    .Y(\i52/n399 ));
 OA21x2_ASAP7_75t_SL \i52/i210  (.A1(\i52/n37 ),
    .A2(\i52/n426 ),
    .B(\i52/n91 ),
    .Y(\i52/n203 ));
 NAND2xp5_ASAP7_75t_SL \i52/i211  (.A(\i52/n146 ),
    .B(\i52/n194 ),
    .Y(\i52/n202 ));
 NAND4xp25_ASAP7_75t_SL \i52/i212  (.A(\i52/n438 ),
    .B(\i52/n109 ),
    .C(\i52/n71 ),
    .D(\i52/n565 ),
    .Y(\i52/n201 ));
 OAI221xp5_ASAP7_75t_SL \i52/i213  (.A1(\i52/n60 ),
    .A2(\i52/n58 ),
    .B1(\i52/n556 ),
    .B2(\i52/n569 ),
    .C(\i52/n76 ),
    .Y(\i52/n226 ));
 OAI222xp33_ASAP7_75t_SL \i52/i214  (.A1(\i52/n498 ),
    .A2(\i52/n42 ),
    .B1(\i52/n496 ),
    .B2(\i52/n50 ),
    .C1(\i52/n556 ),
    .C2(\i52/n55 ),
    .Y(\i52/n200 ));
 AND3x1_ASAP7_75t_SL \i52/i215  (.A(\i52/n90 ),
    .B(\i52/n407 ),
    .C(\i52/n559 ),
    .Y(\i52/n199 ));
 NAND2xp33_ASAP7_75t_SL \i52/i216  (.A(\i52/n148 ),
    .B(\i52/n170 ),
    .Y(\i52/n198 ));
 NAND3x1_ASAP7_75t_SL \i52/i217  (.A(\i52/n561 ),
    .B(\i52/n110 ),
    .C(\i52/n107 ),
    .Y(\i52/n224 ));
 AOI22xp5_ASAP7_75t_SL \i52/i218  (.A1(\i52/n571 ),
    .A2(\i52/n59 ),
    .B1(\i52/n51 ),
    .B2(\i52/n534 ),
    .Y(\i52/n223 ));
 AOI22xp5_ASAP7_75t_SL \i52/i219  (.A1(\i52/n62 ),
    .A2(\i52/n457 ),
    .B1(\i52/n38 ),
    .B2(\i52/n52 ),
    .Y(\i52/n222 ));
 OR3x1_ASAP7_75t_SL \i52/i22  (.A(\i52/n379 ),
    .B(\i52/n377 ),
    .C(\i52/n360 ),
    .Y(\i52/n398 ));
 AOI221x1_ASAP7_75t_SL \i52/i220  (.A1(\i52/n59 ),
    .A2(\i52/n51 ),
    .B1(\i52/n54 ),
    .B2(\i52/n444 ),
    .C(\i52/n432 ),
    .Y(\i52/n220 ));
 AOI211x1_ASAP7_75t_SL \i52/i221  (.A1(\i52/n69 ),
    .A2(\i52/n48 ),
    .B(\i52/n564 ),
    .C(\i52/n138 ),
    .Y(\i52/n219 ));
 OAI21xp5_ASAP7_75t_SL \i52/i222  (.A1(\i52/n36 ),
    .A2(\i52/n58 ),
    .B(\i52/n422 ),
    .Y(\i52/n218 ));
 NOR2x1_ASAP7_75t_SL \i52/i223  (.A(\i52/n92 ),
    .B(\i52/n545 ),
    .Y(\i52/n216 ));
 OAI211xp5_ASAP7_75t_SL \i52/i224  (.A1(\i52/n459 ),
    .A2(\i52/n505 ),
    .B(\i52/n79 ),
    .C(\i52/n510 ),
    .Y(\i52/n215 ));
 NOR2xp33_ASAP7_75t_SL \i52/i225  (.A(\i52/n99 ),
    .B(\i52/n149 ),
    .Y(\i52/n23 ));
 NOR2xp33_ASAP7_75t_SL \i52/i226  (.A(\i52/n100 ),
    .B(\i52/n543 ),
    .Y(\i52/n197 ));
 INVx1_ASAP7_75t_SL \i52/i227  (.A(\i52/n509 ),
    .Y(\i52/n195 ));
 INVx1_ASAP7_75t_SL \i52/i228  (.A(\i52/n193 ),
    .Y(\i52/n194 ));
 INVx1_ASAP7_75t_SL \i52/i229  (.A(\i52/n543 ),
    .Y(\i52/n192 ));
 OR3x1_ASAP7_75t_SL \i52/i23  (.A(\i52/n380 ),
    .B(\i52/n346 ),
    .C(\i52/n320 ),
    .Y(\i52/n397 ));
 INVxp67_ASAP7_75t_SL \i52/i230  (.A(\i52/n187 ),
    .Y(\i52/n188 ));
 INVx1_ASAP7_75t_SL \i52/i231  (.A(\i52/n184 ),
    .Y(\i52/n185 ));
 OAI21xp33_ASAP7_75t_SL \i52/i232  (.A1(\i52/n550 ),
    .A2(\i52/n446 ),
    .B(\i52/n555 ),
    .Y(\i52/n182 ));
 NAND2xp5_ASAP7_75t_SL \i52/i233  (.A(\i52/n500 ),
    .B(\i52/n95 ),
    .Y(\i52/n181 ));
 OAI21xp5_ASAP7_75t_SL \i52/i234  (.A1(\i52/n534 ),
    .A2(\i52/n44 ),
    .B(\i52/n441 ),
    .Y(\i52/n180 ));
 NOR2xp33_ASAP7_75t_SL \i52/i235  (.A(\i52/n101 ),
    .B(\i52/n416 ),
    .Y(\i52/n179 ));
 NAND2xp33_ASAP7_75t_L \i52/i236  (.A(\i52/n502 ),
    .B(\i52/n490 ),
    .Y(\i52/n178 ));
 NOR2xp33_ASAP7_75t_SL \i52/i237  (.A(\i52/n18 ),
    .B(\i52/n85 ),
    .Y(\i52/n177 ));
 OAI21xp5_ASAP7_75t_SL \i52/i238  (.A1(\i52/n45 ),
    .A2(\i52/n427 ),
    .B(\i52/n127 ),
    .Y(\i52/n176 ));
 OAI21xp5_ASAP7_75t_SL \i52/i239  (.A1(\i52/n415 ),
    .A2(\i52/n556 ),
    .B(\i52/n97 ),
    .Y(\i52/n175 ));
 NAND3xp33_ASAP7_75t_SL \i52/i24  (.A(\i52/n391 ),
    .B(\i52/n376 ),
    .C(\i52/n359 ),
    .Y(\i52/n396 ));
 OAI21xp5_ASAP7_75t_SL \i52/i240  (.A1(\i52/n53 ),
    .A2(\i52/n44 ),
    .B(\i52/n49 ),
    .Y(\i52/n174 ));
 AOI22xp5_ASAP7_75t_SL \i52/i241  (.A1(\i52/n35 ),
    .A2(\i52/n62 ),
    .B1(\i52/n38 ),
    .B2(\i52/n53 ),
    .Y(\i52/n173 ));
 OA21x2_ASAP7_75t_SL \i52/i242  (.A1(\i52/n448 ),
    .A2(\i52/n15 ),
    .B(\i52/n487 ),
    .Y(\i52/n196 ));
 AOI21xp33_ASAP7_75t_SL \i52/i243  (.A1(\i52/n50 ),
    .A2(\i52/n448 ),
    .B(\i52/n36 ),
    .Y(\i52/n172 ));
 OAI21xp5_ASAP7_75t_SL \i52/i244  (.A1(\i52/n444 ),
    .A2(\i52/n62 ),
    .B(\i52/n467 ),
    .Y(\i52/n171 ));
 OAI21xp33_ASAP7_75t_SL \i52/i245  (.A1(\i52/n49 ),
    .A2(\i52/n38 ),
    .B(\i52/n467 ),
    .Y(\i52/n170 ));
 AOI21xp33_ASAP7_75t_SL \i52/i246  (.A1(\i52/n480 ),
    .A2(\i52/n58 ),
    .B(\i52/n36 ),
    .Y(\i52/n169 ));
 OAI21xp5_ASAP7_75t_SL \i52/i247  (.A1(\i52/n45 ),
    .A2(\i52/n556 ),
    .B(\i52/n21 ),
    .Y(\i52/n168 ));
 AOI21xp33_ASAP7_75t_SL \i52/i248  (.A1(\i52/n445 ),
    .A2(\i52/n36 ),
    .B(\i52/n459 ),
    .Y(\i52/n167 ));
 NAND2xp5_ASAP7_75t_SL \i52/i249  (.A(\i52/n467 ),
    .B(\i52/n116 ),
    .Y(\i52/n22 ));
 NOR2x1_ASAP7_75t_SL \i52/i25  (.A(\i52/n300 ),
    .B(\i52/n377 ),
    .Y(\i52/n394 ));
 NAND2xp5_ASAP7_75t_L \i52/i250  (.A(\i52/n139 ),
    .B(\i52/n562 ),
    .Y(\i52/n166 ));
 OAI22xp5_ASAP7_75t_L \i52/i251  (.A1(\i52/n515 ),
    .A2(\i52/n556 ),
    .B1(\i52/n16 ),
    .B2(\i52/n50 ),
    .Y(\i52/n193 ));
 AOI22xp5_ASAP7_75t_SL \i52/i252  (.A1(\i52/n48 ),
    .A2(\i52/n59 ),
    .B1(\i52/n5 ),
    .B2(\i52/n57 ),
    .Y(\i52/n191 ));
 OAI22xp5_ASAP7_75t_SL \i52/i253  (.A1(\i52/n515 ),
    .A2(\i52/n60 ),
    .B1(\i52/n37 ),
    .B2(\i52/n498 ),
    .Y(\i52/n190 ));
 NAND2xp33_ASAP7_75t_SL \i52/i254  (.A(\i52/n17 ),
    .B(\i52/n112 ),
    .Y(\i52/n189 ));
 OAI22xp5_ASAP7_75t_SL \i52/i255  (.A1(\i52/n45 ),
    .A2(\i52/n60 ),
    .B1(\i52/n50 ),
    .B2(\i52/n427 ),
    .Y(\i52/n187 ));
 OAI21xp5_ASAP7_75t_SL \i52/i256  (.A1(\i52/n53 ),
    .A2(\i52/n41 ),
    .B(\i52/n441 ),
    .Y(\i52/n186 ));
 NOR2xp33_ASAP7_75t_L \i52/i257  (.A(\i52/n15 ),
    .B(\i52/n484 ),
    .Y(\i52/n184 ));
 NAND2xp33_ASAP7_75t_L \i52/i258  (.A(\i52/n79 ),
    .B(\i52/n510 ),
    .Y(\i52/n165 ));
 OAI21xp33_ASAP7_75t_SL \i52/i259  (.A1(\i52/n459 ),
    .A2(\i52/n496 ),
    .B(\i52/n522 ),
    .Y(\i52/n183 ));
 NOR2x1_ASAP7_75t_SL \i52/i26  (.A(\i52/n361 ),
    .B(\i52/n357 ),
    .Y(\i52/n393 ));
 INVxp67_ASAP7_75t_SL \i52/i260  (.A(\i52/n163 ),
    .Y(\i52/n164 ));
 INVxp67_ASAP7_75t_SL \i52/i261  (.A(\i52/n161 ),
    .Y(\i52/n162 ));
 INVxp67_ASAP7_75t_SL \i52/i262  (.A(\i52/n417 ),
    .Y(\i52/n160 ));
 INVx1_ASAP7_75t_SL \i52/i263  (.A(\i52/n158 ),
    .Y(\i52/n159 ));
 INVxp67_ASAP7_75t_SL \i52/i264  (.A(\i52/n434 ),
    .Y(\i52/n157 ));
 INVxp67_ASAP7_75t_SL \i52/i265  (.A(\i52/n546 ),
    .Y(\i52/n154 ));
 INVxp67_ASAP7_75t_SL \i52/i266  (.A(\i52/n547 ),
    .Y(\i52/n153 ));
 OAI21xp5_ASAP7_75t_SL \i52/i267  (.A1(\i52/n534 ),
    .A2(\i52/n41 ),
    .B(\i52/n46 ),
    .Y(\i52/n150 ));
 OAI22xp5_ASAP7_75t_SL \i52/i268  (.A1(\i52/n60 ),
    .A2(\i52/n42 ),
    .B1(\i52/n460 ),
    .B2(\i52/n15 ),
    .Y(\i52/n149 ));
 OAI21xp5_ASAP7_75t_SL \i52/i269  (.A1(\i52/n35 ),
    .A2(\i52/n41 ),
    .B(\i52/n39 ),
    .Y(\i52/n148 ));
 NAND3xp33_ASAP7_75t_SL \i52/i27  (.A(\i52/n341 ),
    .B(\i52/n580 ),
    .C(\i52/n339 ),
    .Y(\i52/n392 ));
 OAI21xp5_ASAP7_75t_SL \i52/i270  (.A1(\i52/n443 ),
    .A2(\i52/n46 ),
    .B(\i52/n534 ),
    .Y(\i52/n147 ));
 AOI22xp33_ASAP7_75t_SL \i52/i271  (.A1(\i52/n48 ),
    .A2(\i52/n53 ),
    .B1(\i52/n5 ),
    .B2(\i52/n534 ),
    .Y(\i52/n146 ));
 OAI22xp5_ASAP7_75t_SL \i52/i272  (.A1(\i52/n480 ),
    .A2(\i52/n498 ),
    .B1(\i52/n58 ),
    .B2(\i52/n445 ),
    .Y(\i52/n145 ));
 OAI22xp33_ASAP7_75t_SL \i52/i273  (.A1(\i52/n40 ),
    .A2(\i52/n446 ),
    .B1(\i52/n15 ),
    .B2(\i52/n42 ),
    .Y(\i52/n144 ));
 OAI22xp5_ASAP7_75t_SL \i52/i274  (.A1(\i52/n446 ),
    .A2(\i52/n60 ),
    .B1(\i52/n50 ),
    .B2(\i52/n15 ),
    .Y(\i52/n143 ));
 OAI21xp5_ASAP7_75t_SL \i52/i275  (.A1(\i52/n37 ),
    .A2(\i52/n496 ),
    .B(\i52/n86 ),
    .Y(\i52/n163 ));
 AOI22xp5_ASAP7_75t_SL \i52/i276  (.A1(\i52/n35 ),
    .A2(\i52/n49 ),
    .B1(\i52/n38 ),
    .B2(\i52/n44 ),
    .Y(\i52/n161 ));
 OAI22xp5_ASAP7_75t_SL \i52/i277  (.A1(\i52/n36 ),
    .A2(\i52/n569 ),
    .B1(\i52/n446 ),
    .B2(\i52/n447 ),
    .Y(\i52/n142 ));
 NAND2xp33_ASAP7_75t_SL \i52/i278  (.A(\i52/n488 ),
    .B(\i52/n140 ),
    .Y(\i52/n141 ));
 OAI22xp5_ASAP7_75t_SL \i52/i279  (.A1(\i52/n415 ),
    .A2(\i52/n60 ),
    .B1(\i52/n550 ),
    .B2(\i52/n460 ),
    .Y(\i52/n158 ));
 NOR2xp33_ASAP7_75t_L \i52/i28  (.A(\i52/n366 ),
    .B(\i52/n329 ),
    .Y(\i52/n391 ));
 AO22x2_ASAP7_75t_SL \i52/i280  (.A1(\i52/n62 ),
    .A2(\i52/n59 ),
    .B1(\i52/n43 ),
    .B2(\i52/n57 ),
    .Y(\i52/n156 ));
 OAI21xp5_ASAP7_75t_SL \i52/i281  (.A1(\i52/n55 ),
    .A2(\i52/n40 ),
    .B(\i52/n73 ),
    .Y(\i52/n155 ));
 AOI22xp5_ASAP7_75t_SL \i52/i282  (.A1(\i52/n35 ),
    .A2(\i52/n39 ),
    .B1(\i52/n51 ),
    .B2(\i52/n57 ),
    .Y(\i52/n152 ));
 AOI22xp5_ASAP7_75t_SL \i52/i283  (.A1(\i52/n46 ),
    .A2(\i52/n57 ),
    .B1(\i52/n38 ),
    .B2(\i52/n454 ),
    .Y(\i52/n151 ));
 INVxp67_ASAP7_75t_SL \i52/i284  (.A(\i52/n564 ),
    .Y(\i52/n137 ));
 INVx1_ASAP7_75t_SL \i52/i285  (.A(\i52/n514 ),
    .Y(\i52/n136 ));
 INVxp67_ASAP7_75t_SL \i52/i286  (.A(\i52/n437 ),
    .Y(\i52/n135 ));
 INVxp67_ASAP7_75t_SL \i52/i287  (.A(\i52/n133 ),
    .Y(\i52/n134 ));
 INVxp67_ASAP7_75t_SL \i52/i288  (.A(\i52/n555 ),
    .Y(\i52/n132 ));
 INVxp67_ASAP7_75t_SL \i52/i289  (.A(\i52/n527 ),
    .Y(\i52/n130 ));
 NOR5xp2_ASAP7_75t_SL \i52/i29  (.A(\i52/n331 ),
    .B(\i52/n279 ),
    .C(\i52/n322 ),
    .D(\i52/n248 ),
    .E(\i52/n541 ),
    .Y(\i52/n390 ));
 INVxp67_ASAP7_75t_SL \i52/i290  (.A(\i52/n127 ),
    .Y(\i52/n128 ));
 INVxp67_ASAP7_75t_SL \i52/i291  (.A(\i52/n502 ),
    .Y(\i52/n126 ));
 INVxp67_ASAP7_75t_SL \i52/i292  (.A(\i52/n123 ),
    .Y(\i52/n124 ));
 INVxp67_ASAP7_75t_SL \i52/i293  (.A(\i52/n425 ),
    .Y(\i52/n122 ));
 INVxp67_ASAP7_75t_SL \i52/i294  (.A(\i52/n120 ),
    .Y(\i52/n121 ));
 INVxp67_ASAP7_75t_SL \i52/i295  (.A(\i52/n118 ),
    .Y(\i52/n119 ));
 INVxp67_ASAP7_75t_SL \i52/i296  (.A(\i52/n484 ),
    .Y(\i52/n117 ));
 INVx1_ASAP7_75t_SL \i52/i297  (.A(\i52/n116 ),
    .Y(\i52/n115 ));
 NAND2xp5_ASAP7_75t_SL \i52/i298  (.A(\i52/n49 ),
    .B(\i52/n467 ),
    .Y(\i52/n140 ));
 NAND2xp5_ASAP7_75t_SL \i52/i299  (.A(\i52/n441 ),
    .B(\i52/n57 ),
    .Y(\i52/n114 ));
 INVx2_ASAP7_75t_SL \i52/i3  (.A(\i52/n498 ),
    .Y(\i52/n3 ));
 NOR3xp33_ASAP7_75t_SL \i52/i30  (.A(\i52/n327 ),
    .B(\i52/n343 ),
    .C(\i52/n375 ),
    .Y(\i52/n389 ));
 NAND2xp5_ASAP7_75t_SL \i52/i300  (.A(\i52/n58 ),
    .B(\i52/n56 ),
    .Y(\i52/n113 ));
 NAND2xp5_ASAP7_75t_SL \i52/i301  (.A(\i52/n38 ),
    .B(\i52/n59 ),
    .Y(\i52/n112 ));
 NAND2xp33_ASAP7_75t_SL \i52/i302  (.A(\i52/n480 ),
    .B(\i52/n45 ),
    .Y(\i52/n111 ));
 NAND2xp5_ASAP7_75t_SL \i52/i303  (.A(\i52/n3 ),
    .B(\i52/n47 ),
    .Y(\i52/n110 ));
 NAND2xp5_ASAP7_75t_SL \i52/i304  (.A(\i52/n49 ),
    .B(\i52/n3 ),
    .Y(\i52/n109 ));
 NAND2xp5_ASAP7_75t_SL \i52/i305  (.A(\i52/n52 ),
    .B(\i52/n51 ),
    .Y(\i52/n108 ));
 NAND2xp5_ASAP7_75t_SL \i52/i306  (.A(\i52/n35 ),
    .B(\i52/n43 ),
    .Y(\i52/n107 ));
 NAND2xp5_ASAP7_75t_SL \i52/i307  (.A(\i52/n35 ),
    .B(\i52/n444 ),
    .Y(\i52/n139 ));
 AND2x2_ASAP7_75t_SL \i52/i308  (.A(\i52/n43 ),
    .B(\i52/n53 ),
    .Y(\i52/n138 ));
 NAND2xp5_ASAP7_75t_SL \i52/i309  (.A(\i52/n52 ),
    .B(\i52/n5 ),
    .Y(\i52/n21 ));
 NOR2x1_ASAP7_75t_SL \i52/i31  (.A(\i52/n372 ),
    .B(\i52/n332 ),
    .Y(\i52/n388 ));
 NAND2xp5_ASAP7_75t_SL \i52/i310  (.A(\i52/n62 ),
    .B(\i52/n41 ),
    .Y(\i52/n133 ));
 AND2x2_ASAP7_75t_SL \i52/i311  (.A(\i52/n49 ),
    .B(\i52/n454 ),
    .Y(\i52/n131 ));
 NOR2xp67_ASAP7_75t_SL \i52/i312  (.A(\i52/n448 ),
    .B(\i52/n556 ),
    .Y(\i52/n20 ));
 NAND2xp5_ASAP7_75t_SL \i52/i313  (.A(\i52/n48 ),
    .B(\i52/n3 ),
    .Y(\i52/n106 ));
 NAND2xp5_ASAP7_75t_SL \i52/i314  (.A(\i52/n54 ),
    .B(\i52/n48 ),
    .Y(\i52/n129 ));
 NAND2xp5_ASAP7_75t_SL \i52/i315  (.A(\i52/n454 ),
    .B(\i52/n47 ),
    .Y(\i52/n105 ));
 NOR2xp33_ASAP7_75t_SL \i52/i316  (.A(\i52/n415 ),
    .B(\i52/n15 ),
    .Y(\i52/n104 ));
 NAND2xp5_ASAP7_75t_SL \i52/i317  (.A(\i52/n48 ),
    .B(\i52/n41 ),
    .Y(\i52/n127 ));
 NOR2xp33_ASAP7_75t_SL \i52/i318  (.A(\i52/n446 ),
    .B(\i52/n427 ),
    .Y(\i52/n103 ));
 NOR2xp33_ASAP7_75t_L \i52/i319  (.A(\i52/n62 ),
    .B(\i52/n39 ),
    .Y(\i52/n125 ));
 NAND2xp5_ASAP7_75t_SL \i52/i32  (.A(\i52/n330 ),
    .B(\i52/n349 ),
    .Y(\i52/n387 ));
 NAND2xp5_ASAP7_75t_SL \i52/i320  (.A(\i52/n62 ),
    .B(\i52/n44 ),
    .Y(\i52/n123 ));
 NAND2xp5_ASAP7_75t_SL \i52/i321  (.A(\i52/n62 ),
    .B(\i52/n52 ),
    .Y(\i52/n120 ));
 NAND2xp5_ASAP7_75t_SL \i52/i322  (.A(\i52/n49 ),
    .B(\i52/n54 ),
    .Y(\i52/n102 ));
 NOR2xp67_ASAP7_75t_SL \i52/i323  (.A(\i52/n441 ),
    .B(\i52/n49 ),
    .Y(\i52/n118 ));
 NOR2xp33_ASAP7_75t_L \i52/i324  (.A(\i52/n496 ),
    .B(\i52/n58 ),
    .Y(\i52/n101 ));
 OR2x2_ASAP7_75t_SL \i52/i325  (.A(\i52/n39 ),
    .B(\i52/n48 ),
    .Y(\i52/n116 ));
 INVxp67_ASAP7_75t_SL \i52/i326  (.A(\i52/n518 ),
    .Y(\i52/n100 ));
 INVxp67_ASAP7_75t_SL \i52/i327  (.A(\i52/n97 ),
    .Y(\i52/n98 ));
 INVx1_ASAP7_75t_SL \i52/i328  (.A(\i52/n566 ),
    .Y(\i52/n96 ));
 INVxp67_ASAP7_75t_SL \i52/i329  (.A(\i52/n438 ),
    .Y(\i52/n93 ));
 NOR3x1_ASAP7_75t_SL \i52/i33  (.A(\i52/n25 ),
    .B(\i52/n345 ),
    .C(\i52/n272 ),
    .Y(\i52/n395 ));
 INVxp67_ASAP7_75t_SL \i52/i330  (.A(\i52/n91 ),
    .Y(\i52/n92 ));
 INVxp67_ASAP7_75t_SL \i52/i331  (.A(\i52/n476 ),
    .Y(\i52/n90 ));
 INVxp67_ASAP7_75t_SL \i52/i332  (.A(\i52/n88 ),
    .Y(\i52/n89 ));
 INVxp67_ASAP7_75t_R \i52/i333  (.A(\i52/n519 ),
    .Y(\i52/n87 ));
 INVxp33_ASAP7_75t_SL \i52/i334  (.A(\i52/n85 ),
    .Y(\i52/n86 ));
 INVxp67_ASAP7_75t_SL \i52/i335  (.A(\i52/n80 ),
    .Y(\i52/n81 ));
 INVx1_ASAP7_75t_SL \i52/i336  (.A(\i52/n77 ),
    .Y(\i52/n78 ));
 INVx1_ASAP7_75t_SL \i52/i337  (.A(\i52/n17 ),
    .Y(\i52/n18 ));
 NAND2xp5_ASAP7_75t_SL \i52/i338  (.A(\i52/n443 ),
    .B(\i52/n53 ),
    .Y(\i52/n76 ));
 NAND2xp5_ASAP7_75t_SL \i52/i339  (.A(\i52/n39 ),
    .B(\i52/n54 ),
    .Y(\i52/n75 ));
 NOR3xp33_ASAP7_75t_SL \i52/i34  (.A(\i52/n288 ),
    .B(\i52/n25 ),
    .C(\i52/n369 ),
    .Y(\i52/n385 ));
 NAND2xp5_ASAP7_75t_SL \i52/i340  (.A(\i52/n46 ),
    .B(\i52/n53 ),
    .Y(\i52/n19 ));
 NAND2xp5_ASAP7_75t_SL \i52/i341  (.A(\i52/n55 ),
    .B(\i52/n459 ),
    .Y(\i52/n74 ));
 NAND2xp5_ASAP7_75t_SL \i52/i342  (.A(\i52/n46 ),
    .B(\i52/n54 ),
    .Y(\i52/n73 ));
 NAND2xp5_ASAP7_75t_SL \i52/i343  (.A(\i52/n54 ),
    .B(\i52/n38 ),
    .Y(\i52/n72 ));
 NAND2xp5_ASAP7_75t_SL \i52/i344  (.A(\i52/n444 ),
    .B(\i52/n454 ),
    .Y(\i52/n71 ));
 NAND2xp5_ASAP7_75t_SL \i52/i345  (.A(\i52/n51 ),
    .B(\i52/n44 ),
    .Y(\i52/n70 ));
 NAND2xp5_ASAP7_75t_L \i52/i346  (.A(\i52/n16 ),
    .B(\i52/n36 ),
    .Y(\i52/n69 ));
 NOR2xp33_ASAP7_75t_SL \i52/i347  (.A(\i52/n496 ),
    .B(\i52/n45 ),
    .Y(\i52/n68 ));
 AND2x2_ASAP7_75t_SL \i52/i348  (.A(\i52/n5 ),
    .B(\i52/n54 ),
    .Y(\i52/n99 ));
 NAND2xp5_ASAP7_75t_SL \i52/i349  (.A(\i52/n441 ),
    .B(\i52/n454 ),
    .Y(\i52/n97 ));
 NOR2xp33_ASAP7_75t_SL \i52/i35  (.A(\i52/n350 ),
    .B(\i52/n25 ),
    .Y(\i52/n384 ));
 NAND2xp5_ASAP7_75t_SL \i52/i350  (.A(\i52/n444 ),
    .B(\i52/n44 ),
    .Y(\i52/n95 ));
 NAND2xp5_ASAP7_75t_SL \i52/i351  (.A(\i52/n38 ),
    .B(\i52/n53 ),
    .Y(\i52/n67 ));
 AND2x2_ASAP7_75t_SL \i52/i352  (.A(\i52/n5 ),
    .B(\i52/n41 ),
    .Y(\i52/n94 ));
 NAND2xp5_ASAP7_75t_SL \i52/i353  (.A(\i52/n443 ),
    .B(\i52/n41 ),
    .Y(\i52/n91 ));
 NAND2xp5_ASAP7_75t_SL \i52/i354  (.A(\i52/n38 ),
    .B(\i52/n41 ),
    .Y(\i52/n88 ));
 NAND2xp33_ASAP7_75t_L \i52/i355  (.A(\i52/n40 ),
    .B(\i52/n550 ),
    .Y(\i52/n66 ));
 NOR2xp67_ASAP7_75t_L \i52/i356  (.A(\i52/n36 ),
    .B(\i52/n45 ),
    .Y(\i52/n85 ));
 NAND2xp5_ASAP7_75t_SL \i52/i357  (.A(\i52/n39 ),
    .B(\i52/n57 ),
    .Y(\i52/n84 ));
 NAND2xp5_ASAP7_75t_SL \i52/i358  (.A(\i52/n15 ),
    .B(\i52/n16 ),
    .Y(\i52/n83 ));
 NOR2x1_ASAP7_75t_L \i52/i359  (.A(\i52/n534 ),
    .B(\i52/n53 ),
    .Y(\i52/n82 ));
 NOR3xp33_ASAP7_75t_SL \i52/i36  (.A(\i52/n328 ),
    .B(\i52/n323 ),
    .C(\i52/n8 ),
    .Y(\i52/n383 ));
 NAND2xp5_ASAP7_75t_SL \i52/i360  (.A(\i52/n5 ),
    .B(\i52/n57 ),
    .Y(\i52/n65 ));
 NAND2xp5_ASAP7_75t_SL \i52/i361  (.A(\i52/n46 ),
    .B(\i52/n44 ),
    .Y(\i52/n80 ));
 NAND2xp5_ASAP7_75t_SL \i52/i362  (.A(\i52/n444 ),
    .B(\i52/n57 ),
    .Y(\i52/n79 ));
 NOR2xp33_ASAP7_75t_SL \i52/i363  (.A(\i52/n515 ),
    .B(\i52/n15 ),
    .Y(\i52/n64 ));
 NOR2xp33_ASAP7_75t_SL \i52/i364  (.A(\i52/n515 ),
    .B(\i52/n496 ),
    .Y(\i52/n63 ));
 NAND2xp5_ASAP7_75t_SL \i52/i365  (.A(\i52/n46 ),
    .B(\i52/n467 ),
    .Y(\i52/n77 ));
 NAND2xp5_ASAP7_75t_SL \i52/i366  (.A(\i52/n5 ),
    .B(\i52/n44 ),
    .Y(\i52/n17 ));
 INVx1_ASAP7_75t_SL \i52/i367  (.A(\i52/n62 ),
    .Y(\i52/n61 ));
 INVx3_ASAP7_75t_SL \i52/i368  (.A(\i52/n60 ),
    .Y(\i52/n59 ));
 INVx3_ASAP7_75t_SL \i52/i369  (.A(\i52/n441 ),
    .Y(\i52/n58 ));
 NAND4xp25_ASAP7_75t_SL \i52/i37  (.A(\i52/n310 ),
    .B(\i52/n304 ),
    .C(\i52/n303 ),
    .D(\i52/n337 ),
    .Y(\i52/n382 ));
 INVx2_ASAP7_75t_SL \i52/i370  (.A(\i52/n443 ),
    .Y(\i52/n56 ));
 INVx2_ASAP7_75t_SL \i52/i371  (.A(\i52/n444 ),
    .Y(\i52/n55 ));
 INVx3_ASAP7_75t_SL \i52/i372  (.A(\i52/n50 ),
    .Y(\i52/n49 ));
 AND2x4_ASAP7_75t_SL \i52/i373  (.A(\i52/n33 ),
    .B(\i52/n507 ),
    .Y(\i52/n62 ));
 OR2x4_ASAP7_75t_SL \i52/i374  (.A(\i52/n29 ),
    .B(\i52/n6 ),
    .Y(\i52/n60 ));
 AND2x4_ASAP7_75t_SL \i52/i375  (.A(\i52/n551 ),
    .B(\i52/n30 ),
    .Y(\i52/n57 ));
 NAND2x1_ASAP7_75t_SL \i52/i376  (.A(\i52/n551 ),
    .B(\i52/n30 ),
    .Y(\i52/n16 ));
 AND2x4_ASAP7_75t_SL \i52/i377  (.A(\i52/n551 ),
    .B(\i52/n485 ),
    .Y(\i52/n54 ));
 AND2x4_ASAP7_75t_SL \i52/i378  (.A(\i52/n451 ),
    .B(\i52/n14 ),
    .Y(\i52/n53 ));
 AND2x4_ASAP7_75t_SL \i52/i379  (.A(\i52/n451 ),
    .B(\i52/n551 ),
    .Y(\i52/n52 ));
 NAND3xp33_ASAP7_75t_L \i52/i38  (.A(\i52/n286 ),
    .B(\i52/n304 ),
    .C(\i52/n354 ),
    .Y(\i52/n381 ));
 AND2x4_ASAP7_75t_SL \i52/i380  (.A(\i52/n33 ),
    .B(\i52/n477 ),
    .Y(\i52/n51 ));
 OR2x6_ASAP7_75t_SL \i52/i381  (.A(\i52/n34 ),
    .B(\i52/n440 ),
    .Y(\i52/n50 ));
 INVx4_ASAP7_75t_SL \i52/i382  (.A(\i52/n46 ),
    .Y(\i52/n45 ));
 INVx3_ASAP7_75t_SL \i52/i383  (.A(\i52/n44 ),
    .Y(\i52/n15 ));
 INVx4_ASAP7_75t_SL \i52/i384  (.A(\i52/n43 ),
    .Y(\i52/n42 ));
 INVx3_ASAP7_75t_SL \i52/i385  (.A(\i52/n38 ),
    .Y(\i52/n37 ));
 INVx3_ASAP7_75t_SL \i52/i386  (.A(\i52/n36 ),
    .Y(\i52/n35 ));
 AND2x4_ASAP7_75t_SL \i52/i387  (.A(\i52/n33 ),
    .B(\i52/n10 ),
    .Y(\i52/n48 ));
 AND2x4_ASAP7_75t_SL \i52/i388  (.A(\i52/n32 ),
    .B(\i52/n507 ),
    .Y(\i52/n47 ));
 AND2x4_ASAP7_75t_SL \i52/i389  (.A(\i52/n32 ),
    .B(\i52/n10 ),
    .Y(\i52/n46 ));
 NAND3xp33_ASAP7_75t_SL \i52/i39  (.A(\i52/n290 ),
    .B(\i52/n338 ),
    .C(\i52/n324 ),
    .Y(\i52/n380 ));
 AND2x4_ASAP7_75t_SL \i52/i390  (.A(\i52/n552 ),
    .B(\i52/n14 ),
    .Y(\i52/n44 ));
 AND2x4_ASAP7_75t_SL \i52/i391  (.A(\i52/n4 ),
    .B(\i52/n10 ),
    .Y(\i52/n43 ));
 AND2x4_ASAP7_75t_SL \i52/i392  (.A(\i52/n2 ),
    .B(\i52/n30 ),
    .Y(\i52/n41 ));
 NAND2x1_ASAP7_75t_SL \i52/i393  (.A(\i52/n2 ),
    .B(\i52/n30 ),
    .Y(\i52/n40 ));
 AND2x4_ASAP7_75t_SL \i52/i394  (.A(\i52/n32 ),
    .B(\i52/n477 ),
    .Y(\i52/n39 ));
 AND2x4_ASAP7_75t_SL \i52/i395  (.A(\i52/n411 ),
    .B(\i52/n477 ),
    .Y(\i52/n38 ));
 OR2x6_ASAP7_75t_SL \i52/i396  (.A(\i52/n28 ),
    .B(\i52/n31 ),
    .Y(\i52/n36 ));
 NAND2xp5_ASAP7_75t_SL \i52/i397  (.A(\i52/n11 ),
    .B(\i52/n0 ),
    .Y(\i52/n31 ));
 NAND2x1p5_ASAP7_75t_SL \i52/i398  (.A(n17[4]),
    .B(n17[5]),
    .Y(\i52/n34 ));
 AND2x2_ASAP7_75t_SL \i52/i399  (.A(\i52/n26 ),
    .B(\i52/n9 ),
    .Y(\i52/n33 ));
 INVx2_ASAP7_75t_SL \i52/i4  (.A(\i52/n34 ),
    .Y(\i52/n4 ));
 NAND2xp5_ASAP7_75t_L \i52/i40  (.A(\i52/n574 ),
    .B(\i52/n370 ),
    .Y(\i52/n379 ));
 AND2x2_ASAP7_75t_SL \i52/i400  (.A(n17[4]),
    .B(\i52/n26 ),
    .Y(\i52/n32 ));
 INVx2_ASAP7_75t_SL \i52/i401  (.A(\i52/n6 ),
    .Y(\i52/n30 ));
 NAND2xp5_ASAP7_75t_SL \i52/i402  (.A(\i52/n27 ),
    .B(\i52/n1 ),
    .Y(\i52/n28 ));
 NAND2x1_ASAP7_75t_SL \i52/i403  (.A(n17[3]),
    .B(\i52/n0 ),
    .Y(\i52/n29 ));
 INVx1_ASAP7_75t_SL \i52/i404  (.A(n17[1]),
    .Y(\i52/n27 ));
 INVx3_ASAP7_75t_SL \i52/i405  (.A(n17[5]),
    .Y(\i52/n26 ));
 INVx2_ASAP7_75t_SL \i52/i406  (.A(n17[6]),
    .Y(\i52/n13 ));
 INVx2_ASAP7_75t_SL \i52/i407  (.A(n17[7]),
    .Y(\i52/n12 ));
 INVx2_ASAP7_75t_SL \i52/i408  (.A(n17[3]),
    .Y(\i52/n11 ));
 INVx1_ASAP7_75t_SL \i52/i409  (.A(\i52/n338 ),
    .Y(\i52/n8 ));
 NAND2xp33_ASAP7_75t_SL \i52/i41  (.A(\i52/n335 ),
    .B(\i52/n352 ),
    .Y(\i52/n378 ));
 AND2x2_ASAP7_75t_L \i52/i410  (.A(\i52/n12 ),
    .B(n17[6]),
    .Y(\i52/n10 ));
 INVx2_ASAP7_75t_SL \i52/i411  (.A(n17[4]),
    .Y(\i52/n9 ));
 OR2x2_ASAP7_75t_SL \i52/i412  (.A(\i52/n94 ),
    .B(\i52/n537 ),
    .Y(\i52/n7 ));
 OR2x2_ASAP7_75t_SL \i52/i413  (.A(n17[0]),
    .B(n17[1]),
    .Y(\i52/n6 ));
 NAND2xp5_ASAP7_75t_SL \i52/i414  (.A(\i52/n5 ),
    .B(\i52/n409 ),
    .Y(\i52/n407 ));
 NAND2xp5_ASAP7_75t_SL \i52/i415  (.A(\i52/n39 ),
    .B(\i52/n409 ),
    .Y(\i52/n408 ));
 NAND2xp5_ASAP7_75t_SL \i52/i416  (.A(\i52/n46 ),
    .B(\i52/n409 ),
    .Y(\i52/n410 ));
 INVx2_ASAP7_75t_SL \i52/i417  (.A(\i52/n567 ),
    .Y(\i52/n411 ));
 AND2x4_ASAP7_75t_SL \i52/i418  (.A(\i52/n507 ),
    .B(\i52/n411 ),
    .Y(\i52/n412 ));
 AOI22xp5_ASAP7_75t_SL \i52/i419  (.A1(\i52/n412 ),
    .A2(\i52/n409 ),
    .B1(\i52/n38 ),
    .B2(\i52/n57 ),
    .Y(\i52/n413 ));
 NOR2x1_ASAP7_75t_SL \i52/i42  (.A(\i52/n351 ),
    .B(\i52/n360 ),
    .Y(\i52/n386 ));
 NAND2xp5_ASAP7_75t_SL \i52/i420  (.A(\i52/n412 ),
    .B(\i52/n467 ),
    .Y(\i52/n414 ));
 INVx3_ASAP7_75t_SL \i52/i421  (.A(\i52/n412 ),
    .Y(\i52/n415 ));
 AND2x2_ASAP7_75t_SL \i52/i422  (.A(\i52/n412 ),
    .B(\i52/n3 ),
    .Y(\i52/n416 ));
 AOI22xp5_ASAP7_75t_SL \i52/i423  (.A1(\i52/n39 ),
    .A2(\i52/n41 ),
    .B1(\i52/n454 ),
    .B2(\i52/n412 ),
    .Y(\i52/n417 ));
 AOI222xp33_ASAP7_75t_SL \i52/i424  (.A1(\i52/n54 ),
    .A2(\i52/n412 ),
    .B1(\i52/n5 ),
    .B2(\i52/n35 ),
    .C1(\i52/n52 ),
    .C2(\i52/n47 ),
    .Y(\i52/n418 ));
 NAND2xp5_ASAP7_75t_SL \i52/i425  (.A(\i52/n412 ),
    .B(\i52/n52 ),
    .Y(\i52/n419 ));
 AOI22xp5_ASAP7_75t_SL \i52/i426  (.A1(\i52/n454 ),
    .A2(\i52/n111 ),
    .B1(\i52/n412 ),
    .B2(\i52/n44 ),
    .Y(\i52/n420 ));
 AOI221xp5_ASAP7_75t_SL \i52/i427  (.A1(\i52/n412 ),
    .A2(\i52/n35 ),
    .B1(\i52/n41 ),
    .B2(\i52/n49 ),
    .C(\i52/n528 ),
    .Y(\i52/n421 ));
 OAI21xp5_ASAP7_75t_SL \i52/i428  (.A1(\i52/n53 ),
    .A2(\i52/n57 ),
    .B(\i52/n412 ),
    .Y(\i52/n422 ));
 AOI221xp5_ASAP7_75t_SL \i52/i429  (.A1(\i52/n54 ),
    .A2(\i52/n62 ),
    .B1(\i52/n534 ),
    .B2(\i52/n412 ),
    .C(\i52/n142 ),
    .Y(\i52/n423 ));
 NAND2xp33_ASAP7_75t_L \i52/i43  (.A(\i52/n340 ),
    .B(\i52/n312 ),
    .Y(\i52/n375 ));
 NAND2xp5_ASAP7_75t_SL \i52/i430  (.A(\i52/n424 ),
    .B(\i52/n412 ),
    .Y(\i52/n425 ));
 AND2x4_ASAP7_75t_SL \i52/i431  (.A(\i52/n2 ),
    .B(\i52/n451 ),
    .Y(\i52/n424 ));
 NOR2xp67_ASAP7_75t_L \i52/i432  (.A(\i52/n424 ),
    .B(\i52/n409 ),
    .Y(\i52/n426 ));
 INVx4_ASAP7_75t_SL \i52/i433  (.A(\i52/n424 ),
    .Y(\i52/n427 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i52/i434  (.A1(\i52/n424 ),
    .A2(\i52/n41 ),
    .B(\i52/n51 ),
    .C(\i52/n99 ),
    .Y(\i52/n428 ));
 O2A1O1Ixp33_ASAP7_75t_R \i52/i435  (.A1(\i52/n441 ),
    .A2(\i52/n5 ),
    .B(\i52/n424 ),
    .C(\i52/n18 ),
    .Y(\i52/n429 ));
 AOI21xp5_ASAP7_75t_SL \i52/i436  (.A1(\i52/n116 ),
    .A2(\i52/n424 ),
    .B(\i52/n168 ),
    .Y(\i52/n430 ));
 AOI22xp5_ASAP7_75t_SL \i52/i437  (.A1(\i52/n467 ),
    .A2(\i52/n113 ),
    .B1(\i52/n47 ),
    .B2(\i52/n424 ),
    .Y(\i52/n431 ));
 OA21x2_ASAP7_75t_SL \i52/i438  (.A1(\i52/n5 ),
    .A2(\i52/n62 ),
    .B(\i52/n424 ),
    .Y(\i52/n432 ));
 OAI21xp33_ASAP7_75t_SL \i52/i439  (.A1(\i52/n424 ),
    .A2(\i52/n53 ),
    .B(\i52/n39 ),
    .Y(\i52/n433 ));
 NAND2xp33_ASAP7_75t_L \i52/i44  (.A(\i52/n574 ),
    .B(\i52/n318 ),
    .Y(\i52/n374 ));
 AOI22xp5_ASAP7_75t_SL \i52/i440  (.A1(\i52/n39 ),
    .A2(\i52/n454 ),
    .B1(\i52/n38 ),
    .B2(\i52/n424 ),
    .Y(\i52/n434 ));
 NAND2xp5_ASAP7_75t_SL \i52/i441  (.A(\i52/n441 ),
    .B(\i52/n424 ),
    .Y(\i52/n435 ));
 NAND2xp5_ASAP7_75t_SL \i52/i442  (.A(\i52/n49 ),
    .B(\i52/n424 ),
    .Y(\i52/n436 ));
 NAND2xp5_ASAP7_75t_SL \i52/i443  (.A(\i52/n444 ),
    .B(\i52/n424 ),
    .Y(\i52/n437 ));
 NAND2xp5_ASAP7_75t_SL \i52/i444  (.A(\i52/n443 ),
    .B(\i52/n424 ),
    .Y(\i52/n438 ));
 INVx2_ASAP7_75t_SL \i52/i445  (.A(\i52/n439 ),
    .Y(\i52/n440 ));
 AND2x2_ASAP7_75t_SL \i52/i446  (.A(n17[7]),
    .B(n17[6]),
    .Y(\i52/n439 ));
 AND2x4_ASAP7_75t_SL \i52/i447  (.A(\i52/n439 ),
    .B(\i52/n411 ),
    .Y(\i52/n441 ));
 AOI211xp5_ASAP7_75t_SL \i52/i448  (.A1(\i52/n59 ),
    .A2(\i52/n439 ),
    .B(\i52/n520 ),
    .C(\i52/n89 ),
    .Y(\i52/n442 ));
 AND2x4_ASAP7_75t_SL \i52/i449  (.A(\i52/n439 ),
    .B(\i52/n33 ),
    .Y(\i52/n443 ));
 NOR2xp67_ASAP7_75t_SL \i52/i45  (.A(\i52/n317 ),
    .B(\i52/n342 ),
    .Y(\i52/n373 ));
 AND2x4_ASAP7_75t_SL \i52/i450  (.A(\i52/n439 ),
    .B(\i52/n32 ),
    .Y(\i52/n444 ));
 INVx3_ASAP7_75t_SL \i52/i451  (.A(\i52/n54 ),
    .Y(\i52/n445 ));
 INVx3_ASAP7_75t_SL \i52/i452  (.A(\i52/n47 ),
    .Y(\i52/n446 ));
 INVx2_ASAP7_75t_SL \i52/i453  (.A(\i52/n52 ),
    .Y(\i52/n447 ));
 INVx3_ASAP7_75t_SL \i52/i454  (.A(\i52/n48 ),
    .Y(\i52/n448 ));
 OAI22xp5_ASAP7_75t_SL \i52/i455  (.A1(\i52/n445 ),
    .A2(\i52/n446 ),
    .B1(\i52/n447 ),
    .B2(\i52/n448 ),
    .Y(\i52/n449 ));
 AOI22xp33_ASAP7_75t_SL \i52/i456  (.A1(\i52/n62 ),
    .A2(\i52/n534 ),
    .B1(\i52/n48 ),
    .B2(\i52/n3 ),
    .Y(\i52/n450 ));
 AND2x2_ASAP7_75t_SL \i52/i457  (.A(n17[0]),
    .B(n17[1]),
    .Y(\i52/n451 ));
 AND2x2_ASAP7_75t_SL \i52/i458  (.A(\i52/n11 ),
    .B(\i52/n0 ),
    .Y(\i52/n452 ));
 INVx4_ASAP7_75t_SL \i52/i459  (.A(\i52/n453 ),
    .Y(\i52/n454 ));
 NAND3xp33_ASAP7_75t_SL \i52/i46  (.A(\i52/n307 ),
    .B(\i52/n315 ),
    .C(\i52/n558 ),
    .Y(\i52/n372 ));
 NAND2x1p5_ASAP7_75t_SL \i52/i460  (.A(\i52/n451 ),
    .B(\i52/n452 ),
    .Y(\i52/n453 ));
 OAI22xp5_ASAP7_75t_SL \i52/i461  (.A1(\i52/n42 ),
    .A2(\i52/n453 ),
    .B1(\i52/n50 ),
    .B2(\i52/n550 ),
    .Y(\i52/n455 ));
 OAI221xp5_ASAP7_75t_SL \i52/i462  (.A1(\i52/n484 ),
    .A2(\i52/n60 ),
    .B1(\i52/n453 ),
    .B2(\i52/n459 ),
    .C(\i52/n425 ),
    .Y(\i52/n456 ));
 NAND2xp33_ASAP7_75t_R \i52/i463  (.A(\i52/n453 ),
    .B(\i52/n498 ),
    .Y(\i52/n457 ));
 NOR2xp33_ASAP7_75t_SL \i52/i464  (.A(\i52/n453 ),
    .B(\i52/n37 ),
    .Y(\i52/n458 ));
 INVx2_ASAP7_75t_SL \i52/i465  (.A(\i52/n51 ),
    .Y(\i52/n459 ));
 INVx2_ASAP7_75t_SL \i52/i466  (.A(\i52/n39 ),
    .Y(\i52/n460 ));
 NOR2xp33_ASAP7_75t_SL \i52/i467  (.A(\i52/n176 ),
    .B(\i52/n539 ),
    .Y(\i52/n461 ));
 NOR4xp25_ASAP7_75t_SL \i52/i468  (.A(\i52/n539 ),
    .B(\i52/n128 ),
    .C(\i52/n544 ),
    .D(\i52/n131 ),
    .Y(\i52/n462 ));
 OA21x2_ASAP7_75t_SL \i52/i469  (.A1(\i52/n42 ),
    .A2(\i52/n525 ),
    .B(\i52/n19 ),
    .Y(\i52/n463 ));
 NOR2x1_ASAP7_75t_SL \i52/i47  (.A(\i52/n265 ),
    .B(\i52/n326 ),
    .Y(\i52/n371 ));
 INVx5_ASAP7_75t_SL \i52/i470  (.A(\i52/n466 ),
    .Y(\i52/n467 ));
 OR2x6_ASAP7_75t_SL \i52/i471  (.A(\i52/n464 ),
    .B(\i52/n465 ),
    .Y(\i52/n466 ));
 INVx1_ASAP7_75t_SL \i52/i472  (.A(\i52/n485 ),
    .Y(\i52/n464 ));
 INVx2_ASAP7_75t_SL \i52/i473  (.A(\i52/n452 ),
    .Y(\i52/n465 ));
 A2O1A1Ixp33_ASAP7_75t_R \i52/i474  (.A1(\i52/n466 ),
    .A2(\i52/n40 ),
    .B(\i52/n459 ),
    .C(\i52/n84 ),
    .Y(\i52/n468 ));
 AOI21xp5_ASAP7_75t_L \i52/i475  (.A1(\i52/n480 ),
    .A2(\i52/n125 ),
    .B(\i52/n466 ),
    .Y(\i52/n469 ));
 OAI222xp33_ASAP7_75t_SL \i52/i476  (.A1(\i52/n466 ),
    .A2(\i52/n37 ),
    .B1(\i52/n40 ),
    .B2(\i52/n415 ),
    .C1(\i52/n447 ),
    .C2(\i52/n50 ),
    .Y(\i52/n470 ));
 OAI221xp5_ASAP7_75t_SL \i52/i477  (.A1(\i52/n466 ),
    .A2(\i52/n55 ),
    .B1(\i52/n556 ),
    .B2(\i52/n459 ),
    .C(\i52/n154 ),
    .Y(\i52/n471 ));
 OAI221xp5_ASAP7_75t_SL \i52/i478  (.A1(\i52/n466 ),
    .A2(\i52/n56 ),
    .B1(\i52/n16 ),
    .B2(\i52/n415 ),
    .C(\i52/n179 ),
    .Y(\i52/n472 ));
 OAI22x1_ASAP7_75t_L \i52/i479  (.A1(\i52/n446 ),
    .A2(\i52/n466 ),
    .B1(\i52/n515 ),
    .B2(\i52/n15 ),
    .Y(\i52/n473 ));
 NOR2xp33_ASAP7_75t_SL \i52/i48  (.A(\i52/n333 ),
    .B(\i52/n248 ),
    .Y(\i52/n370 ));
 OAI22xp33_ASAP7_75t_SL \i52/i480  (.A1(\i52/n446 ),
    .A2(\i52/n36 ),
    .B1(\i52/n466 ),
    .B2(\i52/n480 ),
    .Y(\i52/n474 ));
 OAI22xp5_ASAP7_75t_SL \i52/i481  (.A1(\i52/n61 ),
    .A2(\i52/n498 ),
    .B1(\i52/n569 ),
    .B2(\i52/n466 ),
    .Y(\i52/n475 ));
 NOR2xp67_ASAP7_75t_SL \i52/i482  (.A(\i52/n42 ),
    .B(\i52/n466 ),
    .Y(\i52/n476 ));
 AND2x4_ASAP7_75t_SL \i52/i483  (.A(n17[7]),
    .B(\i52/n13 ),
    .Y(\i52/n477 ));
 AND2x4_ASAP7_75t_SL \i52/i484  (.A(\i52/n4 ),
    .B(\i52/n477 ),
    .Y(\i52/n478 ));
 NAND2xp5_ASAP7_75t_SL \i52/i485  (.A(\i52/n478 ),
    .B(\i52/n409 ),
    .Y(\i52/n479 ));
 INVx3_ASAP7_75t_SL \i52/i486  (.A(\i52/n478 ),
    .Y(\i52/n480 ));
 OAI31xp33_ASAP7_75t_SL \i52/i487  (.A1(\i52/n454 ),
    .A2(\i52/n534 ),
    .A3(\i52/n59 ),
    .B(\i52/n478 ),
    .Y(\i52/n481 ));
 AOI21xp5_ASAP7_75t_SL \i52/i488  (.A1(\i52/n53 ),
    .A2(\i52/n478 ),
    .B(\i52/n187 ),
    .Y(\i52/n482 ));
 NOR2xp33_ASAP7_75t_SL \i52/i489  (.A(\i52/n478 ),
    .B(\i52/n441 ),
    .Y(\i52/n483 ));
 NAND2xp67_ASAP7_75t_SL \i52/i49  (.A(\i52/n340 ),
    .B(\i52/n336 ),
    .Y(\i52/n369 ));
 NOR2x1_ASAP7_75t_SL \i52/i490  (.A(\i52/n478 ),
    .B(\i52/n443 ),
    .Y(\i52/n484 ));
 AND2x4_ASAP7_75t_SL \i52/i491  (.A(n17[0]),
    .B(\i52/n27 ),
    .Y(\i52/n485 ));
 INVx2_ASAP7_75t_SL \i52/i492  (.A(\i52/n29 ),
    .Y(\i52/n14 ));
 NAND2xp5_ASAP7_75t_SL \i52/i493  (.A(\i52/n478 ),
    .B(\i52/n486 ),
    .Y(\i52/n487 ));
 AND2x4_ASAP7_75t_SL \i52/i494  (.A(\i52/n485 ),
    .B(\i52/n14 ),
    .Y(\i52/n486 ));
 NAND2xp5_ASAP7_75t_SL \i52/i495  (.A(\i52/n486 ),
    .B(\i52/n412 ),
    .Y(\i52/n488 ));
 NAND2xp5_ASAP7_75t_SL \i52/i496  (.A(\i52/n43 ),
    .B(\i52/n486 ),
    .Y(\i52/n489 ));
 NAND2xp5_ASAP7_75t_SL \i52/i497  (.A(\i52/n443 ),
    .B(\i52/n486 ),
    .Y(\i52/n490 ));
 NAND2xp5_ASAP7_75t_SL \i52/i498  (.A(\i52/n5 ),
    .B(\i52/n486 ),
    .Y(\i52/n491 ));
 NAND2xp5_ASAP7_75t_SL \i52/i499  (.A(\i52/n486 ),
    .B(\i52/n47 ),
    .Y(\i52/n492 ));
 INVx2_ASAP7_75t_SL \i52/i5  (.A(\i52/n569 ),
    .Y(\i52/n5 ));
 NOR2x1_ASAP7_75t_SL \i52/i50  (.A(\i52/n541 ),
    .B(\i52/n342 ),
    .Y(\i52/n368 ));
 AOI22xp5_ASAP7_75t_SL \i52/i500  (.A1(\i52/n47 ),
    .A2(\i52/n454 ),
    .B1(\i52/n444 ),
    .B2(\i52/n486 ),
    .Y(\i52/n493 ));
 AOI22xp5_ASAP7_75t_SL \i52/i501  (.A1(\i52/n441 ),
    .A2(\i52/n486 ),
    .B1(\i52/n444 ),
    .B2(\i52/n52 ),
    .Y(\i52/n494 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i52/i502  (.A1(\i52/n454 ),
    .A2(\i52/n486 ),
    .B(\i52/n5 ),
    .C(\i52/n126 ),
    .Y(\i52/n495 ));
 INVx3_ASAP7_75t_SL \i52/i503  (.A(\i52/n486 ),
    .Y(\i52/n496 ));
 OAI21xp5_ASAP7_75t_SL \i52/i504  (.A1(\i52/n486 ),
    .A2(\i52/n409 ),
    .B(\i52/n444 ),
    .Y(\i52/n497 ));
 NAND2x1p5_ASAP7_75t_SL \i52/i505  (.A(\i52/n2 ),
    .B(\i52/n485 ),
    .Y(\i52/n498 ));
 NAND2xp5_ASAP7_75t_SL \i52/i506  (.A(\i52/n38 ),
    .B(\i52/n3 ),
    .Y(\i52/n499 ));
 NAND2xp33_ASAP7_75t_L \i52/i507  (.A(\i52/n3 ),
    .B(\i52/n444 ),
    .Y(\i52/n500 ));
 NAND2xp5_ASAP7_75t_SL \i52/i508  (.A(\i52/n3 ),
    .B(\i52/n46 ),
    .Y(\i52/n501 ));
 NAND2xp5_ASAP7_75t_SL \i52/i509  (.A(\i52/n441 ),
    .B(\i52/n3 ),
    .Y(\i52/n502 ));
 NOR2x1_ASAP7_75t_SL \i52/i51  (.A(\i52/n316 ),
    .B(\i52/n327 ),
    .Y(\i52/n367 ));
 AOI22xp5_ASAP7_75t_SL \i52/i510  (.A1(\i52/n443 ),
    .A2(\i52/n454 ),
    .B1(\i52/n39 ),
    .B2(\i52/n3 ),
    .Y(\i52/n503 ));
 OAI31xp33_ASAP7_75t_SL \i52/i511  (.A1(\i52/n52 ),
    .A2(\i52/n3 ),
    .A3(\i52/n44 ),
    .B(\i52/n39 ),
    .Y(\i52/n504 ));
 NOR2xp33_ASAP7_75t_SL \i52/i512  (.A(\i52/n424 ),
    .B(\i52/n3 ),
    .Y(\i52/n505 ));
 AO21x2_ASAP7_75t_SL \i52/i513  (.A1(\i52/n443 ),
    .A2(\i52/n3 ),
    .B(\i52/n449 ),
    .Y(\i52/n506 ));
 AND2x2_ASAP7_75t_SL \i52/i514  (.A(\i52/n12 ),
    .B(\i52/n13 ),
    .Y(\i52/n507 ));
 AOI22xp5_ASAP7_75t_SL \i52/i515  (.A1(\i52/n508 ),
    .A2(\i52/n409 ),
    .B1(\i52/n444 ),
    .B2(\i52/n3 ),
    .Y(\i52/n509 ));
 AND2x4_ASAP7_75t_SL \i52/i516  (.A(\i52/n507 ),
    .B(\i52/n4 ),
    .Y(\i52/n508 ));
 NAND2xp5_ASAP7_75t_SL \i52/i517  (.A(\i52/n508 ),
    .B(\i52/n3 ),
    .Y(\i52/n510 ));
 AOI22xp33_ASAP7_75t_SL \i52/i518  (.A1(\i52/n48 ),
    .A2(\i52/n454 ),
    .B1(\i52/n508 ),
    .B2(\i52/n486 ),
    .Y(\i52/n511 ));
 AOI22xp5_ASAP7_75t_SL \i52/i519  (.A1(\i52/n508 ),
    .A2(\i52/n41 ),
    .B1(\i52/n478 ),
    .B2(\i52/n52 ),
    .Y(\i52/n512 ));
 NAND2xp5_ASAP7_75t_SL \i52/i52  (.A(\i52/n281 ),
    .B(\i52/n321 ),
    .Y(\i52/n366 ));
 AOI22xp5_ASAP7_75t_SL \i52/i520  (.A1(\i52/n508 ),
    .A2(\i52/n424 ),
    .B1(\i52/n443 ),
    .B2(\i52/n52 ),
    .Y(\i52/n513 ));
 AND2x2_ASAP7_75t_SL \i52/i521  (.A(\i52/n508 ),
    .B(\i52/n52 ),
    .Y(\i52/n514 ));
 INVx2_ASAP7_75t_SL \i52/i522  (.A(\i52/n508 ),
    .Y(\i52/n515 ));
 AOI22xp5_ASAP7_75t_SL \i52/i523  (.A1(\i52/n508 ),
    .A2(\i52/n467 ),
    .B1(\i52/n441 ),
    .B2(\i52/n44 ),
    .Y(\i52/n516 ));
 AOI22xp5_ASAP7_75t_SL \i52/i524  (.A1(\i52/n35 ),
    .A2(\i52/n38 ),
    .B1(\i52/n508 ),
    .B2(\i52/n53 ),
    .Y(\i52/n517 ));
 NAND2xp5_ASAP7_75t_SL \i52/i525  (.A(\i52/n508 ),
    .B(\i52/n534 ),
    .Y(\i52/n518 ));
 NAND2xp5_ASAP7_75t_SL \i52/i526  (.A(\i52/n35 ),
    .B(\i52/n508 ),
    .Y(\i52/n519 ));
 AND2x2_ASAP7_75t_SL \i52/i527  (.A(\i52/n508 ),
    .B(\i52/n57 ),
    .Y(\i52/n520 ));
 AND2x2_ASAP7_75t_SL \i52/i528  (.A(\i52/n508 ),
    .B(\i52/n454 ),
    .Y(\i52/n521 ));
 NAND2xp5_ASAP7_75t_SL \i52/i529  (.A(\i52/n508 ),
    .B(\i52/n54 ),
    .Y(\i52/n522 ));
 NOR5xp2_ASAP7_75t_SL \i52/i53  (.A(\i52/n215 ),
    .B(\i52/n533 ),
    .C(\i52/n226 ),
    .D(\i52/n24 ),
    .E(\i52/n471 ),
    .Y(\i52/n365 ));
 OR2x2_ASAP7_75t_SL \i52/i530  (.A(\i52/n0 ),
    .B(n17[3]),
    .Y(\i52/n523 ));
 NAND2xp5_ASAP7_75t_SL \i52/i531  (.A(n17[1]),
    .B(\i52/n1 ),
    .Y(\i52/n524 ));
 NOR2xp33_ASAP7_75t_SL \i52/i532  (.A(\i52/n525 ),
    .B(\i52/n460 ),
    .Y(\i52/n526 ));
 OR2x4_ASAP7_75t_SL \i52/i533  (.A(\i52/n523 ),
    .B(\i52/n524 ),
    .Y(\i52/n525 ));
 NOR2xp67_ASAP7_75t_L \i52/i534  (.A(\i52/n525 ),
    .B(\i52/n448 ),
    .Y(\i52/n527 ));
 OAI22xp5_ASAP7_75t_SL \i52/i535  (.A1(\i52/n42 ),
    .A2(\i52/n40 ),
    .B1(\i52/n525 ),
    .B2(\i52/n460 ),
    .Y(\i52/n528 ));
 OAI21xp5_ASAP7_75t_SL \i52/i536  (.A1(\i52/n55 ),
    .A2(\i52/n525 ),
    .B(\i52/n489 ),
    .Y(\i52/n529 ));
 OAI22xp33_ASAP7_75t_SL \i52/i537  (.A1(\i52/n460 ),
    .A2(\i52/n60 ),
    .B1(\i52/n525 ),
    .B2(\i52/n446 ),
    .Y(\i52/n530 ));
 AOI31xp33_ASAP7_75t_SL \i52/i538  (.A1(\i52/n42 ),
    .A2(\i52/n56 ),
    .A3(\i52/n459 ),
    .B(\i52/n525 ),
    .Y(\i52/n531 ));
 AO21x1_ASAP7_75t_SL \i52/i539  (.A1(\i52/n525 ),
    .A2(\i52/n114 ),
    .B(\i52/n483 ),
    .Y(\i52/n532 ));
 NOR2x1_ASAP7_75t_SL \i52/i54  (.A(\i52/n8 ),
    .B(\i52/n328 ),
    .Y(\i52/n364 ));
 OAI221xp5_ASAP7_75t_SL \i52/i540  (.A1(\i52/n496 ),
    .A2(\i52/n448 ),
    .B1(\i52/n42 ),
    .B2(\i52/n525 ),
    .C(\i52/n19 ),
    .Y(\i52/n533 ));
 INVx4_ASAP7_75t_SL \i52/i541  (.A(\i52/n525 ),
    .Y(\i52/n534 ));
 OAI221xp5_ASAP7_75t_SL \i52/i542  (.A1(\i52/n45 ),
    .A2(\i52/n40 ),
    .B1(\i52/n525 ),
    .B2(\i52/n37 ),
    .C(\i52/n519 ),
    .Y(\i52/n535 ));
 AND2x4_ASAP7_75t_SL \i52/i543  (.A(\i52/n452 ),
    .B(\i52/n552 ),
    .Y(\i52/n409 ));
 OAI22xp5_ASAP7_75t_SL \i52/i544  (.A1(\i52/n42 ),
    .A2(\i52/n536 ),
    .B1(\i52/n50 ),
    .B2(\i52/n525 ),
    .Y(\i52/n537 ));
 INVx4_ASAP7_75t_SL \i52/i545  (.A(\i52/n409 ),
    .Y(\i52/n536 ));
 OAI22x1_ASAP7_75t_SL \i52/i546  (.A1(\i52/n448 ),
    .A2(\i52/n536 ),
    .B1(\i52/n459 ),
    .B2(\i52/n466 ),
    .Y(\i52/n538 ));
 OAI22xp5_ASAP7_75t_SL \i52/i547  (.A1(\i52/n459 ),
    .A2(\i52/n536 ),
    .B1(\i52/n556 ),
    .B2(\i52/n460 ),
    .Y(\i52/n539 ));
 OAI22xp5_ASAP7_75t_SL \i52/i548  (.A1(\i52/n536 ),
    .A2(\i52/n118 ),
    .B1(\i52/n50 ),
    .B2(\i52/n554 ),
    .Y(\i52/n540 ));
 OAI211xp5_ASAP7_75t_SL \i52/i549  (.A1(\i52/n61 ),
    .A2(\i52/n536 ),
    .B(\i52/n136 ),
    .C(\i52/n95 ),
    .Y(\i52/n541 ));
 NAND2x1_ASAP7_75t_SL \i52/i55  (.A(\i52/n325 ),
    .B(\i52/n305 ),
    .Y(\i52/n377 ));
 OAI222xp33_ASAP7_75t_SL \i52/i550  (.A1(\i52/n536 ),
    .A2(\i52/n56 ),
    .B1(\i52/n60 ),
    .B2(\i52/n55 ),
    .C1(\i52/n16 ),
    .C2(\i52/n480 ),
    .Y(\i52/n542 ));
 OAI22xp5_ASAP7_75t_SL \i52/i551  (.A1(\i52/n61 ),
    .A2(\i52/n496 ),
    .B1(\i52/n45 ),
    .B2(\i52/n536 ),
    .Y(\i52/n543 ));
 AOI21xp33_ASAP7_75t_SL \i52/i552  (.A1(\i52/n556 ),
    .A2(\i52/n536 ),
    .B(\i52/n56 ),
    .Y(\i52/n544 ));
 OAI22xp33_ASAP7_75t_SL \i52/i553  (.A1(\i52/n16 ),
    .A2(\i52/n446 ),
    .B1(\i52/n536 ),
    .B2(\i52/n58 ),
    .Y(\i52/n545 ));
 OAI22xp33_ASAP7_75t_SL \i52/i554  (.A1(\i52/n56 ),
    .A2(\i52/n36 ),
    .B1(\i52/n536 ),
    .B2(\i52/n37 ),
    .Y(\i52/n546 ));
 OAI22xp5_ASAP7_75t_SL \i52/i555  (.A1(\i52/n480 ),
    .A2(\i52/n40 ),
    .B1(\i52/n50 ),
    .B2(\i52/n536 ),
    .Y(\i52/n547 ));
 NOR2xp33_ASAP7_75t_SL \i52/i556  (.A(\i52/n459 ),
    .B(\i52/n536 ),
    .Y(\i52/n548 ));
 NOR2xp33_ASAP7_75t_SL \i52/i557  (.A(\i52/n446 ),
    .B(\i52/n536 ),
    .Y(\i52/n549 ));
 INVx1_ASAP7_75t_SL \i52/i558  (.A(\i52/n53 ),
    .Y(\i52/n550 ));
 AND2x4_ASAP7_75t_SL \i52/i559  (.A(n17[3]),
    .B(n17[2]),
    .Y(\i52/n551 ));
 NOR2x1_ASAP7_75t_SL \i52/i56  (.A(\i52/n343 ),
    .B(\i52/n327 ),
    .Y(\i52/n363 ));
 INVx2_ASAP7_75t_SL \i52/i560  (.A(\i52/n524 ),
    .Y(\i52/n552 ));
 NOR2xp33_ASAP7_75t_SL \i52/i561  (.A(\i52/n553 ),
    .B(\i52/n486 ),
    .Y(\i52/n554 ));
 AND2x4_ASAP7_75t_SL \i52/i562  (.A(\i52/n551 ),
    .B(\i52/n552 ),
    .Y(\i52/n553 ));
 NAND2xp5_ASAP7_75t_SL \i52/i563  (.A(\i52/n478 ),
    .B(\i52/n553 ),
    .Y(\i52/n555 ));
 INVx3_ASAP7_75t_SL \i52/i564  (.A(\i52/n553 ),
    .Y(\i52/n556 ));
 OAI21xp5_ASAP7_75t_SL \i52/i565  (.A1(\i52/n553 ),
    .A2(\i52/n486 ),
    .B(\i52/n39 ),
    .Y(\i52/n557 ));
 AOI211xp5_ASAP7_75t_SL \i52/i566  (.A1(\i52/n553 ),
    .A2(\i52/n49 ),
    .B(\i52/n416 ),
    .C(\i52/n506 ),
    .Y(\i52/n558 ));
 OAI21xp5_ASAP7_75t_SL \i52/i567  (.A1(\i52/n53 ),
    .A2(\i52/n553 ),
    .B(\i52/n62 ),
    .Y(\i52/n559 ));
 OAI21xp5_ASAP7_75t_SL \i52/i568  (.A1(\i52/n553 ),
    .A2(\i52/n454 ),
    .B(\i52/n444 ),
    .Y(\i52/n560 ));
 OAI21xp5_ASAP7_75t_SL \i52/i569  (.A1(\i52/n46 ),
    .A2(\i52/n51 ),
    .B(\i52/n553 ),
    .Y(\i52/n561 ));
 NOR2x1_ASAP7_75t_SL \i52/i57  (.A(\i52/n264 ),
    .B(\i52/n326 ),
    .Y(\i52/n376 ));
 NAND2xp5_ASAP7_75t_SL \i52/i570  (.A(\i52/n47 ),
    .B(\i52/n553 ),
    .Y(\i52/n562 ));
 NAND2xp5_ASAP7_75t_SL \i52/i571  (.A(\i52/n43 ),
    .B(\i52/n553 ),
    .Y(\i52/n563 ));
 AND2x2_ASAP7_75t_SL \i52/i572  (.A(\i52/n441 ),
    .B(\i52/n553 ),
    .Y(\i52/n564 ));
 NAND2xp5_ASAP7_75t_SL \i52/i573  (.A(\i52/n38 ),
    .B(\i52/n553 ),
    .Y(\i52/n565 ));
 NOR2xp33_ASAP7_75t_SL \i52/i574  (.A(\i52/n553 ),
    .B(\i52/n57 ),
    .Y(\i52/n566 ));
 NAND2xp5_ASAP7_75t_SL \i52/i575  (.A(\i52/n9 ),
    .B(n17[5]),
    .Y(\i52/n567 ));
 OAI221xp5_ASAP7_75t_SL \i52/i576  (.A1(\i52/n82 ),
    .A2(\i52/n61 ),
    .B1(\i52/n82 ),
    .B2(\i52/n569 ),
    .C(\i52/n219 ),
    .Y(\i52/n570 ));
 OR2x2_ASAP7_75t_SL \i52/i577  (.A(\i52/n568 ),
    .B(\i52/n567 ),
    .Y(\i52/n569 ));
 NAND2xp5_ASAP7_75t_SL \i52/i578  (.A(\i52/n12 ),
    .B(n17[6]),
    .Y(\i52/n568 ));
 NAND2xp5_ASAP7_75t_SL \i52/i579  (.A(\i52/n50 ),
    .B(\i52/n569 ),
    .Y(\i52/n571 ));
 INVxp67_ASAP7_75t_SL \i52/i58  (.A(\i52/n361 ),
    .Y(\i52/n362 ));
 OAI21xp5_ASAP7_75t_SL \i52/i580  (.A1(\i52/n569 ),
    .A2(\i52/n498 ),
    .B(\i52/n88 ),
    .Y(\i52/n572 ));
 AND4x1_ASAP7_75t_SL \i52/i581  (.A(\i52/n418 ),
    .B(\i52/n250 ),
    .C(\i52/n581 ),
    .D(\i52/n196 ),
    .Y(\i52/n573 ));
 AND4x1_ASAP7_75t_SL \i52/i582  (.A(\i52/n208 ),
    .B(\i52/n482 ),
    .C(\i52/n431 ),
    .D(\i52/n418 ),
    .Y(\i52/n574 ));
 AND2x2_ASAP7_75t_SL \i52/i583  (.A(\i52/n575 ),
    .B(\i52/n339 ),
    .Y(\i52/n576 ));
 AOI21xp33_ASAP7_75t_SL \i52/i584  (.A1(\i52/n35 ),
    .A2(\i52/n51 ),
    .B(\i52/n520 ),
    .Y(\i52/n575 ));
 NAND3xp33_ASAP7_75t_SL \i52/i585  (.A(\i52/n577 ),
    .B(\i52/n191 ),
    .C(\i52/n242 ),
    .Y(\i52/n578 ));
 AO21x1_ASAP7_75t_SL \i52/i586  (.A1(\i52/n448 ),
    .A2(\i52/n42 ),
    .B(\i52/n427 ),
    .Y(\i52/n577 ));
 NOR3xp33_ASAP7_75t_SL \i52/i587  (.A(\i52/n579 ),
    .B(\i52/n240 ),
    .C(\i52/n449 ),
    .Y(\i52/n580 ));
 OAI21xp5_ASAP7_75t_SL \i52/i588  (.A1(\i52/n50 ),
    .A2(\i52/n16 ),
    .B(\i52/n501 ),
    .Y(\i52/n579 ));
 AOI21xp5_ASAP7_75t_SL \i52/i589  (.A1(\i52/n43 ),
    .A2(\i52/n52 ),
    .B(\i52/n528 ),
    .Y(\i52/n581 ));
 INVxp67_ASAP7_75t_SL \i52/i59  (.A(\i52/n357 ),
    .Y(\i52/n358 ));
 NOR2x2_ASAP7_75t_SL \i52/i6  (.A(\i52/n402 ),
    .B(\i52/n401 ),
    .Y(n16[4]));
 AND5x1_ASAP7_75t_SL \i52/i60  (.A(\i52/n277 ),
    .B(\i52/n581 ),
    .C(\i52/n270 ),
    .D(\i52/n495 ),
    .E(\i52/n186 ),
    .Y(\i52/n356 ));
 NOR3xp33_ASAP7_75t_SL \i52/i61  (.A(\i52/n287 ),
    .B(\i52/n269 ),
    .C(\i52/n252 ),
    .Y(\i52/n355 ));
 NOR3xp33_ASAP7_75t_SL \i52/i62  (.A(\i52/n313 ),
    .B(\i52/n253 ),
    .C(\i52/n214 ),
    .Y(\i52/n354 ));
 AND5x1_ASAP7_75t_SL \i52/i63  (.A(\i52/n244 ),
    .B(\i52/n256 ),
    .C(\i52/n442 ),
    .D(\i52/n247 ),
    .E(\i52/n192 ),
    .Y(\i52/n353 ));
 NOR2xp33_ASAP7_75t_SL \i52/i64  (.A(\i52/n314 ),
    .B(\i52/n319 ),
    .Y(\i52/n352 ));
 NAND4xp25_ASAP7_75t_SL \i52/i65  (.A(\i52/n296 ),
    .B(\i52/n304 ),
    .C(\i52/n309 ),
    .D(\i52/n292 ),
    .Y(\i52/n351 ));
 NAND5xp2_ASAP7_75t_SL \i52/i66  (.A(\i52/n276 ),
    .B(\i52/n237 ),
    .C(\i52/n164 ),
    .D(\i52/n153 ),
    .E(\i52/n223 ),
    .Y(\i52/n350 ));
 NOR4xp25_ASAP7_75t_SL \i52/i67  (.A(\i52/n267 ),
    .B(\i52/n533 ),
    .C(\i52/n227 ),
    .D(\i52/n209 ),
    .Y(\i52/n349 ));
 NAND4xp25_ASAP7_75t_SL \i52/i68  (.A(\i52/n284 ),
    .B(\i52/n298 ),
    .C(\i52/n301 ),
    .D(\i52/n303 ),
    .Y(\i52/n348 ));
 NAND4xp25_ASAP7_75t_SL \i52/i69  (.A(\i52/n311 ),
    .B(\i52/n309 ),
    .C(\i52/n463 ),
    .D(\i52/n185 ),
    .Y(\i52/n347 ));
 NOR2x2_ASAP7_75t_SL \i52/i7  (.A(\i52/n397 ),
    .B(\i52/n403 ),
    .Y(n16[3]));
 NAND3xp33_ASAP7_75t_SL \i52/i70  (.A(\i52/n303 ),
    .B(\i52/n275 ),
    .C(\i52/n408 ),
    .Y(\i52/n361 ));
 NAND4xp75_ASAP7_75t_SL \i52/i71  (.A(\i52/n219 ),
    .B(\i52/n199 ),
    .C(\i52/n263 ),
    .D(\i52/n21 ),
    .Y(\i52/n360 ));
 NAND2xp33_ASAP7_75t_L \i52/i72  (.A(\i52/n283 ),
    .B(\i52/n344 ),
    .Y(\i52/n346 ));
 AND2x2_ASAP7_75t_SL \i52/i73  (.A(\i52/n286 ),
    .B(\i52/n334 ),
    .Y(\i52/n359 ));
 NAND2x1p5_ASAP7_75t_SL \i52/i74  (.A(\i52/n341 ),
    .B(\i52/n297 ),
    .Y(\i52/n357 ));
 INVxp67_ASAP7_75t_SL \i52/i75  (.A(\i52/n344 ),
    .Y(\i52/n345 ));
 NOR5xp2_ASAP7_75t_SL \i52/i76  (.A(\i52/n469 ),
    .B(\i52/n213 ),
    .C(\i52/n158 ),
    .D(\i52/n514 ),
    .E(\i52/n526 ),
    .Y(\i52/n337 ));
 NOR3xp33_ASAP7_75t_SL \i52/i77  (.A(\i52/n308 ),
    .B(\i52/n230 ),
    .C(\i52/n542 ),
    .Y(\i52/n336 ));
 NOR2xp33_ASAP7_75t_SL \i52/i78  (.A(\i52/n266 ),
    .B(\i52/n285 ),
    .Y(\i52/n335 ));
 NOR2xp33_ASAP7_75t_SL \i52/i79  (.A(\i52/n306 ),
    .B(\i52/n257 ),
    .Y(\i52/n334 ));
 AND5x2_ASAP7_75t_SL \i52/i8  (.A(\i52/n395 ),
    .B(\i52/n386 ),
    .C(\i52/n388 ),
    .D(\i52/n373 ),
    .E(\i52/n365 ),
    .Y(n16[6]));
 NOR2x1_ASAP7_75t_SL \i52/i80  (.A(\i52/n271 ),
    .B(\i52/n245 ),
    .Y(\i52/n344 ));
 NAND3xp33_ASAP7_75t_SL \i52/i81  (.A(\i52/n222 ),
    .B(\i52/n504 ),
    .C(\i52/n513 ),
    .Y(\i52/n333 ));
 NAND2xp5_ASAP7_75t_L \i52/i82  (.A(\i52/n305 ),
    .B(\i52/n462 ),
    .Y(\i52/n332 ));
 NAND2xp67_ASAP7_75t_SL \i52/i83  (.A(\i52/n461 ),
    .B(\i52/n295 ),
    .Y(\i52/n331 ));
 NAND3xp33_ASAP7_75t_SL \i52/i84  (.A(\i52/n581 ),
    .B(\i52/n210 ),
    .C(\i52/n196 ),
    .Y(\i52/n343 ));
 NOR3xp33_ASAP7_75t_SL \i52/i85  (.A(\i52/n570 ),
    .B(\i52/n7 ),
    .C(\i52/n472 ),
    .Y(\i52/n330 ));
 NAND2xp5_ASAP7_75t_SL \i52/i86  (.A(\i52/n479 ),
    .B(\i52/n284 ),
    .Y(\i52/n342 ));
 OR3x1_ASAP7_75t_SL \i52/i87  (.A(\i52/n215 ),
    .B(\i52/n226 ),
    .C(\i52/n24 ),
    .Y(\i52/n329 ));
 NOR2x1_ASAP7_75t_SL \i52/i88  (.A(\i52/n542 ),
    .B(\i52/n308 ),
    .Y(\i52/n341 ));
 NOR2xp33_ASAP7_75t_SL \i52/i89  (.A(\i52/n268 ),
    .B(\i52/n255 ),
    .Y(\i52/n340 ));
 AND3x4_ASAP7_75t_SL \i52/i9  (.A(\i52/n395 ),
    .B(\i52/n404 ),
    .C(\i52/n383 ),
    .Y(n16[1]));
 NOR2xp33_ASAP7_75t_SL \i52/i90  (.A(\i52/n456 ),
    .B(\i52/n294 ),
    .Y(\i52/n339 ));
 NOR3x1_ASAP7_75t_SL \i52/i91  (.A(\i52/n221 ),
    .B(\i52/n145 ),
    .C(\i52/n260 ),
    .Y(\i52/n338 ));
 NOR3xp33_ASAP7_75t_SL \i52/i92  (.A(\i52/n228 ),
    .B(\i52/n163 ),
    .C(\i52/n218 ),
    .Y(\i52/n325 ));
 NOR2xp33_ASAP7_75t_SL \i52/i93  (.A(\i52/n578 ),
    .B(\i52/n280 ),
    .Y(\i52/n324 ));
 NAND3xp33_ASAP7_75t_SL \i52/i94  (.A(\i52/n418 ),
    .B(\i52/n273 ),
    .C(\i52/n431 ),
    .Y(\i52/n323 ));
 NAND4xp25_ASAP7_75t_SL \i52/i95  (.A(\i52/n203 ),
    .B(\i52/n428 ),
    .C(\i52/n234 ),
    .D(\i52/n481 ),
    .Y(\i52/n322 ));
 NAND2x1_ASAP7_75t_SL \i52/i96  (.A(\i52/n293 ),
    .B(\i52/n307 ),
    .Y(\i52/n328 ));
 NOR5xp2_ASAP7_75t_SL \i52/i97  (.A(\i52/n302 ),
    .B(\i52/n468 ),
    .C(\i52/n93 ),
    .D(\i52/n172 ),
    .E(\i52/n122 ),
    .Y(\i52/n321 ));
 NAND3xp33_ASAP7_75t_SL \i52/i98  (.A(\i52/n259 ),
    .B(\i52/n278 ),
    .C(\i52/n516 ),
    .Y(\i52/n320 ));
 NAND2xp33_ASAP7_75t_SL \i52/i99  (.A(\i52/n430 ),
    .B(\i52/n299 ),
    .Y(\i52/n319 ));
 AOI22xp5_ASAP7_75t_SL i520 (.A1(n875),
    .A2(n1153),
    .B1(n876),
    .B2(n227),
    .Y(n952));
 OAI22xp5_ASAP7_75t_SL i521 (.A1(n1180),
    .A2(n800),
    .B1(n801),
    .B2(n543),
    .Y(n951));
 AOI22xp5_ASAP7_75t_SL i522 (.A1(n568),
    .A2(n500),
    .B1(n567),
    .B2(n499),
    .Y(n950));
 XNOR2xp5_ASAP7_75t_SL i523 (.A(n322),
    .B(n321),
    .Y(n949));
 XOR2xp5_ASAP7_75t_SL i524 (.A(n1210),
    .B(n323),
    .Y(n948));
 XOR2xp5_ASAP7_75t_SL i525 (.A(n603),
    .B(n1212),
    .Y(n947));
 AOI22xp5_ASAP7_75t_SL i526 (.A1(n513),
    .A2(n796),
    .B1(n797),
    .B2(n514),
    .Y(n946));
 XOR2xp5_ASAP7_75t_SL i527 (.A(n324),
    .B(n325),
    .Y(n945));
 XOR2xp5_ASAP7_75t_SL i528 (.A(n796),
    .B(n626),
    .Y(n944));
 XOR2xp5_ASAP7_75t_SL i529 (.A(n327),
    .B(n1179),
    .Y(n943));
 INVx2_ASAP7_75t_SL \i53/i0  (.A(n15[7]),
    .Y(\i53/n0 ));
 INVx2_ASAP7_75t_SL \i53/i1  (.A(n15[2]),
    .Y(\i53/n1 ));
 NOR2x2_ASAP7_75t_SL \i53/i10  (.A(\i53/n404 ),
    .B(\i53/n410 ),
    .Y(n14[3]));
 NAND2x1_ASAP7_75t_SL \i53/i100  (.A(\i53/n300 ),
    .B(\i53/n314 ),
    .Y(\i53/n334 ));
 NOR5xp2_ASAP7_75t_SL \i53/i101  (.A(\i53/n309 ),
    .B(\i53/n553 ),
    .C(\i53/n100 ),
    .D(\i53/n179 ),
    .E(\i53/n127 ),
    .Y(\i53/n327 ));
 NAND3xp33_ASAP7_75t_SL \i53/i102  (.A(\i53/n264 ),
    .B(\i53/n576 ),
    .C(\i53/n540 ),
    .Y(\i53/n326 ));
 NAND2xp33_ASAP7_75t_SL \i53/i103  (.A(\i53/n476 ),
    .B(\i53/n306 ),
    .Y(\i53/n325 ));
 NOR5xp2_ASAP7_75t_SL \i53/i104  (.A(\i53/n250 ),
    .B(\i53/n220 ),
    .C(\i53/n237 ),
    .D(\i53/n197 ),
    .E(\i53/n163 ),
    .Y(\i53/n324 ));
 NAND5xp2_ASAP7_75t_SL \i53/i105  (.A(\i53/n440 ),
    .B(\i53/n541 ),
    .C(\i53/n154 ),
    .D(\i53/n475 ),
    .E(\i53/n559 ),
    .Y(\i53/n323 ));
 NAND3xp33_ASAP7_75t_SL \i53/i106  (.A(\i53/n201 ),
    .B(\i53/n464 ),
    .C(\i53/n287 ),
    .Y(\i53/n322 ));
 NOR5xp2_ASAP7_75t_SL \i53/i107  (.A(\i53/n199 ),
    .B(\i53/n86 ),
    .C(\i53/n193 ),
    .D(\i53/n208 ),
    .E(\i53/n76 ),
    .Y(\i53/n321 ));
 NAND5xp2_ASAP7_75t_SL \i53/i108  (.A(\i53/n21 ),
    .B(\i53/n516 ),
    .C(\i53/n154 ),
    .D(\i53/n435 ),
    .E(\i53/n142 ),
    .Y(\i53/n320 ));
 NOR5xp2_ASAP7_75t_SL \i53/i109  (.A(\i53/n172 ),
    .B(\i53/n517 ),
    .C(\i53/n162 ),
    .D(\i53/n138 ),
    .E(\i53/n136 ),
    .Y(\i53/n319 ));
 AND5x2_ASAP7_75t_SL \i53/i11  (.A(\i53/n402 ),
    .B(\i53/n393 ),
    .C(\i53/n395 ),
    .D(\i53/n380 ),
    .E(\i53/n372 ),
    .Y(n14[6]));
 NOR2xp33_ASAP7_75t_SL \i53/i110  (.A(\i53/n279 ),
    .B(\i53/n313 ),
    .Y(\i53/n318 ));
 NOR2xp33_ASAP7_75t_SL \i53/i111  (.A(\i53/n268 ),
    .B(\i53/n297 ),
    .Y(\i53/n317 ));
 NAND3x1_ASAP7_75t_SL \i53/i112  (.A(\i53/n500 ),
    .B(\i53/n541 ),
    .C(\i53/n295 ),
    .Y(\i53/n333 ));
 NAND3x1_ASAP7_75t_SL \i53/i113  (.A(\i53/n259 ),
    .B(\i53/n239 ),
    .C(\i53/n215 ),
    .Y(\i53/n332 ));
 AOI21xp5_ASAP7_75t_L \i53/i114  (.A1(\i53/n56 ),
    .A2(\i53/n487 ),
    .B(\i53/n123 ),
    .Y(\i53/n309 ));
 NOR2xp33_ASAP7_75t_SL \i53/i115  (.A(\i53/n250 ),
    .B(\i53/n518 ),
    .Y(\i53/n308 ));
 NAND2xp5_ASAP7_75t_SL \i53/i116  (.A(\i53/n460 ),
    .B(\i53/n267 ),
    .Y(\i53/n307 ));
 NOR2xp33_ASAP7_75t_SL \i53/i117  (.A(\i53/n266 ),
    .B(\i53/n22 ),
    .Y(\i53/n306 ));
 NOR2xp33_ASAP7_75t_SL \i53/i118  (.A(\i53/n245 ),
    .B(\i53/n255 ),
    .Y(\i53/n305 ));
 NOR2xp67_ASAP7_75t_SL \i53/i119  (.A(\i53/n129 ),
    .B(\i53/n252 ),
    .Y(\i53/n304 ));
 AND3x4_ASAP7_75t_SL \i53/i12  (.A(\i53/n402 ),
    .B(\i53/n411 ),
    .C(\i53/n390 ),
    .Y(n14[1]));
 NOR2xp33_ASAP7_75t_SL \i53/i120  (.A(\i53/n18 ),
    .B(\i53/n250 ),
    .Y(\i53/n303 ));
 NOR4xp25_ASAP7_75t_SL \i53/i121  (.A(\i53/n227 ),
    .B(\i53/n18 ),
    .C(\i53/n546 ),
    .D(\i53/n524 ),
    .Y(\i53/n302 ));
 NAND2xp5_ASAP7_75t_SL \i53/i122  (.A(\i53/n499 ),
    .B(\i53/n538 ),
    .Y(\i53/n301 ));
 NOR4xp25_ASAP7_75t_SL \i53/i123  (.A(\i53/n84 ),
    .B(\i53/n183 ),
    .C(\i53/n164 ),
    .D(\i53/n174 ),
    .Y(\i53/n300 ));
 NOR3xp33_ASAP7_75t_SL \i53/i124  (.A(\i53/n188 ),
    .B(\i53/n155 ),
    .C(\i53/n187 ),
    .Y(\i53/n299 ));
 NAND2xp5_ASAP7_75t_SL \i53/i125  (.A(\i53/n210 ),
    .B(\i53/n495 ),
    .Y(\i53/n298 ));
 NAND2xp33_ASAP7_75t_SL \i53/i126  (.A(\i53/n417 ),
    .B(\i53/n19 ),
    .Y(\i53/n297 ));
 NOR2xp33_ASAP7_75t_SL \i53/i127  (.A(\i53/n518 ),
    .B(\i53/n219 ),
    .Y(\i53/n296 ));
 NOR2x1p5_ASAP7_75t_SL \i53/i128  (.A(\i53/n205 ),
    .B(\i53/n534 ),
    .Y(\i53/n295 ));
 NAND2xp33_ASAP7_75t_SL \i53/i129  (.A(\i53/n264 ),
    .B(\i53/n248 ),
    .Y(\i53/n294 ));
 NOR2x1p5_ASAP7_75t_SL \i53/i13  (.A(\i53/n412 ),
    .B(\i53/n403 ),
    .Y(n14[5]));
 NAND3xp33_ASAP7_75t_SL \i53/i130  (.A(\i53/n20 ),
    .B(\i53/n451 ),
    .C(\i53/n529 ),
    .Y(\i53/n293 ));
 NOR3xp33_ASAP7_75t_SL \i53/i131  (.A(\i53/n158 ),
    .B(\i53/n169 ),
    .C(\i53/n147 ),
    .Y(\i53/n316 ));
 NAND2xp5_ASAP7_75t_SL \i53/i132  (.A(\i53/n226 ),
    .B(\i53/n157 ),
    .Y(\i53/n315 ));
 NOR2x1_ASAP7_75t_SL \i53/i133  (.A(\i53/n204 ),
    .B(\i53/n222 ),
    .Y(\i53/n314 ));
 NAND2xp5_ASAP7_75t_SL \i53/i134  (.A(\i53/n154 ),
    .B(\i53/n228 ),
    .Y(\i53/n313 ));
 NOR2x1_ASAP7_75t_SL \i53/i135  (.A(\i53/n206 ),
    .B(\i53/n253 ),
    .Y(\i53/n312 ));
 NAND2xp5_ASAP7_75t_SL \i53/i136  (.A(\i53/n477 ),
    .B(\i53/n459 ),
    .Y(\i53/n292 ));
 NOR2x1_ASAP7_75t_SL \i53/i137  (.A(\i53/n546 ),
    .B(\i53/n518 ),
    .Y(\i53/n311 ));
 NOR3x1_ASAP7_75t_SL \i53/i138  (.A(\i53/n162 ),
    .B(\i53/n508 ),
    .C(\i53/n135 ),
    .Y(\i53/n310 ));
 INVx1_ASAP7_75t_SL \i53/i139  (.A(\i53/n289 ),
    .Y(\i53/n290 ));
 AND2x4_ASAP7_75t_SL \i53/i14  (.A(\i53/n413 ),
    .B(\i53/n396 ),
    .Y(n14[0]));
 INVx1_ASAP7_75t_SL \i53/i140  (.A(\i53/n23 ),
    .Y(\i53/n288 ));
 NOR4xp25_ASAP7_75t_SL \i53/i141  (.A(\i53/n547 ),
    .B(\i53/n176 ),
    .C(\i53/n167 ),
    .D(\i53/n145 ),
    .Y(\i53/n287 ));
 AOI211xp5_ASAP7_75t_SL \i53/i142  (.A1(\i53/n88 ),
    .A2(\i53/n45 ),
    .B(\i53/n236 ),
    .C(\i53/n186 ),
    .Y(\i53/n286 ));
 NAND2xp33_ASAP7_75t_L \i53/i143  (.A(\i53/n216 ),
    .B(\i53/n235 ),
    .Y(\i53/n285 ));
 NAND5xp2_ASAP7_75t_SL \i53/i144  (.A(\i53/n566 ),
    .B(\i53/n182 ),
    .C(\i53/n192 ),
    .D(\i53/n563 ),
    .E(\i53/n469 ),
    .Y(\i53/n284 ));
 NOR2xp33_ASAP7_75t_SL \i53/i145  (.A(\i53/n209 ),
    .B(\i53/n211 ),
    .Y(\i53/n283 ));
 AOI211xp5_ASAP7_75t_SL \i53/i146  (.A1(\i53/n57 ),
    .A2(\i53/n126 ),
    .B(\i53/n549 ),
    .C(\i53/n139 ),
    .Y(\i53/n282 ));
 OA21x2_ASAP7_75t_SL \i53/i147  (.A1(\i53/n454 ),
    .A2(\i53/n56 ),
    .B(\i53/n516 ),
    .Y(\i53/n281 ));
 NOR4xp25_ASAP7_75t_SL \i53/i148  (.A(\i53/n194 ),
    .B(\i53/n132 ),
    .C(\i53/n152 ),
    .D(\i53/n135 ),
    .Y(\i53/n280 ));
 NAND5xp2_ASAP7_75t_SL \i53/i149  (.A(\i53/n112 ),
    .B(\i53/n562 ),
    .C(\i53/n445 ),
    .D(\i53/n481 ),
    .E(\i53/n75 ),
    .Y(\i53/n279 ));
 NOR3xp33_ASAP7_75t_SL \i53/i15  (.A(\i53/n385 ),
    .B(\i53/n381 ),
    .C(\i53/n388 ),
    .Y(\i53/n413 ));
 NOR3xp33_ASAP7_75t_SL \i53/i150  (.A(\i53/n223 ),
    .B(\i53/n133 ),
    .C(\i53/n74 ),
    .Y(\i53/n278 ));
 NAND2xp5_ASAP7_75t_SL \i53/i151  (.A(\i53/n488 ),
    .B(\i53/n21 ),
    .Y(\i53/n277 ));
 NAND5xp2_ASAP7_75t_SL \i53/i152  (.A(\i53/n565 ),
    .B(\i53/n467 ),
    .C(\i53/n452 ),
    .D(\i53/n144 ),
    .E(\i53/n557 ),
    .Y(\i53/n276 ));
 NAND4xp25_ASAP7_75t_SL \i53/i153  (.A(\i53/n233 ),
    .B(\i53/n424 ),
    .C(\i53/n85 ),
    .D(\i53/n461 ),
    .Y(\i53/n275 ));
 NAND5xp2_ASAP7_75t_SL \i53/i154  (.A(\i53/n577 ),
    .B(\i53/n419 ),
    .C(\i53/n178 ),
    .D(\i53/n466 ),
    .E(\i53/n81 ),
    .Y(\i53/n274 ));
 NAND2xp5_ASAP7_75t_SL \i53/i155  (.A(\i53/n496 ),
    .B(\i53/n225 ),
    .Y(\i53/n273 ));
 NAND3xp33_ASAP7_75t_SL \i53/i156  (.A(\i53/n221 ),
    .B(\i53/n536 ),
    .C(\i53/n503 ),
    .Y(\i53/n272 ));
 NAND2xp5_ASAP7_75t_SL \i53/i157  (.A(\i53/n500 ),
    .B(\i53/n541 ),
    .Y(\i53/n271 ));
 NOR2xp33_ASAP7_75t_L \i53/i158  (.A(\i53/n243 ),
    .B(\i53/n255 ),
    .Y(\i53/n291 ));
 NAND2xp5_ASAP7_75t_SL \i53/i159  (.A(\i53/n540 ),
    .B(\i53/n264 ),
    .Y(\i53/n270 ));
 NOR2x2_ASAP7_75t_SL \i53/i16  (.A(\i53/n405 ),
    .B(\i53/n406 ),
    .Y(n14[2]));
 NOR2x1p5_ASAP7_75t_SL \i53/i160  (.A(\i53/n551 ),
    .B(\i53/n247 ),
    .Y(\i53/n289 ));
 NAND3x1_ASAP7_75t_SL \i53/i161  (.A(\i53/n196 ),
    .B(\i53/n106 ),
    .C(\i53/n441 ),
    .Y(\i53/n23 ));
 INVxp67_ASAP7_75t_SL \i53/i162  (.A(\i53/n268 ),
    .Y(\i53/n269 ));
 INVxp67_ASAP7_75t_SL \i53/i163  (.A(\i53/n10 ),
    .Y(\i53/n267 ));
 INVxp67_ASAP7_75t_SL \i53/i164  (.A(\i53/n262 ),
    .Y(\i53/n263 ));
 INVxp67_ASAP7_75t_SL \i53/i165  (.A(\i53/n260 ),
    .Y(\i53/n261 ));
 INVx1_ASAP7_75t_SL \i53/i166  (.A(\i53/n258 ),
    .Y(\i53/n259 ));
 INVxp67_ASAP7_75t_SL \i53/i167  (.A(\i53/n495 ),
    .Y(\i53/n257 ));
 INVxp67_ASAP7_75t_SL \i53/i168  (.A(\i53/n253 ),
    .Y(\i53/n254 ));
 INVxp67_ASAP7_75t_SL \i53/i169  (.A(\i53/n515 ),
    .Y(\i53/n251 ));
 NAND4xp75_ASAP7_75t_SL \i53/i17  (.A(\i53/n371 ),
    .B(\i53/n391 ),
    .C(\i53/n369 ),
    .D(\i53/n578 ),
    .Y(\i53/n412 ));
 INVx1_ASAP7_75t_SL \i53/i170  (.A(\i53/n248 ),
    .Y(\i53/n249 ));
 NAND2x1_ASAP7_75t_SL \i53/i171  (.A(\i53/n442 ),
    .B(\i53/n166 ),
    .Y(\i53/n247 ));
 NOR2xp33_ASAP7_75t_SL \i53/i172  (.A(\i53/n574 ),
    .B(\i53/n188 ),
    .Y(\i53/n246 ));
 NAND2xp33_ASAP7_75t_SL \i53/i173  (.A(\i53/n451 ),
    .B(\i53/n154 ),
    .Y(\i53/n245 ));
 OAI21xp5_ASAP7_75t_SL \i53/i174  (.A1(\i53/n44 ),
    .A2(\i53/n483 ),
    .B(\i53/n143 ),
    .Y(\i53/n244 ));
 NAND2xp5_ASAP7_75t_SL \i53/i175  (.A(\i53/n134 ),
    .B(\i53/n451 ),
    .Y(\i53/n243 ));
 AOI211xp5_ASAP7_75t_SL \i53/i176  (.A1(\i53/n67 ),
    .A2(\i53/n28 ),
    .B(\i53/n89 ),
    .C(\i53/n96 ),
    .Y(\i53/n242 ));
 AOI31xp33_ASAP7_75t_SL \i53/i177  (.A1(\i53/n44 ),
    .A2(\i53/n444 ),
    .A3(\i53/n50 ),
    .B(\i53/n37 ),
    .Y(\i53/n241 ));
 NOR3xp33_ASAP7_75t_SL \i53/i178  (.A(\i53/n155 ),
    .B(\i53/n105 ),
    .C(\i53/n94 ),
    .Y(\i53/n240 ));
 NOR3xp33_ASAP7_75t_SL \i53/i179  (.A(\i53/n87 ),
    .B(\i53/n101 ),
    .C(\i53/n574 ),
    .Y(\i53/n239 ));
 NOR3xp33_ASAP7_75t_SL \i53/i18  (.A(\i53/n389 ),
    .B(\i53/n354 ),
    .C(\i53/n399 ),
    .Y(\i53/n411 ));
 OAI31xp33_ASAP7_75t_SL \i53/i180  (.A1(\i53/n39 ),
    .A2(\i53/n41 ),
    .A3(\i53/n55 ),
    .B(\i53/n67 ),
    .Y(\i53/n238 ));
 AOI21xp5_ASAP7_75t_SL \i53/i181  (.A1(\i53/n123 ),
    .A2(\i53/n50 ),
    .B(\i53/n473 ),
    .Y(\i53/n268 ));
 OAI221xp5_ASAP7_75t_SL \i53/i182  (.A1(\i53/n14 ),
    .A2(\i53/n69 ),
    .B1(\i53/n40 ),
    .B2(\i53/n569 ),
    .C(\i53/n479 ),
    .Y(\i53/n237 ));
 AOI21xp33_ASAP7_75t_SL \i53/i183  (.A1(\i53/n130 ),
    .A2(\i53/n38 ),
    .B(\i53/n462 ),
    .Y(\i53/n236 ));
 NOR3xp33_ASAP7_75t_SL \i53/i184  (.A(\i53/n173 ),
    .B(\i53/n87 ),
    .C(\i53/n109 ),
    .Y(\i53/n235 ));
 NAND3xp33_ASAP7_75t_SL \i53/i185  (.A(\i53/n15 ),
    .B(\i53/n17 ),
    .C(\i53/n128 ),
    .Y(\i53/n234 ));
 OAI21xp5_ASAP7_75t_SL \i53/i186  (.A1(\i53/n49 ),
    .A2(\i53/n124 ),
    .B(\i53/n57 ),
    .Y(\i53/n233 ));
 NAND4xp25_ASAP7_75t_SL \i53/i187  (.A(\i53/n137 ),
    .B(\i53/n461 ),
    .C(\i53/n429 ),
    .D(\i53/n115 ),
    .Y(\i53/n232 ));
 NAND2xp33_ASAP7_75t_SL \i53/i188  (.A(\i53/n497 ),
    .B(\i53/n465 ),
    .Y(\i53/n231 ));
 OAI211xp5_ASAP7_75t_SL \i53/i189  (.A1(\i53/n53 ),
    .A2(\i53/n462 ),
    .B(\i53/n480 ),
    .C(\i53/n564 ),
    .Y(\i53/n266 ));
 NAND4xp75_ASAP7_75t_SL \i53/i19  (.A(\i53/n370 ),
    .B(\i53/n401 ),
    .C(\i53/n375 ),
    .D(\i53/n365 ),
    .Y(\i53/n410 ));
 NOR2x1_ASAP7_75t_SL \i53/i190  (.A(\i53/n122 ),
    .B(\i53/n523 ),
    .Y(\i53/n265 ));
 NOR2xp67_ASAP7_75t_SL \i53/i191  (.A(\i53/n519 ),
    .B(\i53/n193 ),
    .Y(\i53/n264 ));
 NAND2xp5_ASAP7_75t_SL \i53/i192  (.A(\i53/n567 ),
    .B(\i53/n472 ),
    .Y(\i53/n22 ));
 NOR2xp33_ASAP7_75t_SL \i53/i193  (.A(\i53/n181 ),
    .B(\i53/n194 ),
    .Y(\i53/n262 ));
 OAI211xp5_ASAP7_75t_SL \i53/i194  (.A1(\i53/n50 ),
    .A2(\i53/n462 ),
    .B(\i53/n143 ),
    .C(\i53/n428 ),
    .Y(\i53/n260 ));
 OR2x2_ASAP7_75t_SL \i53/i195  (.A(\i53/n548 ),
    .B(\i53/n522 ),
    .Y(\i53/n258 ));
 OAI211xp5_ASAP7_75t_SL \i53/i196  (.A1(\i53/n69 ),
    .A2(\i53/n60 ),
    .B(\i53/n141 ),
    .C(\i53/n539 ),
    .Y(\i53/n256 ));
 NAND2xp5_ASAP7_75t_SL \i53/i197  (.A(\i53/n559 ),
    .B(\i53/n418 ),
    .Y(\i53/n255 ));
 NAND2xp5_ASAP7_75t_SL \i53/i198  (.A(\i53/n20 ),
    .B(\i53/n439 ),
    .Y(\i53/n253 ));
 NAND2xp5_ASAP7_75t_SL \i53/i199  (.A(\i53/n498 ),
    .B(\i53/n533 ),
    .Y(\i53/n252 ));
 INVx2_ASAP7_75t_SL \i53/i2  (.A(n15[0]),
    .Y(\i53/n2 ));
 AND3x4_ASAP7_75t_SL \i53/i20  (.A(\i53/n392 ),
    .B(\i53/n407 ),
    .C(\i53/n397 ),
    .Y(n14[7]));
 NAND2xp5_ASAP7_75t_SL \i53/i200  (.A(\i53/n482 ),
    .B(\i53/n530 ),
    .Y(\i53/n250 ));
 NOR2x1_ASAP7_75t_SL \i53/i201  (.A(\i53/n180 ),
    .B(\i53/n163 ),
    .Y(\i53/n248 ));
 INVxp67_ASAP7_75t_SL \i53/i202  (.A(\i53/n227 ),
    .Y(\i53/n228 ));
 INVx1_ASAP7_75t_SL \i53/i203  (.A(\i53/n464 ),
    .Y(\i53/n224 ));
 INVx1_ASAP7_75t_SL \i53/i204  (.A(\i53/n221 ),
    .Y(\i53/n222 ));
 NAND4xp25_ASAP7_75t_SL \i53/i205  (.A(\i53/n450 ),
    .B(\i53/n102 ),
    .C(\i53/n90 ),
    .D(\i53/n528 ),
    .Y(\i53/n218 ));
 AOI31xp33_ASAP7_75t_SL \i53/i206  (.A1(\i53/n433 ),
    .A2(\i53/n56 ),
    .A3(\i53/n37 ),
    .B(\i53/n38 ),
    .Y(\i53/n217 ));
 NOR4xp25_ASAP7_75t_SL \i53/i207  (.A(\i53/n84 ),
    .B(\i53/n545 ),
    .C(\i53/n501 ),
    .D(\i53/n73 ),
    .Y(\i53/n216 ));
 AOI211xp5_ASAP7_75t_SL \i53/i208  (.A1(\i53/n103 ),
    .A2(\i53/n63 ),
    .B(\i53/n133 ),
    .C(\i53/n78 ),
    .Y(\i53/n215 ));
 NOR2x1_ASAP7_75t_SL \i53/i209  (.A(\i53/n520 ),
    .B(\i53/n189 ),
    .Y(\i53/n214 ));
 NAND4xp75_ASAP7_75t_SL \i53/i21  (.A(\i53/n580 ),
    .B(\i53/n374 ),
    .C(\i53/n383 ),
    .D(\i53/n400 ),
    .Y(\i53/n409 ));
 OAI31xp33_ASAP7_75t_SL \i53/i210  (.A1(\i53/n46 ),
    .A2(\i53/n514 ),
    .A3(\i53/n67 ),
    .B(\i53/n51 ),
    .Y(\i53/n213 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i53/i211  (.A1(\i53/n462 ),
    .A2(\i53/n42 ),
    .B(\i53/n65 ),
    .C(\i53/n427 ),
    .Y(\i53/n212 ));
 OAI22xp5_ASAP7_75t_SL \i53/i212  (.A1(\i53/n60 ),
    .A2(\i53/n125 ),
    .B1(\i53/n53 ),
    .B2(\i53/n558 ),
    .Y(\i53/n211 ));
 NOR2xp33_ASAP7_75t_SL \i53/i213  (.A(\i53/n160 ),
    .B(\i53/n148 ),
    .Y(\i53/n210 ));
 NAND2xp33_ASAP7_75t_L \i53/i214  (.A(\i53/n449 ),
    .B(\i53/n453 ),
    .Y(\i53/n209 ));
 NAND2xp33_ASAP7_75t_SL \i53/i215  (.A(\i53/n185 ),
    .B(\i53/n560 ),
    .Y(\i53/n208 ));
 OA21x2_ASAP7_75t_SL \i53/i216  (.A1(\i53/n38 ),
    .A2(\i53/n483 ),
    .B(\i53/n98 ),
    .Y(\i53/n207 ));
 NAND2xp5_ASAP7_75t_SL \i53/i217  (.A(\i53/n198 ),
    .B(\i53/n493 ),
    .Y(\i53/n206 ));
 NAND4xp25_ASAP7_75t_SL \i53/i218  (.A(\i53/n484 ),
    .B(\i53/n116 ),
    .C(\i53/n82 ),
    .D(\i53/n432 ),
    .Y(\i53/n205 ));
 OAI221xp5_ASAP7_75t_SL \i53/i219  (.A1(\i53/n68 ),
    .A2(\i53/n65 ),
    .B1(\i53/n425 ),
    .B2(\i53/n507 ),
    .C(\i53/n502 ),
    .Y(\i53/n230 ));
 NAND2x1_ASAP7_75t_SL \i53/i22  (.A(\i53/n362 ),
    .B(\i53/n393 ),
    .Y(\i53/n408 ));
 OAI222xp33_ASAP7_75t_SL \i53/i220  (.A1(\i53/n526 ),
    .A2(\i53/n44 ),
    .B1(\i53/n569 ),
    .B2(\i53/n53 ),
    .C1(\i53/n425 ),
    .C2(\i53/n58 ),
    .Y(\i53/n204 ));
 AND3x1_ASAP7_75t_SL \i53/i221  (.A(\i53/n97 ),
    .B(\i53/n102 ),
    .C(\i53/n492 ),
    .Y(\i53/n203 ));
 NAND2xp33_ASAP7_75t_SL \i53/i222  (.A(\i53/n151 ),
    .B(\i53/n177 ),
    .Y(\i53/n202 ));
 OAI222xp33_ASAP7_75t_SL \i53/i223  (.A1(\i53/n60 ),
    .A2(\i53/n62 ),
    .B1(\i53/n68 ),
    .B2(\i53/n58 ),
    .C1(\i53/n14 ),
    .C2(\i53/n50 ),
    .Y(\i53/n229 ));
 NAND3x1_ASAP7_75t_SL \i53/i224  (.A(\i53/n455 ),
    .B(\i53/n117 ),
    .C(\i53/n114 ),
    .Y(\i53/n227 ));
 AOI22xp5_ASAP7_75t_SL \i53/i225  (.A1(\i53/n509 ),
    .A2(\i53/n67 ),
    .B1(\i53/n55 ),
    .B2(\i53/n514 ),
    .Y(\i53/n226 ));
 AOI22xp5_ASAP7_75t_SL \i53/i226  (.A1(\i53/n70 ),
    .A2(\i53/n79 ),
    .B1(\i53/n39 ),
    .B2(\i53/n57 ),
    .Y(\i53/n225 ));
 OAI21xp5_ASAP7_75t_SL \i53/i227  (.A1(\i53/n37 ),
    .A2(\i53/n65 ),
    .B(\i53/n491 ),
    .Y(\i53/n223 ));
 NOR2x1_ASAP7_75t_SL \i53/i228  (.A(\i53/n99 ),
    .B(\i53/n150 ),
    .Y(\i53/n221 ));
 OAI221xp5_ASAP7_75t_SL \i53/i229  (.A1(\i53/n16 ),
    .A2(\i53/n68 ),
    .B1(\i53/n47 ),
    .B2(\i53/n54 ),
    .C(\i53/n471 ),
    .Y(\i53/n220 ));
 NOR2xp67_ASAP7_75t_SL \i53/i23  (.A(\i53/n355 ),
    .B(\i53/n394 ),
    .Y(\i53/n407 ));
 OAI211xp5_ASAP7_75t_SL \i53/i230  (.A1(\i53/n54 ),
    .A2(\i53/n527 ),
    .B(\i53/n85 ),
    .C(\i53/n531 ),
    .Y(\i53/n219 ));
 NOR2x1_ASAP7_75t_SL \i53/i231  (.A(\i53/n468 ),
    .B(\i53/n153 ),
    .Y(\i53/n21 ));
 NOR2xp33_ASAP7_75t_SL \i53/i232  (.A(\i53/n107 ),
    .B(\i53/n195 ),
    .Y(\i53/n201 ));
 INVx1_ASAP7_75t_SL \i53/i233  (.A(\i53/n533 ),
    .Y(\i53/n199 ));
 INVx1_ASAP7_75t_SL \i53/i234  (.A(\i53/n197 ),
    .Y(\i53/n198 ));
 INVx1_ASAP7_75t_SL \i53/i235  (.A(\i53/n195 ),
    .Y(\i53/n196 ));
 INVxp67_ASAP7_75t_SL \i53/i236  (.A(\i53/n191 ),
    .Y(\i53/n192 ));
 INVx1_ASAP7_75t_SL \i53/i237  (.A(\i53/n189 ),
    .Y(\i53/n190 ));
 OAI21xp33_ASAP7_75t_SL \i53/i238  (.A1(\i53/n494 ),
    .A2(\i53/n48 ),
    .B(\i53/n431 ),
    .Y(\i53/n187 ));
 NAND2xp5_ASAP7_75t_SL \i53/i239  (.A(\i53/n535 ),
    .B(\i53/n539 ),
    .Y(\i53/n186 ));
 NAND4xp75_ASAP7_75t_SL \i53/i24  (.A(\i53/n366 ),
    .B(\i53/n378 ),
    .C(\i53/n360 ),
    .D(\i53/n363 ),
    .Y(\i53/n406 ));
 OAI21xp5_ASAP7_75t_SL \i53/i240  (.A1(\i53/n514 ),
    .A2(\i53/n570 ),
    .B(\i53/n66 ),
    .Y(\i53/n185 ));
 NOR2xp33_ASAP7_75t_SL \i53/i241  (.A(\i53/n108 ),
    .B(\i53/n443 ),
    .Y(\i53/n184 ));
 NAND2xp33_ASAP7_75t_L \i53/i242  (.A(\i53/n532 ),
    .B(\i53/n561 ),
    .Y(\i53/n183 ));
 NOR2xp33_ASAP7_75t_SL \i53/i243  (.A(\i53/n573 ),
    .B(\i53/n91 ),
    .Y(\i53/n182 ));
 OAI21xp5_ASAP7_75t_SL \i53/i244  (.A1(\i53/n454 ),
    .A2(\i53/n473 ),
    .B(\i53/n420 ),
    .Y(\i53/n181 ));
 OAI21xp5_ASAP7_75t_SL \i53/i245  (.A1(\i53/n444 ),
    .A2(\i53/n425 ),
    .B(\i53/n104 ),
    .Y(\i53/n180 ));
 OA21x2_ASAP7_75t_SL \i53/i246  (.A1(\i53/n416 ),
    .A2(\i53/n8 ),
    .B(\i53/n563 ),
    .Y(\i53/n200 ));
 AOI21xp33_ASAP7_75t_SL \i53/i247  (.A1(\i53/n53 ),
    .A2(\i53/n416 ),
    .B(\i53/n37 ),
    .Y(\i53/n179 ));
 OAI21xp5_ASAP7_75t_SL \i53/i248  (.A1(\i53/n59 ),
    .A2(\i53/n70 ),
    .B(\i53/n554 ),
    .Y(\i53/n178 ));
 OAI21xp5_ASAP7_75t_SL \i53/i249  (.A1(\i53/n52 ),
    .A2(\i53/n39 ),
    .B(\i53/n554 ),
    .Y(\i53/n177 ));
 OR3x1_ASAP7_75t_SL \i53/i25  (.A(\i53/n386 ),
    .B(\i53/n384 ),
    .C(\i53/n367 ),
    .Y(\i53/n405 ));
 AOI21xp33_ASAP7_75t_SL \i53/i250  (.A1(\i53/n50 ),
    .A2(\i53/n65 ),
    .B(\i53/n37 ),
    .Y(\i53/n176 ));
 OAI21xp5_ASAP7_75t_SL \i53/i251  (.A1(\i53/n454 ),
    .A2(\i53/n425 ),
    .B(\i53/n19 ),
    .Y(\i53/n175 ));
 AOI21xp33_ASAP7_75t_SL \i53/i252  (.A1(\i53/n462 ),
    .A2(\i53/n37 ),
    .B(\i53/n54 ),
    .Y(\i53/n174 ));
 NAND2xp5_ASAP7_75t_SL \i53/i253  (.A(\i53/n554 ),
    .B(\i53/n421 ),
    .Y(\i53/n20 ));
 NAND2xp5_ASAP7_75t_L \i53/i254  (.A(\i53/n143 ),
    .B(\i53/n428 ),
    .Y(\i53/n173 ));
 OAI22xp33_ASAP7_75t_SL \i53/i255  (.A1(\i53/n71 ),
    .A2(\i53/n425 ),
    .B1(\i53/n14 ),
    .B2(\i53/n53 ),
    .Y(\i53/n197 ));
 OAI22xp5_ASAP7_75t_SL \i53/i256  (.A1(\i53/n69 ),
    .A2(\i53/n569 ),
    .B1(\i53/n454 ),
    .B2(\i53/n60 ),
    .Y(\i53/n195 ));
 OAI22xp5_ASAP7_75t_SL \i53/i257  (.A1(\i53/n54 ),
    .A2(\i53/n60 ),
    .B1(\i53/n425 ),
    .B2(\i53/n40 ),
    .Y(\i53/n194 ));
 OAI22xp5_ASAP7_75t_SL \i53/i258  (.A1(\i53/n71 ),
    .A2(\i53/n68 ),
    .B1(\i53/n38 ),
    .B2(\i53/n526 ),
    .Y(\i53/n193 ));
 OAI22xp5_ASAP7_75t_SL \i53/i259  (.A1(\i53/n454 ),
    .A2(\i53/n68 ),
    .B1(\i53/n53 ),
    .B2(\i53/n473 ),
    .Y(\i53/n191 ));
 OR3x1_ASAP7_75t_SL \i53/i26  (.A(\i53/n387 ),
    .B(\i53/n353 ),
    .C(\i53/n326 ),
    .Y(\i53/n404 ));
 NOR2x1_ASAP7_75t_SL \i53/i260  (.A(\i53/n8 ),
    .B(\i53/n16 ),
    .Y(\i53/n189 ));
 NAND2xp33_ASAP7_75t_L \i53/i261  (.A(\i53/n85 ),
    .B(\i53/n531 ),
    .Y(\i53/n172 ));
 OAI21xp5_ASAP7_75t_SL \i53/i262  (.A1(\i53/n54 ),
    .A2(\i53/n569 ),
    .B(\i53/n469 ),
    .Y(\i53/n188 ));
 INVxp67_ASAP7_75t_SL \i53/i263  (.A(\i53/n170 ),
    .Y(\i53/n171 ));
 INVxp67_ASAP7_75t_SL \i53/i264  (.A(\i53/n168 ),
    .Y(\i53/n169 ));
 INVx1_ASAP7_75t_R \i53/i265  (.A(\i53/n442 ),
    .Y(\i53/n167 ));
 INVx1_ASAP7_75t_SL \i53/i266  (.A(\i53/n165 ),
    .Y(\i53/n166 ));
 INVxp67_ASAP7_75t_SL \i53/i267  (.A(\i53/n479 ),
    .Y(\i53/n164 ));
 INVxp67_ASAP7_75t_SL \i53/i268  (.A(\i53/n160 ),
    .Y(\i53/n161 ));
 INVxp67_ASAP7_75t_SL \i53/i269  (.A(\i53/n158 ),
    .Y(\i53/n159 ));
 NAND3xp33_ASAP7_75t_SL \i53/i27  (.A(\i53/n398 ),
    .B(\i53/n383 ),
    .C(\i53/n366 ),
    .Y(\i53/n403 ));
 OAI22xp5_ASAP7_75t_SL \i53/i270  (.A1(\i53/n68 ),
    .A2(\i53/n44 ),
    .B1(\i53/n40 ),
    .B2(\i53/n8 ),
    .Y(\i53/n153 ));
 AOI21xp33_ASAP7_75t_SL \i53/i271  (.A1(\i53/n425 ),
    .A2(\i53/n60 ),
    .B(\i53/n62 ),
    .Y(\i53/n152 ));
 OAI21xp5_ASAP7_75t_SL \i53/i272  (.A1(\i53/n36 ),
    .A2(\i53/n43 ),
    .B(\i53/n41 ),
    .Y(\i53/n151 ));
 OAI22xp33_ASAP7_75t_SL \i53/i273  (.A1(\i53/n14 ),
    .A2(\i53/n48 ),
    .B1(\i53/n60 ),
    .B2(\i53/n65 ),
    .Y(\i53/n150 ));
 OAI22xp5_ASAP7_75t_SL \i53/i274  (.A1(\i53/n50 ),
    .A2(\i53/n526 ),
    .B1(\i53/n65 ),
    .B2(\i53/n462 ),
    .Y(\i53/n149 ));
 OAI22xp33_ASAP7_75t_SL \i53/i275  (.A1(\i53/n42 ),
    .A2(\i53/n48 ),
    .B1(\i53/n8 ),
    .B2(\i53/n44 ),
    .Y(\i53/n148 ));
 OAI22xp5_ASAP7_75t_SL \i53/i276  (.A1(\i53/n48 ),
    .A2(\i53/n68 ),
    .B1(\i53/n53 ),
    .B2(\i53/n8 ),
    .Y(\i53/n147 ));
 OAI21xp5_ASAP7_75t_SL \i53/i277  (.A1(\i53/n38 ),
    .A2(\i53/n569 ),
    .B(\i53/n92 ),
    .Y(\i53/n170 ));
 AOI22xp5_ASAP7_75t_SL \i53/i278  (.A1(\i53/n36 ),
    .A2(\i53/n52 ),
    .B1(\i53/n39 ),
    .B2(\i53/n570 ),
    .Y(\i53/n168 ));
 OAI22xp5_ASAP7_75t_R \i53/i279  (.A1(\i53/n37 ),
    .A2(\i53/n507 ),
    .B1(\i53/n48 ),
    .B2(\i53/n56 ),
    .Y(\i53/n146 ));
 NOR2x1_ASAP7_75t_SL \i53/i28  (.A(\i53/n307 ),
    .B(\i53/n384 ),
    .Y(\i53/n401 ));
 NAND2xp33_ASAP7_75t_SL \i53/i280  (.A(\i53/n557 ),
    .B(\i53/n144 ),
    .Y(\i53/n145 ));
 OAI22xp5_ASAP7_75t_SL \i53/i281  (.A1(\i53/n444 ),
    .A2(\i53/n68 ),
    .B1(\i53/n494 ),
    .B2(\i53/n40 ),
    .Y(\i53/n165 ));
 AO22x2_ASAP7_75t_SL \i53/i282  (.A1(\i53/n70 ),
    .A2(\i53/n67 ),
    .B1(\i53/n45 ),
    .B2(\i53/n64 ),
    .Y(\i53/n163 ));
 OAI21xp5_ASAP7_75t_SL \i53/i283  (.A1(\i53/n58 ),
    .A2(\i53/n42 ),
    .B(\i53/n458 ),
    .Y(\i53/n162 ));
 OAI22xp33_ASAP7_75t_SL \i53/i284  (.A1(\i53/n62 ),
    .A2(\i53/n37 ),
    .B1(\i53/n60 ),
    .B2(\i53/n38 ),
    .Y(\i53/n160 ));
 OAI22xp5_ASAP7_75t_SL \i53/i285  (.A1(\i53/n50 ),
    .A2(\i53/n42 ),
    .B1(\i53/n53 ),
    .B2(\i53/n60 ),
    .Y(\i53/n158 ));
 AOI22xp5_ASAP7_75t_SL \i53/i286  (.A1(\i53/n36 ),
    .A2(\i53/n41 ),
    .B1(\i53/n55 ),
    .B2(\i53/n64 ),
    .Y(\i53/n157 ));
 OAI22xp5_ASAP7_75t_SL \i53/i287  (.A1(\i53/n462 ),
    .A2(\i53/n48 ),
    .B1(\i53/n56 ),
    .B2(\i53/n416 ),
    .Y(\i53/n156 ));
 OAI22xp33_ASAP7_75t_SL \i53/i288  (.A1(\i53/n44 ),
    .A2(\i53/n47 ),
    .B1(\i53/n53 ),
    .B2(\i53/n494 ),
    .Y(\i53/n155 ));
 AOI22xp5_ASAP7_75t_SL \i53/i289  (.A1(\i53/n72 ),
    .A2(\i53/n43 ),
    .B1(\i53/n51 ),
    .B2(\i53/n57 ),
    .Y(\i53/n154 ));
 NOR2x1_ASAP7_75t_SL \i53/i29  (.A(\i53/n368 ),
    .B(\i53/n364 ),
    .Y(\i53/n400 ));
 INVxp67_ASAP7_75t_SL \i53/i290  (.A(\i53/n430 ),
    .Y(\i53/n142 ));
 INVx1_ASAP7_75t_SL \i53/i291  (.A(\i53/n140 ),
    .Y(\i53/n141 ));
 INVxp67_ASAP7_75t_SL \i53/i292  (.A(\i53/n482 ),
    .Y(\i53/n139 ));
 INVxp67_ASAP7_75t_SL \i53/i293  (.A(\i53/n137 ),
    .Y(\i53/n138 ));
 INVxp67_ASAP7_75t_SL \i53/i294  (.A(\i53/n431 ),
    .Y(\i53/n136 ));
 INVxp67_ASAP7_75t_SL \i53/i295  (.A(\i53/n524 ),
    .Y(\i53/n134 ));
 INVxp67_ASAP7_75t_SL \i53/i296  (.A(\i53/n420 ),
    .Y(\i53/n132 ));
 INVxp67_ASAP7_75t_SL \i53/i297  (.A(\i53/n532 ),
    .Y(\i53/n131 ));
 INVxp67_ASAP7_75t_SL \i53/i298  (.A(\i53/n128 ),
    .Y(\i53/n129 ));
 INVxp67_ASAP7_75t_SL \i53/i299  (.A(\i53/n471 ),
    .Y(\i53/n127 ));
 INVx1_ASAP7_75t_SL \i53/i3  (.A(\i53/n345 ),
    .Y(\i53/n3 ));
 NAND3xp33_ASAP7_75t_SL \i53/i30  (.A(\i53/n348 ),
    .B(\i53/n584 ),
    .C(\i53/n346 ),
    .Y(\i53/n399 ));
 INVxp67_ASAP7_75t_SL \i53/i300  (.A(\i53/n125 ),
    .Y(\i53/n126 ));
 INVxp67_ASAP7_75t_SL \i53/i301  (.A(\i53/n16 ),
    .Y(\i53/n124 ));
 INVx1_ASAP7_75t_SL \i53/i302  (.A(\i53/n421 ),
    .Y(\i53/n123 ));
 NAND2xp5_ASAP7_75t_SL \i53/i303  (.A(\i53/n52 ),
    .B(\i53/n554 ),
    .Y(\i53/n144 ));
 AND2x2_ASAP7_75t_SL \i53/i304  (.A(\i53/n45 ),
    .B(\i53/n57 ),
    .Y(\i53/n122 ));
 NAND2xp5_ASAP7_75t_SL \i53/i305  (.A(\i53/n66 ),
    .B(\i53/n64 ),
    .Y(\i53/n121 ));
 NAND2xp5_ASAP7_75t_SL \i53/i306  (.A(\i53/n65 ),
    .B(\i53/n62 ),
    .Y(\i53/n120 ));
 NAND2xp5_ASAP7_75t_SL \i53/i307  (.A(\i53/n39 ),
    .B(\i53/n67 ),
    .Y(\i53/n119 ));
 NAND2xp33_ASAP7_75t_SL \i53/i308  (.A(\i53/n50 ),
    .B(\i53/n454 ),
    .Y(\i53/n118 ));
 NAND2xp5_ASAP7_75t_SL \i53/i309  (.A(\i53/n5 ),
    .B(\i53/n49 ),
    .Y(\i53/n117 ));
 NOR2xp33_ASAP7_75t_L \i53/i31  (.A(\i53/n373 ),
    .B(\i53/n335 ),
    .Y(\i53/n398 ));
 NAND2xp5_ASAP7_75t_SL \i53/i310  (.A(\i53/n52 ),
    .B(\i53/n5 ),
    .Y(\i53/n116 ));
 NAND2xp5_ASAP7_75t_SL \i53/i311  (.A(\i53/n57 ),
    .B(\i53/n55 ),
    .Y(\i53/n115 ));
 NAND2xp5_ASAP7_75t_SL \i53/i312  (.A(\i53/n36 ),
    .B(\i53/n45 ),
    .Y(\i53/n114 ));
 NAND2xp5_ASAP7_75t_SL \i53/i313  (.A(\i53/n36 ),
    .B(\i53/n59 ),
    .Y(\i53/n143 ));
 AND2x2_ASAP7_75t_SL \i53/i314  (.A(\i53/n72 ),
    .B(\i53/n57 ),
    .Y(\i53/n140 ));
 NAND2xp5_ASAP7_75t_SL \i53/i315  (.A(\i53/n57 ),
    .B(\i53/n7 ),
    .Y(\i53/n19 ));
 NAND2xp5_ASAP7_75t_SL \i53/i316  (.A(\i53/n70 ),
    .B(\i53/n43 ),
    .Y(\i53/n137 ));
 AND2x2_ASAP7_75t_SL \i53/i317  (.A(\i53/n52 ),
    .B(\i53/n46 ),
    .Y(\i53/n135 ));
 NOR2xp67_ASAP7_75t_SL \i53/i318  (.A(\i53/n416 ),
    .B(\i53/n425 ),
    .Y(\i53/n18 ));
 NOR2xp33_ASAP7_75t_SL \i53/i319  (.A(\i53/n54 ),
    .B(\i53/n60 ),
    .Y(\i53/n113 ));
 NOR5xp2_ASAP7_75t_SL \i53/i32  (.A(\i53/n337 ),
    .B(\i53/n284 ),
    .C(\i53/n328 ),
    .D(\i53/n252 ),
    .E(\i53/n256 ),
    .Y(\i53/n397 ));
 NAND2xp5_ASAP7_75t_SL \i53/i320  (.A(\i53/n46 ),
    .B(\i53/n49 ),
    .Y(\i53/n112 ));
 NOR2xp33_ASAP7_75t_SL \i53/i321  (.A(\i53/n48 ),
    .B(\i53/n60 ),
    .Y(\i53/n133 ));
 NOR2xp33_ASAP7_75t_SL \i53/i322  (.A(\i53/n444 ),
    .B(\i53/n8 ),
    .Y(\i53/n111 ));
 NOR2xp33_ASAP7_75t_SL \i53/i323  (.A(\i53/n51 ),
    .B(\i53/n66 ),
    .Y(\i53/n110 ));
 NOR2xp33_ASAP7_75t_SL \i53/i324  (.A(\i53/n48 ),
    .B(\i53/n473 ),
    .Y(\i53/n109 ));
 NOR2xp33_ASAP7_75t_L \i53/i325  (.A(\i53/n70 ),
    .B(\i53/n41 ),
    .Y(\i53/n130 ));
 NAND2xp5_ASAP7_75t_SL \i53/i326  (.A(\i53/n51 ),
    .B(\i53/n61 ),
    .Y(\i53/n17 ));
 NAND2xp5_ASAP7_75t_SL \i53/i327  (.A(\i53/n70 ),
    .B(\i53/n570 ),
    .Y(\i53/n128 ));
 NOR2xp67_ASAP7_75t_SL \i53/i328  (.A(\i53/n66 ),
    .B(\i53/n52 ),
    .Y(\i53/n125 ));
 NOR2xp33_ASAP7_75t_SL \i53/i329  (.A(\i53/n569 ),
    .B(\i53/n65 ),
    .Y(\i53/n108 ));
 NOR3xp33_ASAP7_75t_SL \i53/i33  (.A(\i53/n333 ),
    .B(\i53/n350 ),
    .C(\i53/n382 ),
    .Y(\i53/n396 ));
 NOR2x1_ASAP7_75t_SL \i53/i330  (.A(\i53/n51 ),
    .B(\i53/n63 ),
    .Y(\i53/n16 ));
 INVxp67_ASAP7_75t_SL \i53/i331  (.A(\i53/n106 ),
    .Y(\i53/n107 ));
 INVxp67_ASAP7_75t_SL \i53/i332  (.A(\i53/n104 ),
    .Y(\i53/n105 ));
 INVx1_ASAP7_75t_SL \i53/i333  (.A(\i53/n433 ),
    .Y(\i53/n103 ));
 INVxp67_ASAP7_75t_SL \i53/i334  (.A(\i53/n484 ),
    .Y(\i53/n100 ));
 INVxp67_ASAP7_75t_SL \i53/i335  (.A(\i53/n98 ),
    .Y(\i53/n99 ));
 INVxp67_ASAP7_75t_SL \i53/i336  (.A(\i53/n545 ),
    .Y(\i53/n97 ));
 INVxp67_ASAP7_75t_SL \i53/i337  (.A(\i53/n95 ),
    .Y(\i53/n96 ));
 INVxp67_ASAP7_75t_SL \i53/i338  (.A(\i53/n93 ),
    .Y(\i53/n94 ));
 INVxp67_ASAP7_75t_SL \i53/i339  (.A(\i53/n91 ),
    .Y(\i53/n92 ));
 NOR2x1_ASAP7_75t_SL \i53/i34  (.A(\i53/n379 ),
    .B(\i53/n338 ),
    .Y(\i53/n395 ));
 INVxp67_ASAP7_75t_SL \i53/i340  (.A(\i53/n450 ),
    .Y(\i53/n86 ));
 INVx1_ASAP7_75t_SL \i53/i341  (.A(\i53/n449 ),
    .Y(\i53/n84 ));
 NAND2xp5_ASAP7_75t_SL \i53/i342  (.A(\i53/n58 ),
    .B(\i53/n54 ),
    .Y(\i53/n83 ));
 NAND2xp5_ASAP7_75t_SL \i53/i343  (.A(\i53/n59 ),
    .B(\i53/n46 ),
    .Y(\i53/n82 ));
 NAND2xp5_ASAP7_75t_SL \i53/i344  (.A(\i53/n55 ),
    .B(\i53/n570 ),
    .Y(\i53/n81 ));
 NAND2xp5_ASAP7_75t_L \i53/i345  (.A(\i53/n14 ),
    .B(\i53/n37 ),
    .Y(\i53/n80 ));
 NAND2xp33_ASAP7_75t_SL \i53/i346  (.A(\i53/n47 ),
    .B(\i53/n526 ),
    .Y(\i53/n79 ));
 NAND2xp5_ASAP7_75t_SL \i53/i347  (.A(\i53/n72 ),
    .B(\i53/n514 ),
    .Y(\i53/n106 ));
 NOR2xp33_ASAP7_75t_SL \i53/i348  (.A(\i53/n569 ),
    .B(\i53/n454 ),
    .Y(\i53/n78 ));
 NAND2xp5_ASAP7_75t_SL \i53/i349  (.A(\i53/n66 ),
    .B(\i53/n46 ),
    .Y(\i53/n104 ));
 NAND2xp5_ASAP7_75t_SL \i53/i35  (.A(\i53/n336 ),
    .B(\i53/n356 ),
    .Y(\i53/n394 ));
 NAND2xp5_ASAP7_75t_SL \i53/i350  (.A(\i53/n7 ),
    .B(\i53/n61 ),
    .Y(\i53/n102 ));
 AND2x2_ASAP7_75t_SL \i53/i351  (.A(\i53/n7 ),
    .B(\i53/n43 ),
    .Y(\i53/n101 ));
 NAND2xp5_ASAP7_75t_SL \i53/i352  (.A(\i53/n63 ),
    .B(\i53/n43 ),
    .Y(\i53/n98 ));
 NAND2xp5_ASAP7_75t_SL \i53/i353  (.A(\i53/n39 ),
    .B(\i53/n43 ),
    .Y(\i53/n95 ));
 NAND2xp33_ASAP7_75t_L \i53/i354  (.A(\i53/n42 ),
    .B(\i53/n494 ),
    .Y(\i53/n77 ));
 NAND2xp5_ASAP7_75t_SL \i53/i355  (.A(\i53/n36 ),
    .B(\i53/n72 ),
    .Y(\i53/n93 ));
 NOR2xp67_ASAP7_75t_L \i53/i356  (.A(\i53/n37 ),
    .B(\i53/n454 ),
    .Y(\i53/n91 ));
 NAND2xp5_ASAP7_75t_SL \i53/i357  (.A(\i53/n41 ),
    .B(\i53/n61 ),
    .Y(\i53/n15 ));
 NAND2xp5_ASAP7_75t_SL \i53/i358  (.A(\i53/n41 ),
    .B(\i53/n64 ),
    .Y(\i53/n90 ));
 AND2x2_ASAP7_75t_SL \i53/i359  (.A(\i53/n72 ),
    .B(\i53/n64 ),
    .Y(\i53/n89 ));
 NOR3x1_ASAP7_75t_SL \i53/i36  (.A(\i53/n23 ),
    .B(\i53/n352 ),
    .C(\i53/n277 ),
    .Y(\i53/n402 ));
 NAND2xp5_ASAP7_75t_L \i53/i360  (.A(\i53/n8 ),
    .B(\i53/n14 ),
    .Y(\i53/n88 ));
 AND2x2_ASAP7_75t_SL \i53/i361  (.A(\i53/n72 ),
    .B(\i53/n46 ),
    .Y(\i53/n87 ));
 NOR2xp33_ASAP7_75t_SL \i53/i362  (.A(\i53/n47 ),
    .B(\i53/n38 ),
    .Y(\i53/n76 ));
 NAND2xp5_ASAP7_75t_SL \i53/i363  (.A(\i53/n7 ),
    .B(\i53/n64 ),
    .Y(\i53/n75 ));
 NAND2xp5_ASAP7_75t_SL \i53/i364  (.A(\i53/n59 ),
    .B(\i53/n64 ),
    .Y(\i53/n85 ));
 NOR2xp33_ASAP7_75t_SL \i53/i365  (.A(\i53/n71 ),
    .B(\i53/n8 ),
    .Y(\i53/n74 ));
 NOR2xp33_ASAP7_75t_SL \i53/i366  (.A(\i53/n71 ),
    .B(\i53/n569 ),
    .Y(\i53/n73 ));
 INVx2_ASAP7_75t_SL \i53/i367  (.A(\i53/n72 ),
    .Y(\i53/n71 ));
 INVx1_ASAP7_75t_SL \i53/i368  (.A(\i53/n70 ),
    .Y(\i53/n69 ));
 INVx3_ASAP7_75t_SL \i53/i369  (.A(\i53/n68 ),
    .Y(\i53/n67 ));
 NOR3xp33_ASAP7_75t_SL \i53/i37  (.A(\i53/n294 ),
    .B(\i53/n23 ),
    .C(\i53/n376 ),
    .Y(\i53/n392 ));
 INVx3_ASAP7_75t_SL \i53/i370  (.A(\i53/n66 ),
    .Y(\i53/n65 ));
 INVx2_ASAP7_75t_SL \i53/i371  (.A(\i53/n63 ),
    .Y(\i53/n62 ));
 INVx4_ASAP7_75t_SL \i53/i372  (.A(\i53/n61 ),
    .Y(\i53/n60 ));
 INVx2_ASAP7_75t_SL \i53/i373  (.A(\i53/n59 ),
    .Y(\i53/n58 ));
 INVx3_ASAP7_75t_SL \i53/i374  (.A(\i53/n57 ),
    .Y(\i53/n56 ));
 INVx3_ASAP7_75t_SL \i53/i375  (.A(\i53/n55 ),
    .Y(\i53/n54 ));
 INVx3_ASAP7_75t_SL \i53/i376  (.A(\i53/n53 ),
    .Y(\i53/n52 ));
 AND2x4_ASAP7_75t_SL \i53/i377  (.A(\i53/n436 ),
    .B(\i53/n34 ),
    .Y(\i53/n72 ));
 AND2x4_ASAP7_75t_SL \i53/i378  (.A(\i53/n414 ),
    .B(\i53/n436 ),
    .Y(\i53/n70 ));
 OR2x4_ASAP7_75t_SL \i53/i379  (.A(\i53/n29 ),
    .B(\i53/n9 ),
    .Y(\i53/n68 ));
 NOR2xp33_ASAP7_75t_SL \i53/i38  (.A(\i53/n357 ),
    .B(\i53/n23 ),
    .Y(\i53/n391 ));
 AND2x4_ASAP7_75t_SL \i53/i380  (.A(\i53/n28 ),
    .B(\i53/n437 ),
    .Y(\i53/n66 ));
 AND2x4_ASAP7_75t_SL \i53/i381  (.A(\i53/n456 ),
    .B(\i53/n30 ),
    .Y(\i53/n64 ));
 NAND2x1_ASAP7_75t_SL \i53/i382  (.A(\i53/n456 ),
    .B(\i53/n30 ),
    .Y(\i53/n14 ));
 AND2x4_ASAP7_75t_SL \i53/i383  (.A(\i53/n28 ),
    .B(\i53/n414 ),
    .Y(\i53/n63 ));
 AND2x4_ASAP7_75t_SL \i53/i384  (.A(\i53/n35 ),
    .B(\i53/n422 ),
    .Y(\i53/n61 ));
 AND2x4_ASAP7_75t_SL \i53/i385  (.A(\i53/n28 ),
    .B(\i53/n446 ),
    .Y(\i53/n59 ));
 AND2x4_ASAP7_75t_SL \i53/i386  (.A(\i53/n485 ),
    .B(\i53/n456 ),
    .Y(\i53/n57 ));
 AND2x4_ASAP7_75t_SL \i53/i387  (.A(\i53/n414 ),
    .B(\i53/n32 ),
    .Y(\i53/n55 ));
 OR2x6_ASAP7_75t_SL \i53/i388  (.A(\i53/n33 ),
    .B(\i53/n27 ),
    .Y(\i53/n53 ));
 INVx3_ASAP7_75t_SL \i53/i389  (.A(\i53/n51 ),
    .Y(\i53/n50 ));
 NOR3xp33_ASAP7_75t_SL \i53/i39  (.A(\i53/n334 ),
    .B(\i53/n329 ),
    .C(\i53/n3 ),
    .Y(\i53/n390 ));
 INVx3_ASAP7_75t_SL \i53/i390  (.A(\i53/n49 ),
    .Y(\i53/n48 ));
 INVx4_ASAP7_75t_SL \i53/i391  (.A(\i53/n47 ),
    .Y(\i53/n46 ));
 INVx4_ASAP7_75t_SL \i53/i392  (.A(\i53/n45 ),
    .Y(\i53/n44 ));
 INVx3_ASAP7_75t_SL \i53/i393  (.A(\i53/n41 ),
    .Y(\i53/n40 ));
 INVx4_ASAP7_75t_SL \i53/i394  (.A(\i53/n39 ),
    .Y(\i53/n38 ));
 INVx3_ASAP7_75t_SL \i53/i395  (.A(\i53/n37 ),
    .Y(\i53/n36 ));
 AND2x4_ASAP7_75t_SL \i53/i396  (.A(\i53/n34 ),
    .B(\i53/n32 ),
    .Y(\i53/n51 ));
 AND2x4_ASAP7_75t_SL \i53/i397  (.A(\i53/n446 ),
    .B(\i53/n436 ),
    .Y(\i53/n49 ));
 NAND2x1p5_ASAP7_75t_SL \i53/i398  (.A(\i53/n485 ),
    .B(\i53/n35 ),
    .Y(\i53/n47 ));
 AND2x4_ASAP7_75t_SL \i53/i399  (.A(\i53/n34 ),
    .B(\i53/n447 ),
    .Y(\i53/n45 ));
 INVx2_ASAP7_75t_SL \i53/i4  (.A(\i53/n511 ),
    .Y(\i53/n4 ));
 NAND4xp25_ASAP7_75t_SL \i53/i40  (.A(\i53/n317 ),
    .B(\i53/n311 ),
    .C(\i53/n310 ),
    .D(\i53/n343 ),
    .Y(\i53/n389 ));
 AND2x4_ASAP7_75t_SL \i53/i400  (.A(\i53/n4 ),
    .B(\i53/n30 ),
    .Y(\i53/n43 ));
 NAND2x1_ASAP7_75t_SL \i53/i401  (.A(\i53/n4 ),
    .B(\i53/n30 ),
    .Y(\i53/n42 ));
 AND2x4_ASAP7_75t_SL \i53/i402  (.A(\i53/n446 ),
    .B(\i53/n32 ),
    .Y(\i53/n41 ));
 AND2x4_ASAP7_75t_SL \i53/i403  (.A(\i53/n437 ),
    .B(\i53/n32 ),
    .Y(\i53/n39 ));
 OR2x6_ASAP7_75t_SL \i53/i404  (.A(\i53/n26 ),
    .B(\i53/n31 ),
    .Y(\i53/n37 ));
 INVx3_ASAP7_75t_SL \i53/i405  (.A(\i53/n33 ),
    .Y(\i53/n34 ));
 NAND2xp5_ASAP7_75t_SL \i53/i406  (.A(\i53/n12 ),
    .B(\i53/n1 ),
    .Y(\i53/n31 ));
 AND2x2_ASAP7_75t_SL \i53/i407  (.A(\i53/n12 ),
    .B(\i53/n1 ),
    .Y(\i53/n35 ));
 NAND2x1p5_ASAP7_75t_SL \i53/i408  (.A(n15[4]),
    .B(n15[5]),
    .Y(\i53/n33 ));
 AND2x4_ASAP7_75t_SL \i53/i409  (.A(n15[7]),
    .B(\i53/n13 ),
    .Y(\i53/n32 ));
 NAND3xp33_ASAP7_75t_L \i53/i41  (.A(\i53/n291 ),
    .B(\i53/n311 ),
    .C(\i53/n361 ),
    .Y(\i53/n388 ));
 INVx2_ASAP7_75t_SL \i53/i410  (.A(\i53/n9 ),
    .Y(\i53/n30 ));
 INVx2_ASAP7_75t_SL \i53/i411  (.A(\i53/n28 ),
    .Y(\i53/n27 ));
 NAND2xp5_ASAP7_75t_SL \i53/i412  (.A(\i53/n25 ),
    .B(\i53/n2 ),
    .Y(\i53/n26 ));
 NAND2x1_ASAP7_75t_SL \i53/i413  (.A(n15[3]),
    .B(\i53/n1 ),
    .Y(\i53/n29 ));
 AND2x2_ASAP7_75t_SL \i53/i414  (.A(n15[7]),
    .B(n15[6]),
    .Y(\i53/n28 ));
 INVx1_ASAP7_75t_SL \i53/i415  (.A(n15[1]),
    .Y(\i53/n25 ));
 INVx3_ASAP7_75t_SL \i53/i416  (.A(n15[5]),
    .Y(\i53/n24 ));
 INVx2_ASAP7_75t_SL \i53/i417  (.A(n15[6]),
    .Y(\i53/n13 ));
 INVx2_ASAP7_75t_SL \i53/i418  (.A(n15[3]),
    .Y(\i53/n12 ));
 INVx2_ASAP7_75t_SL \i53/i419  (.A(n15[4]),
    .Y(\i53/n11 ));
 NAND3xp33_ASAP7_75t_SL \i53/i42  (.A(\i53/n296 ),
    .B(\i53/n345 ),
    .C(\i53/n330 ),
    .Y(\i53/n387 ));
 OR2x2_ASAP7_75t_SL \i53/i420  (.A(\i53/n101 ),
    .B(\i53/n522 ),
    .Y(\i53/n10 ));
 OR2x2_ASAP7_75t_SL \i53/i421  (.A(n15[0]),
    .B(n15[1]),
    .Y(\i53/n9 ));
 AND2x2_ASAP7_75t_SL \i53/i422  (.A(\i53/n24 ),
    .B(\i53/n11 ),
    .Y(\i53/n414 ));
 AND2x4_ASAP7_75t_SL \i53/i423  (.A(\i53/n414 ),
    .B(\i53/n447 ),
    .Y(\i53/n415 ));
 INVx3_ASAP7_75t_SL \i53/i424  (.A(\i53/n415 ),
    .Y(\i53/n416 ));
 AOI211x1_ASAP7_75t_SL \i53/i425  (.A1(\i53/n80 ),
    .A2(\i53/n415 ),
    .B(\i53/n430 ),
    .C(\i53/n501 ),
    .Y(\i53/n417 ));
 AOI22xp5_ASAP7_75t_SL \i53/i426  (.A1(\i53/n415 ),
    .A2(\i53/n67 ),
    .B1(\i53/n7 ),
    .B2(\i53/n64 ),
    .Y(\i53/n418 ));
 NAND2xp5_ASAP7_75t_SL \i53/i427  (.A(\i53/n415 ),
    .B(\i53/n5 ),
    .Y(\i53/n419 ));
 NAND2xp5_ASAP7_75t_SL \i53/i428  (.A(\i53/n415 ),
    .B(\i53/n43 ),
    .Y(\i53/n420 ));
 OR2x2_ASAP7_75t_SL \i53/i429  (.A(\i53/n41 ),
    .B(\i53/n415 ),
    .Y(\i53/n421 ));
 NAND2xp5_ASAP7_75t_L \i53/i43  (.A(\i53/n344 ),
    .B(\i53/n377 ),
    .Y(\i53/n386 ));
 INVx2_ASAP7_75t_SL \i53/i430  (.A(\i53/n512 ),
    .Y(\i53/n422 ));
 AND2x4_ASAP7_75t_SL \i53/i431  (.A(\i53/n456 ),
    .B(\i53/n422 ),
    .Y(\i53/n423 ));
 OAI21xp5_ASAP7_75t_SL \i53/i432  (.A1(\i53/n423 ),
    .A2(\i53/n556 ),
    .B(\i53/n41 ),
    .Y(\i53/n424 ));
 INVx4_ASAP7_75t_SL \i53/i433  (.A(\i53/n423 ),
    .Y(\i53/n425 ));
 AOI211x1_ASAP7_75t_L \i53/i434  (.A1(\i53/n423 ),
    .A2(\i53/n52 ),
    .B(\i53/n443 ),
    .C(\i53/n534 ),
    .Y(\i53/n426 ));
 OAI21xp5_ASAP7_75t_SL \i53/i435  (.A1(\i53/n423 ),
    .A2(\i53/n46 ),
    .B(\i53/n59 ),
    .Y(\i53/n427 ));
 NAND2xp5_ASAP7_75t_SL \i53/i436  (.A(\i53/n49 ),
    .B(\i53/n423 ),
    .Y(\i53/n428 ));
 NAND2xp5_ASAP7_75t_SL \i53/i437  (.A(\i53/n45 ),
    .B(\i53/n423 ),
    .Y(\i53/n429 ));
 AND2x2_ASAP7_75t_SL \i53/i438  (.A(\i53/n66 ),
    .B(\i53/n423 ),
    .Y(\i53/n430 ));
 NAND2xp5_ASAP7_75t_SL \i53/i439  (.A(\i53/n51 ),
    .B(\i53/n423 ),
    .Y(\i53/n431 ));
 NAND2xp33_ASAP7_75t_SL \i53/i44  (.A(\i53/n341 ),
    .B(\i53/n359 ),
    .Y(\i53/n385 ));
 NAND2xp5_ASAP7_75t_SL \i53/i440  (.A(\i53/n39 ),
    .B(\i53/n423 ),
    .Y(\i53/n432 ));
 NOR2xp33_ASAP7_75t_SL \i53/i441  (.A(\i53/n423 ),
    .B(\i53/n64 ),
    .Y(\i53/n433 ));
 OAI221xp5_ASAP7_75t_SL \i53/i442  (.A1(\i53/n504 ),
    .A2(\i53/n69 ),
    .B1(\i53/n504 ),
    .B2(\i53/n507 ),
    .C(\i53/n417 ),
    .Y(\i53/n434 ));
 NAND2xp5_ASAP7_75t_SL \i53/i443  (.A(\i53/n448 ),
    .B(\i53/n61 ),
    .Y(\i53/n435 ));
 AND2x2_ASAP7_75t_SL \i53/i444  (.A(\i53/n0 ),
    .B(\i53/n13 ),
    .Y(\i53/n436 ));
 INVx2_ASAP7_75t_SL \i53/i445  (.A(\i53/n505 ),
    .Y(\i53/n437 ));
 AND2x4_ASAP7_75t_SL \i53/i446  (.A(\i53/n436 ),
    .B(\i53/n437 ),
    .Y(\i53/n438 ));
 AOI22xp5_ASAP7_75t_SL \i53/i447  (.A1(\i53/n438 ),
    .A2(\i53/n61 ),
    .B1(\i53/n39 ),
    .B2(\i53/n64 ),
    .Y(\i53/n439 ));
 AOI221xp5_ASAP7_75t_SL \i53/i448  (.A1(\i53/n438 ),
    .A2(\i53/n36 ),
    .B1(\i53/n43 ),
    .B2(\i53/n52 ),
    .C(\i53/n523 ),
    .Y(\i53/n440 ));
 NAND2xp5_ASAP7_75t_SL \i53/i449  (.A(\i53/n438 ),
    .B(\i53/n57 ),
    .Y(\i53/n441 ));
 NOR2x1_ASAP7_75t_SL \i53/i45  (.A(\i53/n358 ),
    .B(\i53/n367 ),
    .Y(\i53/n393 ));
 AOI22xp5_ASAP7_75t_SL \i53/i450  (.A1(\i53/n41 ),
    .A2(\i53/n43 ),
    .B1(\i53/n46 ),
    .B2(\i53/n438 ),
    .Y(\i53/n442 ));
 AND2x2_ASAP7_75t_SL \i53/i451  (.A(\i53/n438 ),
    .B(\i53/n5 ),
    .Y(\i53/n443 ));
 INVx3_ASAP7_75t_SL \i53/i452  (.A(\i53/n438 ),
    .Y(\i53/n444 ));
 NAND2xp5_ASAP7_75t_SL \i53/i453  (.A(\i53/n438 ),
    .B(\i53/n554 ),
    .Y(\i53/n445 ));
 AND2x2_ASAP7_75t_SL \i53/i454  (.A(n15[4]),
    .B(\i53/n24 ),
    .Y(\i53/n446 ));
 AND2x2_ASAP7_75t_L \i53/i455  (.A(\i53/n0 ),
    .B(n15[6]),
    .Y(\i53/n447 ));
 NAND2x1_ASAP7_75t_SL \i53/i456  (.A(\i53/n448 ),
    .B(\i53/n554 ),
    .Y(\i53/n449 ));
 AND2x4_ASAP7_75t_SL \i53/i457  (.A(\i53/n446 ),
    .B(\i53/n447 ),
    .Y(\i53/n448 ));
 NAND2xp5_ASAP7_75t_SL \i53/i458  (.A(\i53/n448 ),
    .B(\i53/n570 ),
    .Y(\i53/n450 ));
 AOI22xp5_ASAP7_75t_SL \i53/i459  (.A1(\i53/n448 ),
    .A2(\i53/n64 ),
    .B1(\i53/n39 ),
    .B2(\i53/n46 ),
    .Y(\i53/n451 ));
 NAND2xp33_ASAP7_75t_L \i53/i46  (.A(\i53/n347 ),
    .B(\i53/n319 ),
    .Y(\i53/n382 ));
 OAI21xp5_ASAP7_75t_SL \i53/i460  (.A1(\i53/n63 ),
    .A2(\i53/n448 ),
    .B(\i53/n514 ),
    .Y(\i53/n452 ));
 OAI21xp5_ASAP7_75t_SL \i53/i461  (.A1(\i53/n514 ),
    .A2(\i53/n43 ),
    .B(\i53/n448 ),
    .Y(\i53/n453 ));
 INVx5_ASAP7_75t_SL \i53/i462  (.A(\i53/n448 ),
    .Y(\i53/n454 ));
 OAI21xp5_ASAP7_75t_SL \i53/i463  (.A1(\i53/n448 ),
    .A2(\i53/n55 ),
    .B(\i53/n423 ),
    .Y(\i53/n455 ));
 AND2x4_ASAP7_75t_SL \i53/i464  (.A(n15[2]),
    .B(n15[3]),
    .Y(\i53/n456 ));
 NAND2xp5_ASAP7_75t_SL \i53/i465  (.A(\i53/n448 ),
    .B(\i53/n457 ),
    .Y(\i53/n458 ));
 AND2x4_ASAP7_75t_SL \i53/i466  (.A(\i53/n456 ),
    .B(\i53/n555 ),
    .Y(\i53/n457 ));
 AOI222xp33_ASAP7_75t_SL \i53/i467  (.A1(\i53/n457 ),
    .A2(\i53/n438 ),
    .B1(\i53/n7 ),
    .B2(\i53/n36 ),
    .C1(\i53/n57 ),
    .C2(\i53/n49 ),
    .Y(\i53/n459 ));
 AOI221xp5_ASAP7_75t_SL \i53/i468  (.A1(\i53/n457 ),
    .A2(\i53/n70 ),
    .B1(\i53/n514 ),
    .B2(\i53/n438 ),
    .C(\i53/n146 ),
    .Y(\i53/n460 ));
 NAND2xp5_ASAP7_75t_SL \i53/i469  (.A(\i53/n457 ),
    .B(\i53/n415 ),
    .Y(\i53/n461 ));
 NAND2xp33_ASAP7_75t_L \i53/i47  (.A(\i53/n344 ),
    .B(\i53/n324 ),
    .Y(\i53/n381 ));
 INVx3_ASAP7_75t_SL \i53/i470  (.A(\i53/n457 ),
    .Y(\i53/n462 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i53/i471  (.A1(\i53/n457 ),
    .A2(\i53/n77 ),
    .B(\i53/n59 ),
    .C(\i53/n202 ),
    .Y(\i53/n463 ));
 AOI221x1_ASAP7_75t_SL \i53/i472  (.A1(\i53/n67 ),
    .A2(\i53/n55 ),
    .B1(\i53/n457 ),
    .B2(\i53/n59 ),
    .C(\i53/n478 ),
    .Y(\i53/n464 ));
 NAND2xp5_ASAP7_75t_SL \i53/i473  (.A(\i53/n52 ),
    .B(\i53/n457 ),
    .Y(\i53/n465 ));
 NAND2xp5_ASAP7_75t_SL \i53/i474  (.A(\i53/n41 ),
    .B(\i53/n457 ),
    .Y(\i53/n466 ));
 NAND2xp5_ASAP7_75t_SL \i53/i475  (.A(\i53/n457 ),
    .B(\i53/n39 ),
    .Y(\i53/n467 ));
 AND2x2_ASAP7_75t_SL \i53/i476  (.A(\i53/n7 ),
    .B(\i53/n457 ),
    .Y(\i53/n468 ));
 NAND2xp5_ASAP7_75t_SL \i53/i477  (.A(\i53/n72 ),
    .B(\i53/n457 ),
    .Y(\i53/n469 ));
 NAND2xp5_ASAP7_75t_SL \i53/i478  (.A(\i53/n470 ),
    .B(\i53/n438 ),
    .Y(\i53/n471 ));
 AND2x4_ASAP7_75t_SL \i53/i479  (.A(\i53/n4 ),
    .B(\i53/n485 ),
    .Y(\i53/n470 ));
 NOR2xp67_ASAP7_75t_SL \i53/i48  (.A(\i53/n323 ),
    .B(\i53/n349 ),
    .Y(\i53/n380 ));
 AOI22xp5_ASAP7_75t_SL \i53/i480  (.A1(\i53/n470 ),
    .A2(\i53/n72 ),
    .B1(\i53/n63 ),
    .B2(\i53/n57 ),
    .Y(\i53/n472 ));
 INVx3_ASAP7_75t_SL \i53/i481  (.A(\i53/n470 ),
    .Y(\i53/n473 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i53/i482  (.A1(\i53/n470 ),
    .A2(\i53/n43 ),
    .B(\i53/n55 ),
    .C(\i53/n468 ),
    .Y(\i53/n474 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i53/i483  (.A1(\i53/n66 ),
    .A2(\i53/n7 ),
    .B(\i53/n470 ),
    .C(\i53/n573 ),
    .Y(\i53/n475 ));
 AOI21xp5_ASAP7_75t_SL \i53/i484  (.A1(\i53/n421 ),
    .A2(\i53/n470 ),
    .B(\i53/n175 ),
    .Y(\i53/n476 ));
 AOI22xp5_ASAP7_75t_R \i53/i485  (.A1(\i53/n554 ),
    .A2(\i53/n120 ),
    .B1(\i53/n49 ),
    .B2(\i53/n470 ),
    .Y(\i53/n477 ));
 OA21x2_ASAP7_75t_SL \i53/i486  (.A1(\i53/n7 ),
    .A2(\i53/n70 ),
    .B(\i53/n470 ),
    .Y(\i53/n478 ));
 AOI22xp5_ASAP7_75t_SL \i53/i487  (.A1(\i53/n41 ),
    .A2(\i53/n46 ),
    .B1(\i53/n39 ),
    .B2(\i53/n470 ),
    .Y(\i53/n479 ));
 NAND2xp5_ASAP7_75t_SL \i53/i488  (.A(\i53/n66 ),
    .B(\i53/n470 ),
    .Y(\i53/n480 ));
 NAND2xp5_ASAP7_75t_SL \i53/i489  (.A(\i53/n52 ),
    .B(\i53/n470 ),
    .Y(\i53/n481 ));
 NAND3xp33_ASAP7_75t_SL \i53/i49  (.A(\i53/n314 ),
    .B(\i53/n426 ),
    .C(\i53/n321 ),
    .Y(\i53/n379 ));
 NAND2xp5_ASAP7_75t_SL \i53/i490  (.A(\i53/n59 ),
    .B(\i53/n470 ),
    .Y(\i53/n482 ));
 NOR2xp67_ASAP7_75t_L \i53/i491  (.A(\i53/n470 ),
    .B(\i53/n61 ),
    .Y(\i53/n483 ));
 NAND2xp5_ASAP7_75t_SL \i53/i492  (.A(\i53/n63 ),
    .B(\i53/n470 ),
    .Y(\i53/n484 ));
 AND2x2_ASAP7_75t_SL \i53/i493  (.A(n15[0]),
    .B(n15[1]),
    .Y(\i53/n485 ));
 OAI21xp33_ASAP7_75t_SL \i53/i494  (.A1(\i53/n470 ),
    .A2(\i53/n486 ),
    .B(\i53/n41 ),
    .Y(\i53/n487 ));
 AND2x4_ASAP7_75t_SL \i53/i495  (.A(\i53/n485 ),
    .B(\i53/n6 ),
    .Y(\i53/n486 ));
 AOI22xp5_ASAP7_75t_SL \i53/i496  (.A1(\i53/n486 ),
    .A2(\i53/n83 ),
    .B1(\i53/n63 ),
    .B2(\i53/n457 ),
    .Y(\i53/n488 ));
 OAI31xp33_ASAP7_75t_R \i53/i497  (.A1(\i53/n57 ),
    .A2(\i53/n486 ),
    .A3(\i53/n457 ),
    .B(\i53/n55 ),
    .Y(\i53/n489 ));
 NAND2xp5_ASAP7_75t_SL \i53/i498  (.A(\i53/n448 ),
    .B(\i53/n486 ),
    .Y(\i53/n490 ));
 OAI21xp5_ASAP7_75t_SL \i53/i499  (.A1(\i53/n486 ),
    .A2(\i53/n64 ),
    .B(\i53/n438 ),
    .Y(\i53/n491 ));
 INVx2_ASAP7_75t_SL \i53/i5  (.A(\i53/n526 ),
    .Y(\i53/n5 ));
 NOR2x1_ASAP7_75t_SL \i53/i50  (.A(\i53/n271 ),
    .B(\i53/n332 ),
    .Y(\i53/n378 ));
 OAI21xp5_ASAP7_75t_SL \i53/i500  (.A1(\i53/n486 ),
    .A2(\i53/n423 ),
    .B(\i53/n70 ),
    .Y(\i53/n492 ));
 AOI22xp33_ASAP7_75t_SL \i53/i501  (.A1(\i53/n415 ),
    .A2(\i53/n486 ),
    .B1(\i53/n7 ),
    .B2(\i53/n514 ),
    .Y(\i53/n493 ));
 INVx2_ASAP7_75t_SL \i53/i502  (.A(\i53/n486 ),
    .Y(\i53/n494 ));
 AOI21xp5_ASAP7_75t_SL \i53/i503  (.A1(\i53/n486 ),
    .A2(\i53/n51 ),
    .B(\i53/n191 ),
    .Y(\i53/n495 ));
 OAI21xp5_ASAP7_75t_SL \i53/i504  (.A1(\i53/n88 ),
    .A2(\i53/n486 ),
    .B(\i53/n63 ),
    .Y(\i53/n496 ));
 OAI21xp5_ASAP7_75t_SL \i53/i505  (.A1(\i53/n486 ),
    .A2(\i53/n570 ),
    .B(\i53/n52 ),
    .Y(\i53/n497 ));
 AOI22xp5_ASAP7_75t_R \i53/i506  (.A1(\i53/n36 ),
    .A2(\i53/n70 ),
    .B1(\i53/n39 ),
    .B2(\i53/n486 ),
    .Y(\i53/n498 ));
 OAI21xp33_ASAP7_75t_SL \i53/i507  (.A1(\i53/n486 ),
    .A2(\i53/n43 ),
    .B(\i53/n66 ),
    .Y(\i53/n499 ));
 AOI22xp5_ASAP7_75t_SL \i53/i508  (.A1(\i53/n36 ),
    .A2(\i53/n39 ),
    .B1(\i53/n72 ),
    .B2(\i53/n486 ),
    .Y(\i53/n500 ));
 AND2x2_ASAP7_75t_SL \i53/i509  (.A(\i53/n45 ),
    .B(\i53/n486 ),
    .Y(\i53/n501 ));
 NOR2xp33_ASAP7_75t_SL \i53/i51  (.A(\i53/n339 ),
    .B(\i53/n252 ),
    .Y(\i53/n377 ));
 NAND2xp5_ASAP7_75t_SL \i53/i510  (.A(\i53/n63 ),
    .B(\i53/n486 ),
    .Y(\i53/n502 ));
 NAND2xp5_ASAP7_75t_SL \i53/i511  (.A(\i53/n39 ),
    .B(\i53/n486 ),
    .Y(\i53/n503 ));
 NOR2x1_ASAP7_75t_L \i53/i512  (.A(\i53/n514 ),
    .B(\i53/n486 ),
    .Y(\i53/n504 ));
 NAND2xp5_ASAP7_75t_SL \i53/i513  (.A(\i53/n11 ),
    .B(n15[5]),
    .Y(\i53/n505 ));
 OAI21xp5_ASAP7_75t_SL \i53/i514  (.A1(\i53/n507 ),
    .A2(\i53/n526 ),
    .B(\i53/n95 ),
    .Y(\i53/n508 ));
 OR2x2_ASAP7_75t_SL \i53/i515  (.A(\i53/n506 ),
    .B(\i53/n505 ),
    .Y(\i53/n507 ));
 NAND2xp5_ASAP7_75t_SL \i53/i516  (.A(\i53/n0 ),
    .B(n15[6]),
    .Y(\i53/n506 ));
 NAND2xp5_ASAP7_75t_SL \i53/i517  (.A(\i53/n53 ),
    .B(\i53/n507 ),
    .Y(\i53/n509 ));
 OAI221xp5_ASAP7_75t_SL \i53/i518  (.A1(\i53/n544 ),
    .A2(\i53/n58 ),
    .B1(\i53/n425 ),
    .B2(\i53/n54 ),
    .C(\i53/n161 ),
    .Y(\i53/n510 ));
 OR2x2_ASAP7_75t_SL \i53/i519  (.A(\i53/n1 ),
    .B(n15[3]),
    .Y(\i53/n511 ));
 NAND2xp5_ASAP7_75t_SL \i53/i52  (.A(\i53/n347 ),
    .B(\i53/n342 ),
    .Y(\i53/n376 ));
 NAND2xp5_ASAP7_75t_SL \i53/i520  (.A(\i53/n2 ),
    .B(n15[1]),
    .Y(\i53/n512 ));
 INVx4_ASAP7_75t_SL \i53/i521  (.A(\i53/n513 ),
    .Y(\i53/n514 ));
 OR2x4_ASAP7_75t_SL \i53/i522  (.A(\i53/n511 ),
    .B(\i53/n512 ),
    .Y(\i53/n513 ));
 OAI221xp5_ASAP7_75t_SL \i53/i523  (.A1(\i53/n569 ),
    .A2(\i53/n416 ),
    .B1(\i53/n44 ),
    .B2(\i53/n513 ),
    .C(\i53/n490 ),
    .Y(\i53/n515 ));
 AO21x1_ASAP7_75t_SL \i53/i524  (.A1(\i53/n513 ),
    .A2(\i53/n121 ),
    .B(\i53/n110 ),
    .Y(\i53/n516 ));
 AOI31xp33_ASAP7_75t_SL \i53/i525  (.A1(\i53/n44 ),
    .A2(\i53/n62 ),
    .A3(\i53/n54 ),
    .B(\i53/n513 ),
    .Y(\i53/n517 ));
 OAI221xp5_ASAP7_75t_SL \i53/i526  (.A1(\i53/n454 ),
    .A2(\i53/n42 ),
    .B1(\i53/n38 ),
    .B2(\i53/n513 ),
    .C(\i53/n93 ),
    .Y(\i53/n518 ));
 OAI22xp33_ASAP7_75t_SL \i53/i527  (.A1(\i53/n40 ),
    .A2(\i53/n68 ),
    .B1(\i53/n513 ),
    .B2(\i53/n48 ),
    .Y(\i53/n519 ));
 OAI21xp5_ASAP7_75t_SL \i53/i528  (.A1(\i53/n58 ),
    .A2(\i53/n513 ),
    .B(\i53/n560 ),
    .Y(\i53/n520 ));
 OA21x2_ASAP7_75t_SL \i53/i529  (.A1(\i53/n44 ),
    .A2(\i53/n513 ),
    .B(\i53/n490 ),
    .Y(\i53/n521 ));
 NOR2x1_ASAP7_75t_SL \i53/i53  (.A(\i53/n256 ),
    .B(\i53/n349 ),
    .Y(\i53/n375 ));
 OAI22xp5_ASAP7_75t_SL \i53/i530  (.A1(\i53/n44 ),
    .A2(\i53/n60 ),
    .B1(\i53/n53 ),
    .B2(\i53/n513 ),
    .Y(\i53/n522 ));
 OAI22xp5_ASAP7_75t_SL \i53/i531  (.A1(\i53/n44 ),
    .A2(\i53/n42 ),
    .B1(\i53/n513 ),
    .B2(\i53/n40 ),
    .Y(\i53/n523 ));
 NOR2xp67_ASAP7_75t_L \i53/i532  (.A(\i53/n513 ),
    .B(\i53/n416 ),
    .Y(\i53/n524 ));
 NOR2xp33_ASAP7_75t_SL \i53/i533  (.A(\i53/n513 ),
    .B(\i53/n40 ),
    .Y(\i53/n525 ));
 NAND2x1p5_ASAP7_75t_SL \i53/i534  (.A(\i53/n4 ),
    .B(\i53/n555 ),
    .Y(\i53/n526 ));
 NOR2xp33_ASAP7_75t_SL \i53/i535  (.A(\i53/n470 ),
    .B(\i53/n5 ),
    .Y(\i53/n527 ));
 NAND2xp5_ASAP7_75t_SL \i53/i536  (.A(\i53/n5 ),
    .B(\i53/n448 ),
    .Y(\i53/n528 ));
 AOI22xp33_ASAP7_75t_SL \i53/i537  (.A1(\i53/n70 ),
    .A2(\i53/n514 ),
    .B1(\i53/n415 ),
    .B2(\i53/n5 ),
    .Y(\i53/n529 ));
 AOI22xp5_ASAP7_75t_SL \i53/i538  (.A1(\i53/n63 ),
    .A2(\i53/n46 ),
    .B1(\i53/n41 ),
    .B2(\i53/n5 ),
    .Y(\i53/n530 ));
 NAND2xp5_ASAP7_75t_SL \i53/i539  (.A(\i53/n72 ),
    .B(\i53/n5 ),
    .Y(\i53/n531 ));
 NOR2x1_ASAP7_75t_SL \i53/i54  (.A(\i53/n322 ),
    .B(\i53/n333 ),
    .Y(\i53/n374 ));
 NAND2xp5_ASAP7_75t_SL \i53/i540  (.A(\i53/n66 ),
    .B(\i53/n5 ),
    .Y(\i53/n532 ));
 AOI22xp5_ASAP7_75t_SL \i53/i541  (.A1(\i53/n72 ),
    .A2(\i53/n61 ),
    .B1(\i53/n59 ),
    .B2(\i53/n5 ),
    .Y(\i53/n533 ));
 AO21x2_ASAP7_75t_SL \i53/i542  (.A1(\i53/n63 ),
    .A2(\i53/n5 ),
    .B(\i53/n156 ),
    .Y(\i53/n534 ));
 NAND2xp33_ASAP7_75t_L \i53/i543  (.A(\i53/n5 ),
    .B(\i53/n59 ),
    .Y(\i53/n535 ));
 NAND2xp5_ASAP7_75t_SL \i53/i544  (.A(\i53/n39 ),
    .B(\i53/n5 ),
    .Y(\i53/n536 ));
 OAI31xp33_ASAP7_75t_SL \i53/i545  (.A1(\i53/n57 ),
    .A2(\i53/n5 ),
    .A3(\i53/n570 ),
    .B(\i53/n41 ),
    .Y(\i53/n537 ));
 AOI22xp5_ASAP7_75t_SL \i53/i546  (.A1(\i53/n46 ),
    .A2(\i53/n118 ),
    .B1(\i53/n438 ),
    .B2(\i53/n570 ),
    .Y(\i53/n538 ));
 NAND2xp5_ASAP7_75t_SL \i53/i547  (.A(\i53/n59 ),
    .B(\i53/n570 ),
    .Y(\i53/n539 ));
 AOI22xp5_ASAP7_75t_SL \i53/i548  (.A1(\i53/n72 ),
    .A2(\i53/n554 ),
    .B1(\i53/n66 ),
    .B2(\i53/n570 ),
    .Y(\i53/n540 ));
 AOI21x1_ASAP7_75t_SL \i53/i549  (.A1(\i53/n570 ),
    .A2(\i53/n49 ),
    .B(\i53/n549 ),
    .Y(\i53/n541 ));
 NAND2xp5_ASAP7_75t_SL \i53/i55  (.A(\i53/n286 ),
    .B(\i53/n327 ),
    .Y(\i53/n373 ));
 NOR2xp67_ASAP7_75t_SL \i53/i550  (.A(\i53/n44 ),
    .B(\i53/n544 ),
    .Y(\i53/n545 ));
 OR2x6_ASAP7_75t_SL \i53/i551  (.A(\i53/n542 ),
    .B(\i53/n543 ),
    .Y(\i53/n544 ));
 INVx1_ASAP7_75t_SL \i53/i552  (.A(\i53/n555 ),
    .Y(\i53/n542 ));
 INVx2_ASAP7_75t_SL \i53/i553  (.A(\i53/n35 ),
    .Y(\i53/n543 ));
 OAI22x1_ASAP7_75t_SL \i53/i554  (.A1(\i53/n416 ),
    .A2(\i53/n60 ),
    .B1(\i53/n54 ),
    .B2(\i53/n544 ),
    .Y(\i53/n546 ));
 OAI22xp5_ASAP7_75t_SL \i53/i555  (.A1(\i53/n69 ),
    .A2(\i53/n526 ),
    .B1(\i53/n507 ),
    .B2(\i53/n544 ),
    .Y(\i53/n547 ));
 OAI22xp33_ASAP7_75t_SL \i53/i556  (.A1(\i53/n48 ),
    .A2(\i53/n37 ),
    .B1(\i53/n544 ),
    .B2(\i53/n50 ),
    .Y(\i53/n548 ));
 OAI22xp5_ASAP7_75t_SL \i53/i557  (.A1(\i53/n48 ),
    .A2(\i53/n544 ),
    .B1(\i53/n71 ),
    .B2(\i53/n8 ),
    .Y(\i53/n549 ));
 OAI221xp5_ASAP7_75t_SL \i53/i558  (.A1(\i53/n544 ),
    .A2(\i53/n62 ),
    .B1(\i53/n14 ),
    .B2(\i53/n444 ),
    .C(\i53/n184 ),
    .Y(\i53/n550 ));
 OAI222xp33_ASAP7_75t_SL \i53/i559  (.A1(\i53/n544 ),
    .A2(\i53/n38 ),
    .B1(\i53/n42 ),
    .B2(\i53/n444 ),
    .C1(\i53/n56 ),
    .C2(\i53/n53 ),
    .Y(\i53/n551 ));
 NOR5xp2_ASAP7_75t_SL \i53/i56  (.A(\i53/n219 ),
    .B(\i53/n515 ),
    .C(\i53/n230 ),
    .D(\i53/n22 ),
    .E(\i53/n510 ),
    .Y(\i53/n372 ));
 AOI21xp5_ASAP7_75t_L \i53/i560  (.A1(\i53/n50 ),
    .A2(\i53/n130 ),
    .B(\i53/n544 ),
    .Y(\i53/n552 ));
 A2O1A1Ixp33_ASAP7_75t_R \i53/i561  (.A1(\i53/n544 ),
    .A2(\i53/n42 ),
    .B(\i53/n54 ),
    .C(\i53/n90 ),
    .Y(\i53/n553 ));
 INVx4_ASAP7_75t_SL \i53/i562  (.A(\i53/n544 ),
    .Y(\i53/n554 ));
 AND2x4_ASAP7_75t_SL \i53/i563  (.A(n15[0]),
    .B(\i53/n25 ),
    .Y(\i53/n555 ));
 NAND2xp5_ASAP7_75t_SL \i53/i564  (.A(\i53/n556 ),
    .B(\i53/n438 ),
    .Y(\i53/n557 ));
 AND2x4_ASAP7_75t_SL \i53/i565  (.A(\i53/n555 ),
    .B(\i53/n6 ),
    .Y(\i53/n556 ));
 NOR2xp33_ASAP7_75t_SL \i53/i566  (.A(\i53/n423 ),
    .B(\i53/n556 ),
    .Y(\i53/n558 ));
 AOI22xp5_ASAP7_75t_R \i53/i567  (.A1(\i53/n415 ),
    .A2(\i53/n46 ),
    .B1(\i53/n72 ),
    .B2(\i53/n556 ),
    .Y(\i53/n559 ));
 NAND2xp5_ASAP7_75t_SL \i53/i568  (.A(\i53/n45 ),
    .B(\i53/n556 ),
    .Y(\i53/n560 ));
 NAND2xp5_ASAP7_75t_SL \i53/i569  (.A(\i53/n63 ),
    .B(\i53/n556 ),
    .Y(\i53/n561 ));
 NOR2x1_ASAP7_75t_SL \i53/i57  (.A(\i53/n3 ),
    .B(\i53/n334 ),
    .Y(\i53/n371 ));
 NAND2xp5_ASAP7_75t_SL \i53/i570  (.A(\i53/n7 ),
    .B(\i53/n556 ),
    .Y(\i53/n562 ));
 NAND2xp5_ASAP7_75t_SL \i53/i571  (.A(\i53/n51 ),
    .B(\i53/n556 ),
    .Y(\i53/n563 ));
 NAND2xp5_ASAP7_75t_SL \i53/i572  (.A(\i53/n556 ),
    .B(\i53/n49 ),
    .Y(\i53/n564 ));
 OAI21xp5_ASAP7_75t_SL \i53/i573  (.A1(\i53/n556 ),
    .A2(\i53/n61 ),
    .B(\i53/n59 ),
    .Y(\i53/n565 ));
 AOI22xp33_ASAP7_75t_SL \i53/i574  (.A1(\i53/n49 ),
    .A2(\i53/n46 ),
    .B1(\i53/n59 ),
    .B2(\i53/n556 ),
    .Y(\i53/n566 ));
 AOI22xp5_ASAP7_75t_SL \i53/i575  (.A1(\i53/n66 ),
    .A2(\i53/n556 ),
    .B1(\i53/n59 ),
    .B2(\i53/n57 ),
    .Y(\i53/n567 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i53/i576  (.A1(\i53/n46 ),
    .A2(\i53/n556 ),
    .B(\i53/n7 ),
    .C(\i53/n131 ),
    .Y(\i53/n568 ));
 INVx4_ASAP7_75t_SL \i53/i577  (.A(\i53/n556 ),
    .Y(\i53/n569 ));
 AND2x4_ASAP7_75t_SL \i53/i578  (.A(\i53/n422 ),
    .B(\i53/n6 ),
    .Y(\i53/n570 ));
 NAND4xp25_ASAP7_75t_SL \i53/i579  (.A(\i53/n157 ),
    .B(\i53/n168 ),
    .C(\i53/n238 ),
    .D(\i53/n571 ),
    .Y(\i53/n572 ));
 NAND2x1_ASAP7_75t_SL \i53/i58  (.A(\i53/n331 ),
    .B(\i53/n312 ),
    .Y(\i53/n384 ));
 NAND2x1_ASAP7_75t_SL \i53/i580  (.A(\i53/n7 ),
    .B(\i53/n570 ),
    .Y(\i53/n571 ));
 INVx1_ASAP7_75t_SL \i53/i581  (.A(\i53/n571 ),
    .Y(\i53/n573 ));
 NAND2xp5_ASAP7_75t_L \i53/i582  (.A(\i53/n571 ),
    .B(\i53/n119 ),
    .Y(\i53/n574 ));
 NOR3xp33_ASAP7_75t_SL \i53/i583  (.A(\i53/n575 ),
    .B(\i53/n111 ),
    .C(\i53/n113 ),
    .Y(\i53/n576 ));
 AO21x1_ASAP7_75t_SL \i53/i584  (.A1(\i53/n70 ),
    .A2(\i53/n57 ),
    .B(\i53/n241 ),
    .Y(\i53/n575 ));
 NAND2xp5_ASAP7_75t_SL \i53/i585  (.A(\i53/n70 ),
    .B(\i53/n57 ),
    .Y(\i53/n577 ));
 AND4x1_ASAP7_75t_SL \i53/i586  (.A(\i53/n459 ),
    .B(\i53/n254 ),
    .C(\i53/n265 ),
    .D(\i53/n200 ),
    .Y(\i53/n578 ));
 AND2x2_ASAP7_75t_SL \i53/i587  (.A(\i53/n579 ),
    .B(\i53/n346 ),
    .Y(\i53/n580 ));
 AOI21xp33_ASAP7_75t_SL \i53/i588  (.A1(\i53/n36 ),
    .A2(\i53/n55 ),
    .B(\i53/n89 ),
    .Y(\i53/n579 ));
 NAND3xp33_ASAP7_75t_SL \i53/i589  (.A(\i53/n581 ),
    .B(\i53/n418 ),
    .C(\i53/n246 ),
    .Y(\i53/n582 ));
 NOR2x1_ASAP7_75t_SL \i53/i59  (.A(\i53/n350 ),
    .B(\i53/n333 ),
    .Y(\i53/n370 ));
 AO21x1_ASAP7_75t_SL \i53/i590  (.A1(\i53/n416 ),
    .A2(\i53/n44 ),
    .B(\i53/n473 ),
    .Y(\i53/n581 ));
 NOR3xp33_ASAP7_75t_SL \i53/i591  (.A(\i53/n583 ),
    .B(\i53/n244 ),
    .C(\i53/n156 ),
    .Y(\i53/n584 ));
 OAI21xp5_ASAP7_75t_SL \i53/i592  (.A1(\i53/n53 ),
    .A2(\i53/n14 ),
    .B(\i53/n528 ),
    .Y(\i53/n583 ));
 INVx1_ASAP7_75t_SL \i53/i6  (.A(\i53/n29 ),
    .Y(\i53/n6 ));
 NOR2x1_ASAP7_75t_SL \i53/i60  (.A(\i53/n270 ),
    .B(\i53/n332 ),
    .Y(\i53/n383 ));
 INVxp67_ASAP7_75t_SL \i53/i61  (.A(\i53/n368 ),
    .Y(\i53/n369 ));
 INVxp67_ASAP7_75t_SL \i53/i62  (.A(\i53/n364 ),
    .Y(\i53/n365 ));
 AND5x1_ASAP7_75t_SL \i53/i63  (.A(\i53/n283 ),
    .B(\i53/n265 ),
    .C(\i53/n463 ),
    .D(\i53/n568 ),
    .E(\i53/n499 ),
    .Y(\i53/n363 ));
 NOR3xp33_ASAP7_75t_SL \i53/i64  (.A(\i53/n293 ),
    .B(\i53/n275 ),
    .C(\i53/n257 ),
    .Y(\i53/n362 ));
 NOR3xp33_ASAP7_75t_SL \i53/i65  (.A(\i53/n572 ),
    .B(\i53/n258 ),
    .C(\i53/n218 ),
    .Y(\i53/n361 ));
 AND5x1_ASAP7_75t_SL \i53/i66  (.A(\i53/n248 ),
    .B(\i53/n261 ),
    .C(\i53/n242 ),
    .D(\i53/n251 ),
    .E(\i53/n196 ),
    .Y(\i53/n360 ));
 NOR2xp33_ASAP7_75t_SL \i53/i67  (.A(\i53/n320 ),
    .B(\i53/n325 ),
    .Y(\i53/n359 ));
 NAND4xp25_ASAP7_75t_SL \i53/i68  (.A(\i53/n303 ),
    .B(\i53/n311 ),
    .C(\i53/n316 ),
    .D(\i53/n299 ),
    .Y(\i53/n358 ));
 NAND5xp2_ASAP7_75t_SL \i53/i69  (.A(\i53/n282 ),
    .B(\i53/n240 ),
    .C(\i53/n171 ),
    .D(\i53/n159 ),
    .E(\i53/n226 ),
    .Y(\i53/n357 ));
 INVx2_ASAP7_75t_SL \i53/i7  (.A(\i53/n507 ),
    .Y(\i53/n7 ));
 NOR4xp25_ASAP7_75t_SL \i53/i70  (.A(\i53/n273 ),
    .B(\i53/n515 ),
    .C(\i53/n231 ),
    .D(\i53/n212 ),
    .Y(\i53/n356 ));
 NAND4xp25_ASAP7_75t_SL \i53/i71  (.A(\i53/n305 ),
    .B(\i53/n289 ),
    .C(\i53/n308 ),
    .D(\i53/n310 ),
    .Y(\i53/n355 ));
 NAND4xp25_ASAP7_75t_SL \i53/i72  (.A(\i53/n318 ),
    .B(\i53/n316 ),
    .C(\i53/n521 ),
    .D(\i53/n190 ),
    .Y(\i53/n354 ));
 NAND3xp33_ASAP7_75t_SL \i53/i73  (.A(\i53/n310 ),
    .B(\i53/n281 ),
    .C(\i53/n15 ),
    .Y(\i53/n368 ));
 NAND4xp75_ASAP7_75t_SL \i53/i74  (.A(\i53/n417 ),
    .B(\i53/n203 ),
    .C(\i53/n269 ),
    .D(\i53/n19 ),
    .Y(\i53/n367 ));
 NAND2xp33_ASAP7_75t_L \i53/i75  (.A(\i53/n288 ),
    .B(\i53/n351 ),
    .Y(\i53/n353 ));
 AND2x2_ASAP7_75t_SL \i53/i76  (.A(\i53/n291 ),
    .B(\i53/n340 ),
    .Y(\i53/n366 ));
 NAND2x1p5_ASAP7_75t_SL \i53/i77  (.A(\i53/n348 ),
    .B(\i53/n304 ),
    .Y(\i53/n364 ));
 INVxp67_ASAP7_75t_SL \i53/i78  (.A(\i53/n351 ),
    .Y(\i53/n352 ));
 NOR5xp2_ASAP7_75t_SL \i53/i79  (.A(\i53/n552 ),
    .B(\i53/n217 ),
    .C(\i53/n165 ),
    .D(\i53/n140 ),
    .E(\i53/n525 ),
    .Y(\i53/n343 ));
 INVx2_ASAP7_75t_SL \i53/i8  (.A(\i53/n570 ),
    .Y(\i53/n8 ));
 NOR3xp33_ASAP7_75t_SL \i53/i80  (.A(\i53/n315 ),
    .B(\i53/n234 ),
    .C(\i53/n229 ),
    .Y(\i53/n342 ));
 NOR2xp33_ASAP7_75t_SL \i53/i81  (.A(\i53/n272 ),
    .B(\i53/n290 ),
    .Y(\i53/n341 ));
 NOR2xp33_ASAP7_75t_SL \i53/i82  (.A(\i53/n313 ),
    .B(\i53/n263 ),
    .Y(\i53/n340 ));
 NOR2x1_ASAP7_75t_SL \i53/i83  (.A(\i53/n276 ),
    .B(\i53/n249 ),
    .Y(\i53/n351 ));
 NAND3xp33_ASAP7_75t_SL \i53/i84  (.A(\i53/n225 ),
    .B(\i53/n537 ),
    .C(\i53/n472 ),
    .Y(\i53/n339 ));
 NAND2xp5_ASAP7_75t_L \i53/i85  (.A(\i53/n312 ),
    .B(\i53/n280 ),
    .Y(\i53/n338 ));
 NAND2xp5_ASAP7_75t_SL \i53/i86  (.A(\i53/n262 ),
    .B(\i53/n302 ),
    .Y(\i53/n337 ));
 NAND3xp33_ASAP7_75t_SL \i53/i87  (.A(\i53/n265 ),
    .B(\i53/n214 ),
    .C(\i53/n200 ),
    .Y(\i53/n350 ));
 NOR3xp33_ASAP7_75t_SL \i53/i88  (.A(\i53/n434 ),
    .B(\i53/n10 ),
    .C(\i53/n550 ),
    .Y(\i53/n336 ));
 NAND2xp5_ASAP7_75t_SL \i53/i89  (.A(\i53/n17 ),
    .B(\i53/n289 ),
    .Y(\i53/n349 ));
 NOR2x1p5_ASAP7_75t_SL \i53/i9  (.A(\i53/n409 ),
    .B(\i53/n408 ),
    .Y(n14[4]));
 OR3x1_ASAP7_75t_SL \i53/i90  (.A(\i53/n219 ),
    .B(\i53/n230 ),
    .C(\i53/n22 ),
    .Y(\i53/n335 ));
 NOR2x1_ASAP7_75t_SL \i53/i91  (.A(\i53/n229 ),
    .B(\i53/n315 ),
    .Y(\i53/n348 ));
 NOR2xp33_ASAP7_75t_L \i53/i92  (.A(\i53/n274 ),
    .B(\i53/n260 ),
    .Y(\i53/n347 ));
 NOR2xp33_ASAP7_75t_SL \i53/i93  (.A(\i53/n220 ),
    .B(\i53/n301 ),
    .Y(\i53/n346 ));
 NOR3x1_ASAP7_75t_SL \i53/i94  (.A(\i53/n224 ),
    .B(\i53/n149 ),
    .C(\i53/n266 ),
    .Y(\i53/n345 ));
 NOR2xp33_ASAP7_75t_SL \i53/i95  (.A(\i53/n298 ),
    .B(\i53/n292 ),
    .Y(\i53/n344 ));
 NOR3xp33_ASAP7_75t_SL \i53/i96  (.A(\i53/n232 ),
    .B(\i53/n170 ),
    .C(\i53/n223 ),
    .Y(\i53/n331 ));
 NOR2xp33_ASAP7_75t_SL \i53/i97  (.A(\i53/n285 ),
    .B(\i53/n582 ),
    .Y(\i53/n330 ));
 NAND3xp33_ASAP7_75t_SL \i53/i98  (.A(\i53/n459 ),
    .B(\i53/n278 ),
    .C(\i53/n477 ),
    .Y(\i53/n329 ));
 NAND4xp25_ASAP7_75t_SL \i53/i99  (.A(\i53/n207 ),
    .B(\i53/n474 ),
    .C(\i53/n489 ),
    .D(\i53/n213 ),
    .Y(\i53/n328 ));
 AOI22xp5_ASAP7_75t_SL i530 (.A1(n547),
    .A2(n1155),
    .B1(n546),
    .B2(n226),
    .Y(n942));
 XNOR2xp5_ASAP7_75t_SL i531 (.A(n591),
    .B(n494),
    .Y(n941));
 AOI22xp5_ASAP7_75t_SL i532 (.A1(n520),
    .A2(n794),
    .B1(n519),
    .B2(n793),
    .Y(n940));
 XNOR2xp5_ASAP7_75t_SL i533 (.A(n602),
    .B(n332),
    .Y(n939));
 OAI22xp5_ASAP7_75t_SL i534 (.A1(n218),
    .A2(n1163),
    .B1(n550),
    .B2(n476),
    .Y(n938));
 XOR2xp5_ASAP7_75t_SL i535 (.A(n335),
    .B(n333),
    .Y(n937));
 AOI22xp5_ASAP7_75t_SL i536 (.A1(n551),
    .A2(n812),
    .B1(n813),
    .B2(n552),
    .Y(n936));
 XOR2xp5_ASAP7_75t_SL i537 (.A(n338),
    .B(n339),
    .Y(n935));
 OAI22xp5_ASAP7_75t_SL i538 (.A1(n560),
    .A2(n1175),
    .B1(n559),
    .B2(n792),
    .Y(n934));
 OAI22xp5_ASAP7_75t_SL i539 (.A1(n566),
    .A2(n808),
    .B1(n565),
    .B2(n807),
    .Y(n933));
 INVx2_ASAP7_75t_SL \i54/i0  (.A(n13[2]),
    .Y(\i54/n0 ));
 INVx2_ASAP7_75t_SL \i54/i1  (.A(n13[0]),
    .Y(\i54/n1 ));
 AND3x4_ASAP7_75t_SL \i54/i10  (.A(\i54/n490 ),
    .B(\i54/n499 ),
    .C(\i54/n478 ),
    .Y(n12[1]));
 NAND2xp33_ASAP7_75t_SL \i54/i100  (.A(\i54/n295 ),
    .B(\i54/n394 ),
    .Y(\i54/n414 ));
 NOR5xp2_ASAP7_75t_SL \i54/i101  (.A(\i54/n338 ),
    .B(\i54/n303 ),
    .C(\i54/n324 ),
    .D(\i54/n271 ),
    .E(\i54/n552 ),
    .Y(\i54/n413 ));
 NAND5xp2_ASAP7_75t_SL \i54/i102  (.A(\i54/n281 ),
    .B(\i54/n530 ),
    .C(\i54/n507 ),
    .D(\i54/n322 ),
    .E(\i54/n267 ),
    .Y(\i54/n412 ));
 NAND3xp33_ASAP7_75t_L \i54/i103  (.A(\i54/n276 ),
    .B(\i54/n308 ),
    .C(\i54/n377 ),
    .Y(\i54/n411 ));
 NOR5xp2_ASAP7_75t_SL \i54/i104  (.A(\i54/n274 ),
    .B(\i54/n121 ),
    .C(\i54/n265 ),
    .D(\i54/n287 ),
    .E(\i54/n100 ),
    .Y(\i54/n410 ));
 NAND5xp2_ASAP7_75t_SL \i54/i105  (.A(\i54/n24 ),
    .B(\i54/n352 ),
    .C(\i54/n507 ),
    .D(\i54/n97 ),
    .E(\i54/n191 ),
    .Y(\i54/n409 ));
 NAND4xp25_ASAP7_75t_SL \i54/i106  (.A(\i54/n214 ),
    .B(\i54/n227 ),
    .C(\i54/n328 ),
    .D(\i54/n16 ),
    .Y(\i54/n408 ));
 NOR5xp2_ASAP7_75t_SL \i54/i107  (.A(\i54/n233 ),
    .B(\i54/n545 ),
    .C(\i54/n219 ),
    .D(\i54/n185 ),
    .E(\i54/n183 ),
    .Y(\i54/n407 ));
 NOR2xp33_ASAP7_75t_SL \i54/i108  (.A(\i54/n368 ),
    .B(\i54/n401 ),
    .Y(\i54/n406 ));
 NOR2xp33_ASAP7_75t_SL \i54/i109  (.A(\i54/n356 ),
    .B(\i54/n386 ),
    .Y(\i54/n405 ));
 NOR2x1p5_ASAP7_75t_SL \i54/i11  (.A(\i54/n500 ),
    .B(\i54/n491 ),
    .Y(n12[5]));
 NAND3x1_ASAP7_75t_SL \i54/i110  (.A(\i54/n231 ),
    .B(\i54/n384 ),
    .C(\i54/n530 ),
    .Y(\i54/n422 ));
 NAND3x1_ASAP7_75t_SL \i54/i111  (.A(\i54/n347 ),
    .B(\i54/n329 ),
    .C(\i54/n296 ),
    .Y(\i54/n421 ));
 AOI21xp5_ASAP7_75t_L \i54/i112  (.A1(\i54/n71 ),
    .A2(\i54/n236 ),
    .B(\i54/n163 ),
    .Y(\i54/n397 ));
 NOR2xp33_ASAP7_75t_SL \i54/i113  (.A(\i54/n338 ),
    .B(\i54/n301 ),
    .Y(\i54/n396 ));
 NAND2xp5_ASAP7_75t_SL \i54/i114  (.A(\i54/n327 ),
    .B(\i54/n355 ),
    .Y(\i54/n395 ));
 NOR2xp33_ASAP7_75t_SL \i54/i115  (.A(\i54/n354 ),
    .B(\i54/n25 ),
    .Y(\i54/n394 ));
 NOR2xp33_ASAP7_75t_SL \i54/i116  (.A(\i54/n333 ),
    .B(\i54/n343 ),
    .Y(\i54/n393 ));
 NOR2xp67_ASAP7_75t_SL \i54/i117  (.A(\i54/n173 ),
    .B(\i54/n340 ),
    .Y(\i54/n392 ));
 NOR2xp33_ASAP7_75t_SL \i54/i118  (.A(\i54/n338 ),
    .B(\i54/n20 ),
    .Y(\i54/n391 ));
 NOR4xp25_ASAP7_75t_SL \i54/i119  (.A(\i54/n312 ),
    .B(\i54/n20 ),
    .C(\i54/n22 ),
    .D(\i54/n180 ),
    .Y(\i54/n390 ));
 AND2x4_ASAP7_75t_SL \i54/i12  (.A(\i54/n501 ),
    .B(\i54/n484 ),
    .Y(n12[0]));
 NAND2xp67_ASAP7_75t_SL \i54/i120  (.A(\i54/n261 ),
    .B(\i54/n319 ),
    .Y(\i54/n389 ));
 NOR4xp25_ASAP7_75t_SL \i54/i121  (.A(\i54/n117 ),
    .B(\i54/n253 ),
    .C(\i54/n221 ),
    .D(\i54/n237 ),
    .Y(\i54/n388 ));
 NOR3xp33_ASAP7_75t_SL \i54/i122  (.A(\i54/n258 ),
    .B(\i54/n540 ),
    .C(\i54/n257 ),
    .Y(\i54/n387 ));
 NAND2xp33_ASAP7_75t_SL \i54/i123  (.A(\i54/n307 ),
    .B(\i54/n21 ),
    .Y(\i54/n386 ));
 NOR2xp33_ASAP7_75t_SL \i54/i124  (.A(\i54/n301 ),
    .B(\i54/n302 ),
    .Y(\i54/n385 ));
 NOR2x1_ASAP7_75t_SL \i54/i125  (.A(\i54/n282 ),
    .B(\i54/n569 ),
    .Y(\i54/n384 ));
 NAND2xp33_ASAP7_75t_SL \i54/i126  (.A(\i54/n353 ),
    .B(\i54/n336 ),
    .Y(\i54/n383 ));
 NAND3xp33_ASAP7_75t_SL \i54/i127  (.A(\i54/n23 ),
    .B(\i54/n212 ),
    .C(\i54/n571 ),
    .Y(\i54/n382 ));
 NOR3xp33_ASAP7_75t_SL \i54/i128  (.A(\i54/n215 ),
    .B(\i54/n228 ),
    .C(\i54/n198 ),
    .Y(\i54/n404 ));
 NAND2xp5_ASAP7_75t_SL \i54/i129  (.A(\i54/n311 ),
    .B(\i54/n214 ),
    .Y(\i54/n403 ));
 NOR3xp33_ASAP7_75t_SL \i54/i13  (.A(\i54/n473 ),
    .B(\i54/n469 ),
    .C(\i54/n476 ),
    .Y(\i54/n501 ));
 NOR2x1_ASAP7_75t_SL \i54/i130  (.A(\i54/n546 ),
    .B(\i54/n305 ),
    .Y(\i54/n402 ));
 NAND2xp5_ASAP7_75t_SL \i54/i131  (.A(\i54/n507 ),
    .B(\i54/n313 ),
    .Y(\i54/n401 ));
 NOR2x1_ASAP7_75t_SL \i54/i132  (.A(\i54/n283 ),
    .B(\i54/n341 ),
    .Y(\i54/n400 ));
 NOR2x1_ASAP7_75t_SL \i54/i133  (.A(\i54/n22 ),
    .B(\i54/n301 ),
    .Y(\i54/n399 ));
 NOR3x1_ASAP7_75t_SL \i54/i134  (.A(\i54/n219 ),
    .B(\i54/n524 ),
    .C(\i54/n182 ),
    .Y(\i54/n398 ));
 INVx1_ASAP7_75t_SL \i54/i135  (.A(\i54/n379 ),
    .Y(\i54/n380 ));
 INVx1_ASAP7_75t_SL \i54/i136  (.A(\i54/n26 ),
    .Y(\i54/n378 ));
 NOR4xp25_ASAP7_75t_SL \i54/i137  (.A(\i54/n201 ),
    .B(\i54/n239 ),
    .C(\i54/n226 ),
    .D(\i54/n195 ),
    .Y(\i54/n377 ));
 AOI211xp5_ASAP7_75t_SL \i54/i138  (.A1(\i54/n70 ),
    .A2(\i54/n65 ),
    .B(\i54/n569 ),
    .C(\i54/n559 ),
    .Y(\i54/n376 ));
 NAND2xp33_ASAP7_75t_SL \i54/i139  (.A(\i54/n297 ),
    .B(\i54/n321 ),
    .Y(\i54/n375 ));
 NOR2x1p5_ASAP7_75t_SL \i54/i14  (.A(\i54/n493 ),
    .B(\i54/n494 ),
    .Y(n12[2]));
 NAND5xp2_ASAP7_75t_SL \i54/i140  (.A(\i54/n534 ),
    .B(\i54/n251 ),
    .C(\i54/n263 ),
    .D(\i54/n509 ),
    .E(\i54/n118 ),
    .Y(\i54/n374 ));
 NOR4xp25_ASAP7_75t_SL \i54/i141  (.A(\i54/n549 ),
    .B(\i54/n152 ),
    .C(\i54/n153 ),
    .D(\i54/n169 ),
    .Y(\i54/n373 ));
 NOR2xp33_ASAP7_75t_SL \i54/i142  (.A(\i54/n288 ),
    .B(\i54/n292 ),
    .Y(\i54/n372 ));
 AOI211xp5_ASAP7_75t_SL \i54/i143  (.A1(\i54/n72 ),
    .A2(\i54/n167 ),
    .B(\i54/n273 ),
    .C(\i54/n187 ),
    .Y(\i54/n371 ));
 OA21x2_ASAP7_75t_SL \i54/i144  (.A1(\i54/n58 ),
    .A2(\i54/n71 ),
    .B(\i54/n352 ),
    .Y(\i54/n370 ));
 NOR4xp25_ASAP7_75t_SL \i54/i145  (.A(\i54/n266 ),
    .B(\i54/n177 ),
    .C(\i54/n207 ),
    .D(\i54/n182 ),
    .Y(\i54/n369 ));
 NAND5xp2_ASAP7_75t_SL \i54/i146  (.A(\i54/n537 ),
    .B(\i54/n106 ),
    .C(\i54/n158 ),
    .D(\i54/n154 ),
    .E(\i54/n98 ),
    .Y(\i54/n368 ));
 NOR3xp33_ASAP7_75t_SL \i54/i147  (.A(\i54/n306 ),
    .B(\i54/n178 ),
    .C(\i54/n96 ),
    .Y(\i54/n367 ));
 NAND2xp5_ASAP7_75t_SL \i54/i148  (.A(\i54/n286 ),
    .B(\i54/n24 ),
    .Y(\i54/n366 ));
 NAND5xp2_ASAP7_75t_SL \i54/i149  (.A(\i54/n210 ),
    .B(\i54/n111 ),
    .C(\i54/n205 ),
    .D(\i54/n194 ),
    .E(\i54/n193 ),
    .Y(\i54/n365 ));
 NAND4xp75_ASAP7_75t_SL \i54/i15  (.A(\i54/n459 ),
    .B(\i54/n479 ),
    .C(\i54/n457 ),
    .D(\i54/n573 ),
    .Y(\i54/n500 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i54/i150  (.A1(\i54/n76 ),
    .A2(\i54/n101 ),
    .B(\i54/n78 ),
    .C(\i54/n278 ),
    .Y(\i54/n364 ));
 NAND4xp25_ASAP7_75t_SL \i54/i151  (.A(\i54/n531 ),
    .B(\i54/n252 ),
    .C(\i54/n119 ),
    .D(\i54/n179 ),
    .Y(\i54/n363 ));
 NAND5xp2_ASAP7_75t_SL \i54/i152  (.A(\i54/n168 ),
    .B(\i54/n561 ),
    .C(\i54/n243 ),
    .D(\i54/n114 ),
    .E(\i54/n109 ),
    .Y(\i54/n362 ));
 NAND2xp5_ASAP7_75t_SL \i54/i153  (.A(\i54/n285 ),
    .B(\i54/n310 ),
    .Y(\i54/n361 ));
 NAND3xp33_ASAP7_75t_SL \i54/i154  (.A(\i54/n304 ),
    .B(\i54/n572 ),
    .C(\i54/n103 ),
    .Y(\i54/n360 ));
 NAND2xp5_ASAP7_75t_SL \i54/i155  (.A(\i54/n530 ),
    .B(\i54/n231 ),
    .Y(\i54/n359 ));
 NOR2xp33_ASAP7_75t_L \i54/i156  (.A(\i54/n332 ),
    .B(\i54/n343 ),
    .Y(\i54/n381 ));
 NAND2xp5_ASAP7_75t_SL \i54/i157  (.A(\i54/n232 ),
    .B(\i54/n353 ),
    .Y(\i54/n358 ));
 NOR2x1p5_ASAP7_75t_SL \i54/i158  (.A(\i54/n290 ),
    .B(\i54/n335 ),
    .Y(\i54/n379 ));
 NAND3x1_ASAP7_75t_SL \i54/i159  (.A(\i54/n270 ),
    .B(\i54/n147 ),
    .C(\i54/n155 ),
    .Y(\i54/n26 ));
 NOR3xp33_ASAP7_75t_SL \i54/i16  (.A(\i54/n487 ),
    .B(\i54/n442 ),
    .C(\i54/n477 ),
    .Y(\i54/n499 ));
 INVxp67_ASAP7_75t_SL \i54/i160  (.A(\i54/n356 ),
    .Y(\i54/n357 ));
 INVxp67_ASAP7_75t_SL \i54/i161  (.A(\i54/n8 ),
    .Y(\i54/n355 ));
 INVxp67_ASAP7_75t_SL \i54/i162  (.A(\i54/n350 ),
    .Y(\i54/n351 ));
 INVxp67_ASAP7_75t_SL \i54/i163  (.A(\i54/n348 ),
    .Y(\i54/n349 ));
 INVx2_ASAP7_75t_SL \i54/i164  (.A(\i54/n346 ),
    .Y(\i54/n347 ));
 INVxp67_ASAP7_75t_SL \i54/i165  (.A(\i54/n506 ),
    .Y(\i54/n345 ));
 INVxp67_ASAP7_75t_SL \i54/i166  (.A(\i54/n341 ),
    .Y(\i54/n342 ));
 INVxp67_ASAP7_75t_SL \i54/i167  (.A(\i54/n547 ),
    .Y(\i54/n339 ));
 INVx1_ASAP7_75t_SL \i54/i168  (.A(\i54/n336 ),
    .Y(\i54/n337 ));
 NAND2x1_ASAP7_75t_SL \i54/i169  (.A(\i54/n225 ),
    .B(\i54/n223 ),
    .Y(\i54/n335 ));
 NAND4xp75_ASAP7_75t_SL \i54/i17  (.A(\i54/n489 ),
    .B(\i54/n458 ),
    .C(\i54/n463 ),
    .D(\i54/n453 ),
    .Y(\i54/n498 ));
 NOR2xp33_ASAP7_75t_SL \i54/i170  (.A(\i54/n264 ),
    .B(\i54/n258 ),
    .Y(\i54/n334 ));
 NAND2xp33_ASAP7_75t_SL \i54/i171  (.A(\i54/n212 ),
    .B(\i54/n507 ),
    .Y(\i54/n333 ));
 NAND2xp5_ASAP7_75t_SL \i54/i172  (.A(\i54/n181 ),
    .B(\i54/n212 ),
    .Y(\i54/n332 ));
 AOI211xp5_ASAP7_75t_SL \i54/i173  (.A1(\i54/n90 ),
    .A2(\i54/n31 ),
    .B(\i54/n125 ),
    .C(\i54/n132 ),
    .Y(\i54/n331 ));
 NOR3xp33_ASAP7_75t_SL \i54/i174  (.A(\i54/n540 ),
    .B(\i54/n144 ),
    .C(\i54/n130 ),
    .Y(\i54/n330 ));
 NOR3xp33_ASAP7_75t_SL \i54/i175  (.A(\i54/n123 ),
    .B(\i54/n138 ),
    .C(\i54/n264 ),
    .Y(\i54/n329 ));
 OAI31xp33_ASAP7_75t_SL \i54/i176  (.A1(\i54/n48 ),
    .A2(\i54/n50 ),
    .A3(\i54/n68 ),
    .B(\i54/n90 ),
    .Y(\i54/n328 ));
 AOI221xp5_ASAP7_75t_SL \i54/i177  (.A1(\i54/n76 ),
    .A2(\i54/n93 ),
    .B1(\i54/n54 ),
    .B2(\i54/n62 ),
    .C(\i54/n196 ),
    .Y(\i54/n327 ));
 OAI31xp33_ASAP7_75t_SL \i54/i178  (.A1(\i54/n72 ),
    .A2(\i54/n74 ),
    .A3(\i54/n76 ),
    .B(\i54/n68 ),
    .Y(\i54/n326 ));
 AOI21xp5_ASAP7_75t_SL \i54/i179  (.A1(\i54/n163 ),
    .A2(\i54/n503 ),
    .B(\i54/n88 ),
    .Y(\i54/n356 ));
 AND3x4_ASAP7_75t_SL \i54/i18  (.A(\i54/n480 ),
    .B(\i54/n495 ),
    .C(\i54/n485 ),
    .Y(n12[7]));
 AOI21xp5_ASAP7_75t_L \i54/i180  (.A1(\i54/n503 ),
    .A2(\i54/n174 ),
    .B(\i54/n87 ),
    .Y(\i54/n325 ));
 OAI221xp5_ASAP7_75t_SL \i54/i181  (.A1(\i54/n15 ),
    .A2(\i54/n92 ),
    .B1(\i54/n49 ),
    .B2(\i54/n56 ),
    .C(\i54/n220 ),
    .Y(\i54/n324 ));
 AOI21xp33_ASAP7_75t_SL \i54/i182  (.A1(\i54/n174 ),
    .A2(\i54/n47 ),
    .B(\i54/n75 ),
    .Y(\i54/n323 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i54/i183  (.A1(\i54/n85 ),
    .A2(\i54/n5 ),
    .B(\i54/n89 ),
    .C(\i54/n17 ),
    .Y(\i54/n322 ));
 NOR3xp33_ASAP7_75t_SL \i54/i184  (.A(\i54/n234 ),
    .B(\i54/n123 ),
    .C(\i54/n151 ),
    .Y(\i54/n321 ));
 NAND3xp33_ASAP7_75t_SL \i54/i185  (.A(\i54/n18 ),
    .B(\i54/n511 ),
    .C(\i54/n172 ),
    .Y(\i54/n320 ));
 AOI22xp5_ASAP7_75t_SL \i54/i186  (.A1(\i54/n60 ),
    .A2(\i54/n159 ),
    .B1(\i54/n62 ),
    .B2(\i54/n53 ),
    .Y(\i54/n319 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i54/i187  (.A1(\i54/n87 ),
    .A2(\i54/n51 ),
    .B(\i54/n67 ),
    .C(\i54/n126 ),
    .Y(\i54/n318 ));
 NAND4xp25_ASAP7_75t_SL \i54/i188  (.A(\i54/n184 ),
    .B(\i54/n179 ),
    .C(\i54/n555 ),
    .D(\i54/n156 ),
    .Y(\i54/n317 ));
 NAND2xp33_ASAP7_75t_SL \i54/i189  (.A(\i54/n246 ),
    .B(\i54/n150 ),
    .Y(\i54/n316 ));
 NAND4xp75_ASAP7_75t_SL \i54/i19  (.A(\i54/n577 ),
    .B(\i54/n462 ),
    .C(\i54/n471 ),
    .D(\i54/n488 ),
    .Y(\i54/n497 ));
 OAI211xp5_ASAP7_75t_SL \i54/i190  (.A1(\i54/n66 ),
    .A2(\i54/n75 ),
    .B(\i54/n157 ),
    .C(\i54/n535 ),
    .Y(\i54/n354 ));
 NOR2xp67_ASAP7_75t_SL \i54/i191  (.A(\i54/n211 ),
    .B(\i54/n265 ),
    .Y(\i54/n353 ));
 AO21x1_ASAP7_75t_SL \i54/i192  (.A1(\i54/n55 ),
    .A2(\i54/n162 ),
    .B(\i54/n510 ),
    .Y(\i54/n352 ));
 NAND2xp5_ASAP7_75t_SL \i54/i193  (.A(\i54/n248 ),
    .B(\i54/n224 ),
    .Y(\i54/n25 ));
 NOR2xp33_ASAP7_75t_SL \i54/i194  (.A(\i54/n249 ),
    .B(\i54/n266 ),
    .Y(\i54/n350 ));
 OAI211xp5_ASAP7_75t_SL \i54/i195  (.A1(\i54/n503 ),
    .A2(\i54/n75 ),
    .B(\i54/n192 ),
    .C(\i54/n536 ),
    .Y(\i54/n348 ));
 OR2x2_ASAP7_75t_SL \i54/i196  (.A(\i54/n203 ),
    .B(\i54/n541 ),
    .Y(\i54/n346 ));
 OAI211xp5_ASAP7_75t_SL \i54/i197  (.A1(\i54/n92 ),
    .A2(\i54/n79 ),
    .B(\i54/n189 ),
    .C(\i54/n139 ),
    .Y(\i54/n344 ));
 NAND2xp5_ASAP7_75t_SL \i54/i198  (.A(\i54/n267 ),
    .B(\i54/n268 ),
    .Y(\i54/n343 ));
 NAND2xp5_ASAP7_75t_SL \i54/i199  (.A(\i54/n23 ),
    .B(\i54/n199 ),
    .Y(\i54/n341 ));
 INVx1_ASAP7_75t_SL \i54/i2  (.A(\i54/n433 ),
    .Y(\i54/n2 ));
 NAND2x1_ASAP7_75t_SL \i54/i20  (.A(\i54/n450 ),
    .B(\i54/n481 ),
    .Y(\i54/n496 ));
 NAND2xp5_ASAP7_75t_SL \i54/i200  (.A(\i54/n245 ),
    .B(\i54/n567 ),
    .Y(\i54/n340 ));
 NAND2xp5_ASAP7_75t_SL \i54/i201  (.A(\i54/n186 ),
    .B(\i54/n564 ),
    .Y(\i54/n338 ));
 NOR2x1_ASAP7_75t_SL \i54/i202  (.A(\i54/n247 ),
    .B(\i54/n552 ),
    .Y(\i54/n336 ));
 INVx1_ASAP7_75t_SL \i54/i203  (.A(\i54/n312 ),
    .Y(\i54/n313 ));
 INVx1_ASAP7_75t_SL \i54/i204  (.A(\i54/n308 ),
    .Y(\i54/n309 ));
 INVx1_ASAP7_75t_SL \i54/i205  (.A(\i54/n304 ),
    .Y(\i54/n305 ));
 NAND4xp25_ASAP7_75t_SL \i54/i206  (.A(\i54/n120 ),
    .B(\i54/n140 ),
    .C(\i54/n126 ),
    .D(\i54/n568 ),
    .Y(\i54/n300 ));
 AOI31xp33_ASAP7_75t_SL \i54/i207  (.A1(\i54/n141 ),
    .A2(\i54/n71 ),
    .A3(\i54/n46 ),
    .B(\i54/n47 ),
    .Y(\i54/n299 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i54/i208  (.A1(\i54/n89 ),
    .A2(\i54/n52 ),
    .B(\i54/n68 ),
    .C(\i54/n146 ),
    .Y(\i54/n298 ));
 NOR4xp25_ASAP7_75t_SL \i54/i209  (.A(\i54/n117 ),
    .B(\i54/n538 ),
    .C(\i54/n556 ),
    .D(\i54/n95 ),
    .Y(\i54/n297 ));
 NOR2xp67_ASAP7_75t_SL \i54/i21  (.A(\i54/n443 ),
    .B(\i54/n482 ),
    .Y(\i54/n495 ));
 AOI211xp5_ASAP7_75t_SL \i54/i210  (.A1(\i54/n142 ),
    .A2(\i54/n82 ),
    .B(\i54/n178 ),
    .C(\i54/n104 ),
    .Y(\i54/n296 ));
 AOI21xp5_ASAP7_75t_SL \i54/i211  (.A1(\i54/n164 ),
    .A2(\i54/n89 ),
    .B(\i54/n238 ),
    .Y(\i54/n295 ));
 NOR2xp33_ASAP7_75t_L \i54/i212  (.A(\i54/n197 ),
    .B(\i54/n259 ),
    .Y(\i54/n294 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i54/i213  (.A1(\i54/n75 ),
    .A2(\i54/n51 ),
    .B(\i54/n84 ),
    .C(\i54/n235 ),
    .Y(\i54/n293 ));
 OAI22xp5_ASAP7_75t_SL \i54/i214  (.A1(\i54/n79 ),
    .A2(\i54/n166 ),
    .B1(\i54/n66 ),
    .B2(\i54/n102 ),
    .Y(\i54/n292 ));
 NOR2xp33_ASAP7_75t_SL \i54/i215  (.A(\i54/n217 ),
    .B(\i54/n543 ),
    .Y(\i54/n291 ));
 OAI222xp33_ASAP7_75t_SL \i54/i216  (.A1(\i54/n87 ),
    .A2(\i54/n47 ),
    .B1(\i54/n51 ),
    .B2(\i54/n14 ),
    .C1(\i54/n71 ),
    .C2(\i54/n66 ),
    .Y(\i54/n290 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i54/i217  (.A1(\i54/n60 ),
    .A2(\i54/n57 ),
    .B(\i54/n5 ),
    .C(\i54/n175 ),
    .Y(\i54/n289 ));
 NAND2xp33_ASAP7_75t_L \i54/i218  (.A(\i54/n116 ),
    .B(\i54/n208 ),
    .Y(\i54/n288 ));
 NAND2xp33_ASAP7_75t_SL \i54/i219  (.A(\i54/n255 ),
    .B(\i54/n557 ),
    .Y(\i54/n287 ));
 NAND4xp75_ASAP7_75t_SL \i54/i22  (.A(\i54/n454 ),
    .B(\i54/n466 ),
    .C(\i54/n448 ),
    .D(\i54/n451 ),
    .Y(\i54/n494 ));
 AOI22xp5_ASAP7_75t_SL \i54/i220  (.A1(\i54/n74 ),
    .A2(\i54/n113 ),
    .B1(\i54/n82 ),
    .B2(\i54/n76 ),
    .Y(\i54/n286 ));
 OAI21xp5_ASAP7_75t_SL \i54/i221  (.A1(\i54/n124 ),
    .A2(\i54/n74 ),
    .B(\i54/n82 ),
    .Y(\i54/n285 ));
 OA21x2_ASAP7_75t_SL \i54/i222  (.A1(\i54/n47 ),
    .A2(\i54/n145 ),
    .B(\i54/n134 ),
    .Y(\i54/n284 ));
 NAND2xp5_ASAP7_75t_SL \i54/i223  (.A(\i54/n204 ),
    .B(\i54/n272 ),
    .Y(\i54/n283 ));
 NAND4xp25_ASAP7_75t_SL \i54/i224  (.A(\i54/n136 ),
    .B(\i54/n560 ),
    .C(\i54/n110 ),
    .D(\i54/n108 ),
    .Y(\i54/n282 ));
 AOI221xp5_ASAP7_75t_SL \i54/i225  (.A1(\i54/n62 ),
    .A2(\i54/n45 ),
    .B1(\i54/n52 ),
    .B2(\i54/n65 ),
    .C(\i54/n539 ),
    .Y(\i54/n281 ));
 OAI221xp5_ASAP7_75t_SL \i54/i226  (.A1(\i54/n91 ),
    .A2(\i54/n84 ),
    .B1(\i54/n69 ),
    .B2(\i54/n515 ),
    .C(\i54/n115 ),
    .Y(\i54/n315 ));
 OAI221xp5_ASAP7_75t_SL \i54/i227  (.A1(\i54/n87 ),
    .A2(\i54/n77 ),
    .B1(\i54/n69 ),
    .B2(\i54/n67 ),
    .C(\i54/n218 ),
    .Y(\i54/n280 ));
 AND3x1_ASAP7_75t_SL \i54/i228  (.A(\i54/n133 ),
    .B(\i54/n140 ),
    .C(\i54/n240 ),
    .Y(\i54/n279 ));
 NAND2xp33_ASAP7_75t_SL \i54/i229  (.A(\i54/n206 ),
    .B(\i54/n241 ),
    .Y(\i54/n278 ));
 OR3x1_ASAP7_75t_SL \i54/i23  (.A(\i54/n474 ),
    .B(\i54/n472 ),
    .C(\i54/n455 ),
    .Y(\i54/n493 ));
 OAI221xp5_ASAP7_75t_SL \i54/i230  (.A1(\i54/n87 ),
    .A2(\i54/n81 ),
    .B1(\i54/n15 ),
    .B2(\i54/n14 ),
    .C(\i54/n254 ),
    .Y(\i54/n277 ));
 OAI222xp33_ASAP7_75t_SL \i54/i231  (.A1(\i54/n79 ),
    .A2(\i54/n81 ),
    .B1(\i54/n91 ),
    .B2(\i54/n77 ),
    .C1(\i54/n15 ),
    .C2(\i54/n503 ),
    .Y(\i54/n314 ));
 NAND3x1_ASAP7_75t_SL \i54/i232  (.A(\i54/n209 ),
    .B(\i54/n558 ),
    .C(\i54/n554 ),
    .Y(\i54/n312 ));
 AOI22xp5_ASAP7_75t_SL \i54/i233  (.A1(\i54/n517 ),
    .A2(\i54/n90 ),
    .B1(\i54/n68 ),
    .B2(\i54/n54 ),
    .Y(\i54/n311 ));
 AOI22xp5_ASAP7_75t_SL \i54/i234  (.A1(\i54/n93 ),
    .A2(\i54/n525 ),
    .B1(\i54/n48 ),
    .B2(\i54/n72 ),
    .Y(\i54/n310 ));
 AOI221x1_ASAP7_75t_SL \i54/i235  (.A1(\i54/n90 ),
    .A2(\i54/n68 ),
    .B1(\i54/n76 ),
    .B2(\i54/n78 ),
    .C(\i54/n242 ),
    .Y(\i54/n308 ));
 AOI211x1_ASAP7_75t_SL \i54/i236  (.A1(\i54/n107 ),
    .A2(\i54/n64 ),
    .B(\i54/n190 ),
    .C(\i54/n556 ),
    .Y(\i54/n307 ));
 OAI21xp5_ASAP7_75t_SL \i54/i237  (.A1(\i54/n46 ),
    .A2(\i54/n84 ),
    .B(\i54/n250 ),
    .Y(\i54/n306 ));
 NOR2x1_ASAP7_75t_SL \i54/i238  (.A(\i54/n135 ),
    .B(\i54/n202 ),
    .Y(\i54/n304 ));
 OAI221xp5_ASAP7_75t_SL \i54/i239  (.A1(\i54/n512 ),
    .A2(\i54/n91 ),
    .B1(\i54/n61 ),
    .B2(\i54/n67 ),
    .C(\i54/n170 ),
    .Y(\i54/n303 ));
 OR3x1_ASAP7_75t_SL \i54/i24  (.A(\i54/n475 ),
    .B(\i54/n441 ),
    .C(\i54/n415 ),
    .Y(\i54/n492 ));
 OAI211xp5_ASAP7_75t_SL \i54/i240  (.A1(\i54/n67 ),
    .A2(\i54/n565 ),
    .B(\i54/n119 ),
    .C(\i54/n562 ),
    .Y(\i54/n302 ));
 NOR2x1_ASAP7_75t_SL \i54/i241  (.A(\i54/n146 ),
    .B(\i54/n544 ),
    .Y(\i54/n24 ));
 NOR2xp33_ASAP7_75t_SL \i54/i242  (.A(\i54/n148 ),
    .B(\i54/n269 ),
    .Y(\i54/n276 ));
 OAI221xp5_ASAP7_75t_SL \i54/i243  (.A1(\i54/n58 ),
    .A2(\i54/n51 ),
    .B1(\i54/n47 ),
    .B2(\i54/n55 ),
    .C(\i54/n129 ),
    .Y(\i54/n301 ));
 INVx1_ASAP7_75t_SL \i54/i244  (.A(\i54/n567 ),
    .Y(\i54/n274 ));
 INVx1_ASAP7_75t_SL \i54/i245  (.A(\i54/n271 ),
    .Y(\i54/n272 ));
 INVx1_ASAP7_75t_SL \i54/i246  (.A(\i54/n269 ),
    .Y(\i54/n270 ));
 INVxp67_ASAP7_75t_SL \i54/i247  (.A(\i54/n262 ),
    .Y(\i54/n263 ));
 INVx1_ASAP7_75t_SL \i54/i248  (.A(\i54/n259 ),
    .Y(\i54/n260 ));
 OAI21xp33_ASAP7_75t_SL \i54/i249  (.A1(\i54/n73 ),
    .A2(\i54/n529 ),
    .B(\i54/n508 ),
    .Y(\i54/n257 ));
 NAND3xp33_ASAP7_75t_SL \i54/i25  (.A(\i54/n486 ),
    .B(\i54/n471 ),
    .C(\i54/n454 ),
    .Y(\i54/n491 ));
 NAND2xp5_ASAP7_75t_SL \i54/i250  (.A(\i54/n570 ),
    .B(\i54/n139 ),
    .Y(\i54/n256 ));
 OAI21xp5_ASAP7_75t_SL \i54/i251  (.A1(\i54/n54 ),
    .A2(\i54/n53 ),
    .B(\i54/n85 ),
    .Y(\i54/n255 ));
 NOR2xp33_ASAP7_75t_SL \i54/i252  (.A(\i54/n149 ),
    .B(\i54/n559 ),
    .Y(\i54/n254 ));
 NAND2xp33_ASAP7_75t_L \i54/i253  (.A(\i54/n566 ),
    .B(\i54/n105 ),
    .Y(\i54/n253 ));
 OAI21xp33_ASAP7_75t_SL \i54/i254  (.A1(\i54/n70 ),
    .A2(\i54/n57 ),
    .B(\i54/n50 ),
    .Y(\i54/n252 ));
 NOR2x1_ASAP7_75t_SL \i54/i255  (.A(\i54/n17 ),
    .B(\i54/n127 ),
    .Y(\i54/n251 ));
 OAI21xp5_ASAP7_75t_SL \i54/i256  (.A1(\i54/n74 ),
    .A2(\i54/n83 ),
    .B(\i54/n62 ),
    .Y(\i54/n250 ));
 OAI21xp5_ASAP7_75t_SL \i54/i257  (.A1(\i54/n58 ),
    .A2(\i54/n88 ),
    .B(\i54/n176 ),
    .Y(\i54/n249 ));
 AOI22xp5_ASAP7_75t_SL \i54/i258  (.A1(\i54/n85 ),
    .A2(\i54/n57 ),
    .B1(\i54/n78 ),
    .B2(\i54/n72 ),
    .Y(\i54/n248 ));
 OAI21xp5_ASAP7_75t_SL \i54/i259  (.A1(\i54/n14 ),
    .A2(\i54/n69 ),
    .B(\i54/n143 ),
    .Y(\i54/n247 ));
 NOR2x1_ASAP7_75t_SL \i54/i26  (.A(\i54/n395 ),
    .B(\i54/n472 ),
    .Y(\i54/n489 ));
 OAI21xp5_ASAP7_75t_SL \i54/i260  (.A1(\i54/n74 ),
    .A2(\i54/n53 ),
    .B(\i54/n65 ),
    .Y(\i54/n246 ));
 AOI22xp5_ASAP7_75t_SL \i54/i261  (.A1(\i54/n45 ),
    .A2(\i54/n93 ),
    .B1(\i54/n48 ),
    .B2(\i54/n74 ),
    .Y(\i54/n245 ));
 OA21x2_ASAP7_75t_SL \i54/i262  (.A1(\i54/n63 ),
    .A2(\i54/n13 ),
    .B(\i54/n509 ),
    .Y(\i54/n275 ));
 AOI21xp33_ASAP7_75t_SL \i54/i263  (.A1(\i54/n66 ),
    .A2(\i54/n63 ),
    .B(\i54/n46 ),
    .Y(\i54/n244 ));
 OAI21xp5_ASAP7_75t_SL \i54/i264  (.A1(\i54/n78 ),
    .A2(\i54/n93 ),
    .B(\i54/n86 ),
    .Y(\i54/n243 ));
 OA21x2_ASAP7_75t_SL \i54/i265  (.A1(\i54/n5 ),
    .A2(\i54/n93 ),
    .B(\i54/n89 ),
    .Y(\i54/n242 ));
 OAI21xp5_ASAP7_75t_SL \i54/i266  (.A1(\i54/n65 ),
    .A2(\i54/n48 ),
    .B(\i54/n86 ),
    .Y(\i54/n241 ));
 OAI21xp5_ASAP7_75t_SL \i54/i267  (.A1(\i54/n74 ),
    .A2(\i54/n70 ),
    .B(\i54/n93 ),
    .Y(\i54/n240 ));
 AOI21xp33_ASAP7_75t_SL \i54/i268  (.A1(\i54/n503 ),
    .A2(\i54/n84 ),
    .B(\i54/n46 ),
    .Y(\i54/n239 ));
 OAI21xp5_ASAP7_75t_SL \i54/i269  (.A1(\i54/n58 ),
    .A2(\i54/n69 ),
    .B(\i54/n21 ),
    .Y(\i54/n238 ));
 NOR2x1_ASAP7_75t_SL \i54/i27  (.A(\i54/n456 ),
    .B(\i54/n452 ),
    .Y(\i54/n488 ));
 AOI21xp33_ASAP7_75t_SL \i54/i270  (.A1(\i54/n75 ),
    .A2(\i54/n46 ),
    .B(\i54/n67 ),
    .Y(\i54/n237 ));
 OAI21xp5_ASAP7_75t_SL \i54/i271  (.A1(\i54/n89 ),
    .A2(\i54/n74 ),
    .B(\i54/n50 ),
    .Y(\i54/n236 ));
 OAI21xp5_ASAP7_75t_SL \i54/i272  (.A1(\i54/n70 ),
    .A2(\i54/n60 ),
    .B(\i54/n78 ),
    .Y(\i54/n235 ));
 NAND2xp5_ASAP7_75t_SL \i54/i273  (.A(\i54/n86 ),
    .B(\i54/n164 ),
    .Y(\i54/n23 ));
 NAND2xp5_ASAP7_75t_L \i54/i274  (.A(\i54/n192 ),
    .B(\i54/n536 ),
    .Y(\i54/n234 ));
 OAI22xp5_ASAP7_75t_SL \i54/i275  (.A1(\i54/n529 ),
    .A2(\i54/n87 ),
    .B1(\i54/n94 ),
    .B2(\i54/n13 ),
    .Y(\i54/n273 ));
 OAI22xp33_ASAP7_75t_SL \i54/i276  (.A1(\i54/n94 ),
    .A2(\i54/n69 ),
    .B1(\i54/n15 ),
    .B2(\i54/n66 ),
    .Y(\i54/n271 ));
 OAI22xp5_ASAP7_75t_SL \i54/i277  (.A1(\i54/n92 ),
    .A2(\i54/n56 ),
    .B1(\i54/n58 ),
    .B2(\i54/n79 ),
    .Y(\i54/n269 ));
 AOI22xp5_ASAP7_75t_SL \i54/i278  (.A1(\i54/n64 ),
    .A2(\i54/n90 ),
    .B1(\i54/n5 ),
    .B2(\i54/n83 ),
    .Y(\i54/n268 ));
 AOI22xp5_ASAP7_75t_SL \i54/i279  (.A1(\i54/n64 ),
    .A2(\i54/n60 ),
    .B1(\i54/n520 ),
    .B2(\i54/n57 ),
    .Y(\i54/n267 ));
 NAND3xp33_ASAP7_75t_SL \i54/i28  (.A(\i54/n436 ),
    .B(\i54/n581 ),
    .C(\i54/n434 ),
    .Y(\i54/n487 ));
 OAI22xp5_ASAP7_75t_SL \i54/i280  (.A1(\i54/n67 ),
    .A2(\i54/n79 ),
    .B1(\i54/n69 ),
    .B2(\i54/n49 ),
    .Y(\i54/n266 ));
 OAI22xp33_ASAP7_75t_SL \i54/i281  (.A1(\i54/n94 ),
    .A2(\i54/n91 ),
    .B1(\i54/n47 ),
    .B2(\i54/n523 ),
    .Y(\i54/n265 ));
 NAND2xp5_ASAP7_75t_L \i54/i282  (.A(\i54/n16 ),
    .B(\i54/n160 ),
    .Y(\i54/n264 ));
 OAI22xp5_ASAP7_75t_SL \i54/i283  (.A1(\i54/n58 ),
    .A2(\i54/n91 ),
    .B1(\i54/n66 ),
    .B2(\i54/n88 ),
    .Y(\i54/n262 ));
 OAI21xp5_ASAP7_75t_SL \i54/i284  (.A1(\i54/n74 ),
    .A2(\i54/n52 ),
    .B(\i54/n85 ),
    .Y(\i54/n261 ));
 NOR2xp33_ASAP7_75t_L \i54/i285  (.A(\i54/n13 ),
    .B(\i54/n512 ),
    .Y(\i54/n259 ));
 NAND2xp33_ASAP7_75t_L \i54/i286  (.A(\i54/n119 ),
    .B(\i54/n562 ),
    .Y(\i54/n233 ));
 OAI21xp5_ASAP7_75t_SL \i54/i287  (.A1(\i54/n67 ),
    .A2(\i54/n56 ),
    .B(\i54/n118 ),
    .Y(\i54/n258 ));
 INVxp67_ASAP7_75t_SL \i54/i288  (.A(\i54/n229 ),
    .Y(\i54/n230 ));
 INVxp67_ASAP7_75t_SL \i54/i289  (.A(\i54/n227 ),
    .Y(\i54/n228 ));
 NOR2x1_ASAP7_75t_SL \i54/i29  (.A(\i54/n461 ),
    .B(\i54/n424 ),
    .Y(\i54/n486 ));
 INVx1_ASAP7_75t_SL \i54/i290  (.A(\i54/n225 ),
    .Y(\i54/n226 ));
 INVx1_ASAP7_75t_SL \i54/i291  (.A(\i54/n222 ),
    .Y(\i54/n223 ));
 INVxp67_ASAP7_75t_SL \i54/i292  (.A(\i54/n220 ),
    .Y(\i54/n221 ));
 INVxp67_ASAP7_75t_SL \i54/i293  (.A(\i54/n217 ),
    .Y(\i54/n218 ));
 INVxp67_ASAP7_75t_SL \i54/i294  (.A(\i54/n215 ),
    .Y(\i54/n216 ));
 OAI22xp33_ASAP7_75t_SL \i54/i295  (.A1(\i54/n49 ),
    .A2(\i54/n91 ),
    .B1(\i54/n55 ),
    .B2(\i54/n529 ),
    .Y(\i54/n211 ));
 OAI21xp5_ASAP7_75t_SL \i54/i296  (.A1(\i54/n57 ),
    .A2(\i54/n80 ),
    .B(\i54/n78 ),
    .Y(\i54/n210 ));
 OAI21xp5_ASAP7_75t_SL \i54/i297  (.A1(\i54/n59 ),
    .A2(\i54/n68 ),
    .B(\i54/n70 ),
    .Y(\i54/n209 ));
 OAI21xp5_ASAP7_75t_SL \i54/i298  (.A1(\i54/n54 ),
    .A2(\i54/n52 ),
    .B(\i54/n59 ),
    .Y(\i54/n208 ));
 AOI21xp33_ASAP7_75t_SL \i54/i299  (.A1(\i54/n69 ),
    .A2(\i54/n79 ),
    .B(\i54/n81 ),
    .Y(\i54/n207 ));
 INVx2_ASAP7_75t_SL \i54/i3  (.A(\i54/n33 ),
    .Y(\i54/n3 ));
 NOR5xp2_ASAP7_75t_SL \i54/i30  (.A(\i54/n426 ),
    .B(\i54/n374 ),
    .C(\i54/n417 ),
    .D(\i54/n340 ),
    .E(\i54/n344 ),
    .Y(\i54/n485 ));
 OAI21xp5_ASAP7_75t_SL \i54/i300  (.A1(\i54/n45 ),
    .A2(\i54/n52 ),
    .B(\i54/n50 ),
    .Y(\i54/n206 ));
 OAI21xp5_ASAP7_75t_SL \i54/i301  (.A1(\i54/n82 ),
    .A2(\i54/n59 ),
    .B(\i54/n54 ),
    .Y(\i54/n205 ));
 AOI22xp33_ASAP7_75t_SL \i54/i302  (.A1(\i54/n64 ),
    .A2(\i54/n74 ),
    .B1(\i54/n5 ),
    .B2(\i54/n54 ),
    .Y(\i54/n204 ));
 OAI22xp33_ASAP7_75t_SL \i54/i303  (.A1(\i54/n529 ),
    .A2(\i54/n46 ),
    .B1(\i54/n87 ),
    .B2(\i54/n503 ),
    .Y(\i54/n203 ));
 AOI22xp5_ASAP7_75t_SL \i54/i304  (.A1(\i54/n520 ),
    .A2(\i54/n86 ),
    .B1(\i54/n85 ),
    .B2(\i54/n53 ),
    .Y(\i54/n232 ));
 OAI22xp5_ASAP7_75t_L \i54/i305  (.A1(\i54/n15 ),
    .A2(\i54/n529 ),
    .B1(\i54/n79 ),
    .B2(\i54/n84 ),
    .Y(\i54/n202 ));
 OAI22xp5_ASAP7_75t_SL \i54/i306  (.A1(\i54/n92 ),
    .A2(\i54/n523 ),
    .B1(\i54/n515 ),
    .B2(\i54/n87 ),
    .Y(\i54/n201 ));
 OAI22xp33_ASAP7_75t_SL \i54/i307  (.A1(\i54/n503 ),
    .A2(\i54/n523 ),
    .B1(\i54/n84 ),
    .B2(\i54/n75 ),
    .Y(\i54/n200 ));
 AOI22xp5_ASAP7_75t_SL \i54/i308  (.A1(\i54/n45 ),
    .A2(\i54/n48 ),
    .B1(\i54/n520 ),
    .B2(\i54/n74 ),
    .Y(\i54/n231 ));
 AOI22xp5_ASAP7_75t_SL \i54/i309  (.A1(\i54/n62 ),
    .A2(\i54/n80 ),
    .B1(\i54/n48 ),
    .B2(\i54/n83 ),
    .Y(\i54/n199 ));
 NOR3xp33_ASAP7_75t_SL \i54/i31  (.A(\i54/n422 ),
    .B(\i54/n438 ),
    .C(\i54/n470 ),
    .Y(\i54/n484 ));
 OAI22xp5_ASAP7_75t_SL \i54/i310  (.A1(\i54/n529 ),
    .A2(\i54/n91 ),
    .B1(\i54/n66 ),
    .B2(\i54/n13 ),
    .Y(\i54/n198 ));
 OAI21xp33_ASAP7_75t_SL \i54/i311  (.A1(\i54/n55 ),
    .A2(\i54/n77 ),
    .B(\i54/n557 ),
    .Y(\i54/n197 ));
 OAI21xp5_ASAP7_75t_SL \i54/i312  (.A1(\i54/n47 ),
    .A2(\i54/n56 ),
    .B(\i54/n128 ),
    .Y(\i54/n229 ));
 AOI22xp5_ASAP7_75t_SL \i54/i313  (.A1(\i54/n45 ),
    .A2(\i54/n65 ),
    .B1(\i54/n48 ),
    .B2(\i54/n53 ),
    .Y(\i54/n227 ));
 AOI22xp5_ASAP7_75t_SL \i54/i314  (.A1(\i54/n50 ),
    .A2(\i54/n52 ),
    .B1(\i54/n60 ),
    .B2(\i54/n62 ),
    .Y(\i54/n225 ));
 AOI22xp5_ASAP7_75t_SL \i54/i315  (.A1(\i54/n89 ),
    .A2(\i54/n520 ),
    .B1(\i54/n82 ),
    .B2(\i54/n72 ),
    .Y(\i54/n224 ));
 OAI22xp5_ASAP7_75t_SL \i54/i316  (.A1(\i54/n46 ),
    .A2(\i54/n515 ),
    .B1(\i54/n529 ),
    .B2(\i54/n71 ),
    .Y(\i54/n196 ));
 NAND2xp33_ASAP7_75t_SL \i54/i317  (.A(\i54/n193 ),
    .B(\i54/n194 ),
    .Y(\i54/n195 ));
 OAI22x1_ASAP7_75t_SL \i54/i318  (.A1(\i54/n14 ),
    .A2(\i54/n91 ),
    .B1(\i54/n49 ),
    .B2(\i54/n73 ),
    .Y(\i54/n222 ));
 AOI22xp5_ASAP7_75t_SL \i54/i319  (.A1(\i54/n50 ),
    .A2(\i54/n60 ),
    .B1(\i54/n48 ),
    .B2(\i54/n89 ),
    .Y(\i54/n220 ));
 NOR2x1_ASAP7_75t_SL \i54/i32  (.A(\i54/n467 ),
    .B(\i54/n427 ),
    .Y(\i54/n483 ));
 OAI21xp5_ASAP7_75t_SL \i54/i320  (.A1(\i54/n77 ),
    .A2(\i54/n51 ),
    .B(\i54/n112 ),
    .Y(\i54/n219 ));
 OAI22xp5_ASAP7_75t_L \i54/i321  (.A1(\i54/n81 ),
    .A2(\i54/n46 ),
    .B1(\i54/n79 ),
    .B2(\i54/n47 ),
    .Y(\i54/n217 ));
 OAI22xp5_ASAP7_75t_SL \i54/i322  (.A1(\i54/n503 ),
    .A2(\i54/n51 ),
    .B1(\i54/n66 ),
    .B2(\i54/n79 ),
    .Y(\i54/n215 ));
 AOI22xp5_ASAP7_75t_SL \i54/i323  (.A1(\i54/n45 ),
    .A2(\i54/n50 ),
    .B1(\i54/n68 ),
    .B2(\i54/n83 ),
    .Y(\i54/n214 ));
 OAI22xp5_ASAP7_75t_SL \i54/i324  (.A1(\i54/n75 ),
    .A2(\i54/n529 ),
    .B1(\i54/n71 ),
    .B2(\i54/n63 ),
    .Y(\i54/n213 ));
 OAI22x1_ASAP7_75t_SL \i54/i325  (.A1(\i54/n63 ),
    .A2(\i54/n79 ),
    .B1(\i54/n67 ),
    .B2(\i54/n87 ),
    .Y(\i54/n22 ));
 AOI22xp5_ASAP7_75t_SL \i54/i326  (.A1(\i54/n59 ),
    .A2(\i54/n83 ),
    .B1(\i54/n48 ),
    .B2(\i54/n60 ),
    .Y(\i54/n212 ));
 INVxp67_ASAP7_75t_SL \i54/i327  (.A(\i54/n190 ),
    .Y(\i54/n191 ));
 INVx1_ASAP7_75t_SL \i54/i328  (.A(\i54/n188 ),
    .Y(\i54/n189 ));
 INVxp67_ASAP7_75t_SL \i54/i329  (.A(\i54/n186 ),
    .Y(\i54/n187 ));
 NAND2xp5_ASAP7_75t_SL \i54/i33  (.A(\i54/n425 ),
    .B(\i54/n444 ),
    .Y(\i54/n482 ));
 INVxp67_ASAP7_75t_SL \i54/i330  (.A(\i54/n184 ),
    .Y(\i54/n185 ));
 INVxp67_ASAP7_75t_SL \i54/i331  (.A(\i54/n508 ),
    .Y(\i54/n183 ));
 INVxp67_ASAP7_75t_SL \i54/i332  (.A(\i54/n180 ),
    .Y(\i54/n181 ));
 INVxp67_ASAP7_75t_SL \i54/i333  (.A(\i54/n176 ),
    .Y(\i54/n177 ));
 INVxp67_ASAP7_75t_SL \i54/i334  (.A(\i54/n566 ),
    .Y(\i54/n175 ));
 INVxp67_ASAP7_75t_SL \i54/i335  (.A(\i54/n172 ),
    .Y(\i54/n173 ));
 INVxp67_ASAP7_75t_SL \i54/i336  (.A(\i54/n170 ),
    .Y(\i54/n171 ));
 INVxp67_ASAP7_75t_SL \i54/i337  (.A(\i54/n168 ),
    .Y(\i54/n169 ));
 INVxp67_ASAP7_75t_SL \i54/i338  (.A(\i54/n166 ),
    .Y(\i54/n167 ));
 INVxp67_ASAP7_75t_SL \i54/i339  (.A(\i54/n512 ),
    .Y(\i54/n165 ));
 NOR3x1_ASAP7_75t_SL \i54/i34  (.A(\i54/n26 ),
    .B(\i54/n440 ),
    .C(\i54/n366 ),
    .Y(\i54/n490 ));
 INVx1_ASAP7_75t_SL \i54/i340  (.A(\i54/n164 ),
    .Y(\i54/n163 ));
 NAND2xp5_ASAP7_75t_SL \i54/i341  (.A(\i54/n65 ),
    .B(\i54/n86 ),
    .Y(\i54/n194 ));
 NAND2xp5_ASAP7_75t_SL \i54/i342  (.A(\i54/n85 ),
    .B(\i54/n83 ),
    .Y(\i54/n162 ));
 NAND2xp5_ASAP7_75t_SL \i54/i343  (.A(\i54/n84 ),
    .B(\i54/n81 ),
    .Y(\i54/n161 ));
 NAND2xp5_ASAP7_75t_SL \i54/i344  (.A(\i54/n48 ),
    .B(\i54/n90 ),
    .Y(\i54/n160 ));
 NAND2xp33_ASAP7_75t_SL \i54/i345  (.A(\i54/n503 ),
    .B(\i54/n58 ),
    .Y(\i54/n159 ));
 NAND2xp5_ASAP7_75t_SL \i54/i346  (.A(\i54/n57 ),
    .B(\i54/n62 ),
    .Y(\i54/n193 ));
 NAND2xp5_ASAP7_75t_SL \i54/i347  (.A(\i54/n62 ),
    .B(\i54/n86 ),
    .Y(\i54/n158 ));
 NAND2xp5_ASAP7_75t_SL \i54/i348  (.A(\i54/n85 ),
    .B(\i54/n89 ),
    .Y(\i54/n157 ));
 NAND2xp5_ASAP7_75t_SL \i54/i349  (.A(\i54/n72 ),
    .B(\i54/n68 ),
    .Y(\i54/n156 ));
 NOR3xp33_ASAP7_75t_SL \i54/i35  (.A(\i54/n383 ),
    .B(\i54/n26 ),
    .C(\i54/n464 ),
    .Y(\i54/n480 ));
 NAND2xp5_ASAP7_75t_SL \i54/i350  (.A(\i54/n62 ),
    .B(\i54/n72 ),
    .Y(\i54/n155 ));
 NAND2xp5_ASAP7_75t_SL \i54/i351  (.A(\i54/n65 ),
    .B(\i54/n89 ),
    .Y(\i54/n154 ));
 NAND2xp5_ASAP7_75t_SL \i54/i352  (.A(\i54/n45 ),
    .B(\i54/n78 ),
    .Y(\i54/n192 ));
 AND2x2_ASAP7_75t_SL \i54/i353  (.A(\i54/n85 ),
    .B(\i54/n70 ),
    .Y(\i54/n190 ));
 AND2x2_ASAP7_75t_SL \i54/i354  (.A(\i54/n520 ),
    .B(\i54/n72 ),
    .Y(\i54/n188 ));
 NAND2xp5_ASAP7_75t_SL \i54/i355  (.A(\i54/n72 ),
    .B(\i54/n5 ),
    .Y(\i54/n21 ));
 NAND2xp5_ASAP7_75t_SL \i54/i356  (.A(\i54/n78 ),
    .B(\i54/n89 ),
    .Y(\i54/n186 ));
 NAND2xp5_ASAP7_75t_SL \i54/i357  (.A(\i54/n93 ),
    .B(\i54/n52 ),
    .Y(\i54/n184 ));
 AND2x2_ASAP7_75t_SL \i54/i358  (.A(\i54/n65 ),
    .B(\i54/n60 ),
    .Y(\i54/n182 ));
 NOR2xp67_ASAP7_75t_SL \i54/i359  (.A(\i54/n63 ),
    .B(\i54/n69 ),
    .Y(\i54/n20 ));
 NOR2xp67_ASAP7_75t_SL \i54/i36  (.A(\i54/n445 ),
    .B(\i54/n26 ),
    .Y(\i54/n479 ));
 NOR2xp67_ASAP7_75t_L \i54/i360  (.A(\i54/n55 ),
    .B(\i54/n63 ),
    .Y(\i54/n180 ));
 NAND2xp5_ASAP7_75t_SL \i54/i361  (.A(\i54/n76 ),
    .B(\i54/n64 ),
    .Y(\i54/n179 ));
 NOR2xp33_ASAP7_75t_SL \i54/i362  (.A(\i54/n67 ),
    .B(\i54/n79 ),
    .Y(\i54/n153 ));
 NOR2xp33_ASAP7_75t_SL \i54/i363  (.A(\i54/n529 ),
    .B(\i54/n79 ),
    .Y(\i54/n178 ));
 NOR2xp33_ASAP7_75t_SL \i54/i364  (.A(\i54/n14 ),
    .B(\i54/n13 ),
    .Y(\i54/n152 ));
 NAND2xp5_ASAP7_75t_SL \i54/i365  (.A(\i54/n64 ),
    .B(\i54/n52 ),
    .Y(\i54/n176 ));
 NOR2xp33_ASAP7_75t_SL \i54/i366  (.A(\i54/n529 ),
    .B(\i54/n88 ),
    .Y(\i54/n151 ));
 NOR2xp33_ASAP7_75t_L \i54/i367  (.A(\i54/n93 ),
    .B(\i54/n50 ),
    .Y(\i54/n174 ));
 NAND2xp5_ASAP7_75t_SL \i54/i368  (.A(\i54/n93 ),
    .B(\i54/n53 ),
    .Y(\i54/n172 ));
 NAND2xp5_ASAP7_75t_SL \i54/i369  (.A(\i54/n89 ),
    .B(\i54/n62 ),
    .Y(\i54/n170 ));
 NOR3xp33_ASAP7_75t_SL \i54/i37  (.A(\i54/n423 ),
    .B(\i54/n418 ),
    .C(\i54/n2 ),
    .Y(\i54/n478 ));
 NAND2xp5_ASAP7_75t_SL \i54/i370  (.A(\i54/n93 ),
    .B(\i54/n72 ),
    .Y(\i54/n168 ));
 NAND2xp5_ASAP7_75t_SL \i54/i371  (.A(\i54/n65 ),
    .B(\i54/n76 ),
    .Y(\i54/n150 ));
 NOR2xp33_ASAP7_75t_SL \i54/i372  (.A(\i54/n85 ),
    .B(\i54/n65 ),
    .Y(\i54/n166 ));
 NOR2xp33_ASAP7_75t_SL \i54/i373  (.A(\i54/n56 ),
    .B(\i54/n84 ),
    .Y(\i54/n149 ));
 OR2x2_ASAP7_75t_SL \i54/i374  (.A(\i54/n64 ),
    .B(\i54/n50 ),
    .Y(\i54/n164 ));
 INVxp67_ASAP7_75t_SL \i54/i375  (.A(\i54/n147 ),
    .Y(\i54/n148 ));
 INVxp67_ASAP7_75t_SL \i54/i376  (.A(\i54/n143 ),
    .Y(\i54/n144 ));
 INVx1_ASAP7_75t_SL \i54/i377  (.A(\i54/n141 ),
    .Y(\i54/n142 ));
 INVxp67_ASAP7_75t_SL \i54/i378  (.A(\i54/n136 ),
    .Y(\i54/n137 ));
 INVxp67_ASAP7_75t_SL \i54/i379  (.A(\i54/n134 ),
    .Y(\i54/n135 ));
 NAND4xp25_ASAP7_75t_SL \i54/i38  (.A(\i54/n405 ),
    .B(\i54/n399 ),
    .C(\i54/n398 ),
    .D(\i54/n432 ),
    .Y(\i54/n477 ));
 INVxp67_ASAP7_75t_SL \i54/i380  (.A(\i54/n538 ),
    .Y(\i54/n133 ));
 INVxp67_ASAP7_75t_SL \i54/i381  (.A(\i54/n131 ),
    .Y(\i54/n132 ));
 INVxp67_ASAP7_75t_SL \i54/i382  (.A(\i54/n129 ),
    .Y(\i54/n130 ));
 INVxp67_ASAP7_75t_SL \i54/i383  (.A(\i54/n127 ),
    .Y(\i54/n128 ));
 INVxp67_ASAP7_75t_SL \i54/i384  (.A(\i54/n120 ),
    .Y(\i54/n121 ));
 INVx1_ASAP7_75t_SL \i54/i385  (.A(\i54/n116 ),
    .Y(\i54/n117 ));
 INVx1_ASAP7_75t_SL \i54/i386  (.A(\i54/n16 ),
    .Y(\i54/n17 ));
 NAND2xp5_ASAP7_75t_SL \i54/i387  (.A(\i54/n82 ),
    .B(\i54/n74 ),
    .Y(\i54/n115 ));
 NAND2xp5_ASAP7_75t_SL \i54/i388  (.A(\i54/n50 ),
    .B(\i54/n76 ),
    .Y(\i54/n114 ));
 NAND2xp5_ASAP7_75t_SL \i54/i389  (.A(\i54/n59 ),
    .B(\i54/n74 ),
    .Y(\i54/n19 ));
 NAND3xp33_ASAP7_75t_L \i54/i39  (.A(\i54/n381 ),
    .B(\i54/n399 ),
    .C(\i54/n449 ),
    .Y(\i54/n476 ));
 NAND2xp5_ASAP7_75t_SL \i54/i390  (.A(\i54/n77 ),
    .B(\i54/n67 ),
    .Y(\i54/n113 ));
 NAND2xp5_ASAP7_75t_SL \i54/i391  (.A(\i54/n59 ),
    .B(\i54/n76 ),
    .Y(\i54/n112 ));
 NAND2xp33_ASAP7_75t_SL \i54/i392  (.A(\i54/n76 ),
    .B(\i54/n48 ),
    .Y(\i54/n111 ));
 NAND2xp5_ASAP7_75t_SL \i54/i393  (.A(\i54/n78 ),
    .B(\i54/n60 ),
    .Y(\i54/n110 ));
 NAND2xp5_ASAP7_75t_SL \i54/i394  (.A(\i54/n68 ),
    .B(\i54/n53 ),
    .Y(\i54/n109 ));
 NAND2xp5_ASAP7_75t_SL \i54/i395  (.A(\i54/n48 ),
    .B(\i54/n70 ),
    .Y(\i54/n108 ));
 NAND2xp5_ASAP7_75t_L \i54/i396  (.A(\i54/n15 ),
    .B(\i54/n46 ),
    .Y(\i54/n107 ));
 NAND2xp5_ASAP7_75t_SL \i54/i397  (.A(\i54/n5 ),
    .B(\i54/n57 ),
    .Y(\i54/n106 ));
 NAND2xp5_ASAP7_75t_SL \i54/i398  (.A(\i54/n520 ),
    .B(\i54/n54 ),
    .Y(\i54/n147 ));
 NAND2xp5_ASAP7_75t_SL \i54/i399  (.A(\i54/n82 ),
    .B(\i54/n57 ),
    .Y(\i54/n105 ));
 INVx1_ASAP7_75t_SL \i54/i4  (.A(\i54/n32 ),
    .Y(\i54/n4 ));
 NAND3xp33_ASAP7_75t_SL \i54/i40  (.A(\i54/n385 ),
    .B(\i54/n433 ),
    .C(\i54/n419 ),
    .Y(\i54/n475 ));
 NOR2xp33_ASAP7_75t_SL \i54/i400  (.A(\i54/n56 ),
    .B(\i54/n58 ),
    .Y(\i54/n104 ));
 AND2x2_ASAP7_75t_SL \i54/i401  (.A(\i54/n5 ),
    .B(\i54/n76 ),
    .Y(\i54/n146 ));
 NOR2xp67_ASAP7_75t_SL \i54/i402  (.A(\i54/n89 ),
    .B(\i54/n80 ),
    .Y(\i54/n145 ));
 NAND2xp5_ASAP7_75t_SL \i54/i403  (.A(\i54/n85 ),
    .B(\i54/n60 ),
    .Y(\i54/n143 ));
 NOR2xp33_ASAP7_75t_SL \i54/i404  (.A(\i54/n70 ),
    .B(\i54/n83 ),
    .Y(\i54/n141 ));
 NAND2xp5_ASAP7_75t_SL \i54/i405  (.A(\i54/n5 ),
    .B(\i54/n80 ),
    .Y(\i54/n140 ));
 NAND2xp5_ASAP7_75t_SL \i54/i406  (.A(\i54/n78 ),
    .B(\i54/n53 ),
    .Y(\i54/n139 ));
 NAND2xp5_ASAP7_75t_SL \i54/i407  (.A(\i54/n48 ),
    .B(\i54/n74 ),
    .Y(\i54/n103 ));
 AND2x2_ASAP7_75t_SL \i54/i408  (.A(\i54/n5 ),
    .B(\i54/n52 ),
    .Y(\i54/n138 ));
 NOR2xp33_ASAP7_75t_SL \i54/i409  (.A(\i54/n70 ),
    .B(\i54/n57 ),
    .Y(\i54/n102 ));
 NAND2xp5_ASAP7_75t_L \i54/i41  (.A(\i54/n574 ),
    .B(\i54/n465 ),
    .Y(\i54/n474 ));
 NAND2xp5_ASAP7_75t_SL \i54/i410  (.A(\i54/n82 ),
    .B(\i54/n89 ),
    .Y(\i54/n136 ));
 NAND2xp5_ASAP7_75t_SL \i54/i411  (.A(\i54/n82 ),
    .B(\i54/n52 ),
    .Y(\i54/n134 ));
 NAND2xp5_ASAP7_75t_SL \i54/i412  (.A(\i54/n48 ),
    .B(\i54/n52 ),
    .Y(\i54/n131 ));
 NAND2xp33_ASAP7_75t_L \i54/i413  (.A(\i54/n51 ),
    .B(\i54/n73 ),
    .Y(\i54/n101 ));
 NAND2xp5_ASAP7_75t_SL \i54/i414  (.A(\i54/n45 ),
    .B(\i54/n520 ),
    .Y(\i54/n129 ));
 NOR2xp67_ASAP7_75t_L \i54/i415  (.A(\i54/n46 ),
    .B(\i54/n58 ),
    .Y(\i54/n127 ));
 NAND2xp5_ASAP7_75t_SL \i54/i416  (.A(\i54/n50 ),
    .B(\i54/n80 ),
    .Y(\i54/n18 ));
 NAND2xp5_ASAP7_75t_SL \i54/i417  (.A(\i54/n50 ),
    .B(\i54/n83 ),
    .Y(\i54/n126 ));
 AND2x2_ASAP7_75t_SL \i54/i418  (.A(\i54/n520 ),
    .B(\i54/n83 ),
    .Y(\i54/n125 ));
 NAND2xp5_ASAP7_75t_L \i54/i419  (.A(\i54/n13 ),
    .B(\i54/n15 ),
    .Y(\i54/n124 ));
 NAND2xp33_ASAP7_75t_SL \i54/i42  (.A(\i54/n430 ),
    .B(\i54/n447 ),
    .Y(\i54/n473 ));
 AND2x2_ASAP7_75t_SL \i54/i420  (.A(\i54/n520 ),
    .B(\i54/n60 ),
    .Y(\i54/n123 ));
 NOR2xp33_ASAP7_75t_SL \i54/i421  (.A(\i54/n61 ),
    .B(\i54/n47 ),
    .Y(\i54/n100 ));
 NOR2xp33_ASAP7_75t_SL \i54/i422  (.A(\i54/n55 ),
    .B(\i54/n49 ),
    .Y(\i54/n99 ));
 NOR2xp67_ASAP7_75t_SL \i54/i423  (.A(\i54/n54 ),
    .B(\i54/n74 ),
    .Y(\i54/n122 ));
 NAND2xp5_ASAP7_75t_SL \i54/i424  (.A(\i54/n5 ),
    .B(\i54/n83 ),
    .Y(\i54/n98 ));
 NAND2xp5_ASAP7_75t_SL \i54/i425  (.A(\i54/n59 ),
    .B(\i54/n53 ),
    .Y(\i54/n120 ));
 NAND2xp5_ASAP7_75t_SL \i54/i426  (.A(\i54/n78 ),
    .B(\i54/n83 ),
    .Y(\i54/n119 ));
 NAND2xp5_ASAP7_75t_SL \i54/i427  (.A(\i54/n59 ),
    .B(\i54/n80 ),
    .Y(\i54/n97 ));
 NAND2xp5_ASAP7_75t_SL \i54/i428  (.A(\i54/n520 ),
    .B(\i54/n76 ),
    .Y(\i54/n118 ));
 NOR2xp33_ASAP7_75t_SL \i54/i429  (.A(\i54/n94 ),
    .B(\i54/n13 ),
    .Y(\i54/n96 ));
 NOR2x1_ASAP7_75t_SL \i54/i43  (.A(\i54/n446 ),
    .B(\i54/n455 ),
    .Y(\i54/n481 ));
 NOR2xp33_ASAP7_75t_SL \i54/i430  (.A(\i54/n94 ),
    .B(\i54/n56 ),
    .Y(\i54/n95 ));
 NAND2x1_ASAP7_75t_SL \i54/i431  (.A(\i54/n59 ),
    .B(\i54/n86 ),
    .Y(\i54/n116 ));
 NAND2x1_ASAP7_75t_SL \i54/i432  (.A(\i54/n5 ),
    .B(\i54/n53 ),
    .Y(\i54/n16 ));
 INVx2_ASAP7_75t_SL \i54/i433  (.A(\i54/n520 ),
    .Y(\i54/n94 ));
 INVx1_ASAP7_75t_SL \i54/i434  (.A(\i54/n93 ),
    .Y(\i54/n92 ));
 INVx3_ASAP7_75t_SL \i54/i435  (.A(\i54/n91 ),
    .Y(\i54/n90 ));
 INVx3_ASAP7_75t_SL \i54/i436  (.A(\i54/n89 ),
    .Y(\i54/n88 ));
 INVx4_ASAP7_75t_SL \i54/i437  (.A(\i54/n87 ),
    .Y(\i54/n86 ));
 INVx2_ASAP7_75t_SL \i54/i438  (.A(\i54/n85 ),
    .Y(\i54/n84 ));
 INVx2_ASAP7_75t_SL \i54/i439  (.A(\i54/n82 ),
    .Y(\i54/n81 ));
 NAND2xp33_ASAP7_75t_L \i54/i44  (.A(\i54/n435 ),
    .B(\i54/n407 ),
    .Y(\i54/n470 ));
 INVx4_ASAP7_75t_SL \i54/i440  (.A(\i54/n80 ),
    .Y(\i54/n79 ));
 INVx2_ASAP7_75t_SL \i54/i441  (.A(\i54/n78 ),
    .Y(\i54/n77 ));
 INVx3_ASAP7_75t_SL \i54/i442  (.A(\i54/n76 ),
    .Y(\i54/n75 ));
 INVx2_ASAP7_75t_SL \i54/i443  (.A(\i54/n74 ),
    .Y(\i54/n73 ));
 INVx3_ASAP7_75t_SL \i54/i444  (.A(\i54/n72 ),
    .Y(\i54/n71 ));
 INVx3_ASAP7_75t_SL \i54/i445  (.A(\i54/n70 ),
    .Y(\i54/n69 ));
 INVx3_ASAP7_75t_SL \i54/i446  (.A(\i54/n68 ),
    .Y(\i54/n67 ));
 INVx3_ASAP7_75t_SL \i54/i447  (.A(\i54/n66 ),
    .Y(\i54/n65 ));
 AND2x4_ASAP7_75t_SL \i54/i448  (.A(\i54/n41 ),
    .B(\i54/n527 ),
    .Y(\i54/n93 ));
 OR2x4_ASAP7_75t_SL \i54/i449  (.A(\i54/n32 ),
    .B(\i54/n7 ),
    .Y(\i54/n91 ));
 NAND2xp33_ASAP7_75t_L \i54/i45  (.A(\i54/n574 ),
    .B(\i54/n413 ),
    .Y(\i54/n469 ));
 AND2x4_ASAP7_75t_SL \i54/i450  (.A(\i54/n38 ),
    .B(\i54/n3 ),
    .Y(\i54/n89 ));
 OR2x6_ASAP7_75t_SL \i54/i451  (.A(\i54/n37 ),
    .B(\i54/n44 ),
    .Y(\i54/n87 ));
 AND2x4_ASAP7_75t_SL \i54/i452  (.A(\i54/n31 ),
    .B(\i54/n42 ),
    .Y(\i54/n85 ));
 AND2x4_ASAP7_75t_SL \i54/i453  (.A(\i54/n36 ),
    .B(\i54/n39 ),
    .Y(\i54/n83 ));
 NAND2x1_ASAP7_75t_SL \i54/i454  (.A(\i54/n36 ),
    .B(\i54/n39 ),
    .Y(\i54/n15 ));
 AND2x4_ASAP7_75t_SL \i54/i455  (.A(\i54/n31 ),
    .B(\i54/n41 ),
    .Y(\i54/n82 ));
 AND2x4_ASAP7_75t_SL \i54/i456  (.A(\i54/n43 ),
    .B(\i54/n35 ),
    .Y(\i54/n80 ));
 AND2x4_ASAP7_75t_SL \i54/i457  (.A(\i54/n31 ),
    .B(\i54/n526 ),
    .Y(\i54/n78 ));
 AND2x4_ASAP7_75t_SL \i54/i458  (.A(\i54/n36 ),
    .B(\i54/n522 ),
    .Y(\i54/n76 ));
 AND2x4_ASAP7_75t_SL \i54/i459  (.A(\i54/n38 ),
    .B(\i54/n4 ),
    .Y(\i54/n74 ));
 NOR2xp33_ASAP7_75t_SL \i54/i46  (.A(\i54/n412 ),
    .B(\i54/n437 ),
    .Y(\i54/n468 ));
 AND2x4_ASAP7_75t_SL \i54/i460  (.A(\i54/n38 ),
    .B(\i54/n36 ),
    .Y(\i54/n72 ));
 AND2x4_ASAP7_75t_SL \i54/i461  (.A(\i54/n36 ),
    .B(\i54/n35 ),
    .Y(\i54/n70 ));
 AND2x4_ASAP7_75t_SL \i54/i462  (.A(\i54/n41 ),
    .B(\i54/n502 ),
    .Y(\i54/n68 ));
 OR2x6_ASAP7_75t_SL \i54/i463  (.A(\i54/n518 ),
    .B(\i54/n30 ),
    .Y(\i54/n66 ));
 INVx3_ASAP7_75t_SL \i54/i464  (.A(\i54/n64 ),
    .Y(\i54/n63 ));
 INVx2_ASAP7_75t_SL \i54/i465  (.A(\i54/n62 ),
    .Y(\i54/n14 ));
 INVx4_ASAP7_75t_SL \i54/i466  (.A(\i54/n61 ),
    .Y(\i54/n60 ));
 INVx5_ASAP7_75t_SL \i54/i467  (.A(\i54/n59 ),
    .Y(\i54/n58 ));
 INVx4_ASAP7_75t_SL \i54/i468  (.A(\i54/n57 ),
    .Y(\i54/n56 ));
 INVx4_ASAP7_75t_SL \i54/i469  (.A(\i54/n55 ),
    .Y(\i54/n54 ));
 NAND3xp33_ASAP7_75t_SL \i54/i47  (.A(\i54/n402 ),
    .B(\i54/n410 ),
    .C(\i54/n376 ),
    .Y(\i54/n467 ));
 INVx4_ASAP7_75t_SL \i54/i470  (.A(\i54/n53 ),
    .Y(\i54/n13 ));
 INVx2_ASAP7_75t_SL \i54/i471  (.A(\i54/n50 ),
    .Y(\i54/n49 ));
 INVx4_ASAP7_75t_SL \i54/i472  (.A(\i54/n48 ),
    .Y(\i54/n47 ));
 INVx8_ASAP7_75t_SL \i54/i473  (.A(\i54/n46 ),
    .Y(\i54/n45 ));
 AND2x4_ASAP7_75t_SL \i54/i474  (.A(\i54/n41 ),
    .B(\i54/n550 ),
    .Y(\i54/n64 ));
 AND2x4_ASAP7_75t_SL \i54/i475  (.A(\i54/n527 ),
    .B(\i54/n42 ),
    .Y(\i54/n62 ));
 NAND2x1p5_ASAP7_75t_SL \i54/i476  (.A(\i54/n38 ),
    .B(\i54/n43 ),
    .Y(\i54/n61 ));
 AND2x4_ASAP7_75t_SL \i54/i477  (.A(\i54/n526 ),
    .B(\i54/n550 ),
    .Y(\i54/n59 ));
 AND2x4_ASAP7_75t_SL \i54/i478  (.A(\i54/n522 ),
    .B(\i54/n4 ),
    .Y(\i54/n57 ));
 OR2x4_ASAP7_75t_SL \i54/i479  (.A(\i54/n33 ),
    .B(\i54/n34 ),
    .Y(\i54/n55 ));
 NOR2x1_ASAP7_75t_SL \i54/i48  (.A(\i54/n359 ),
    .B(\i54/n421 ),
    .Y(\i54/n466 ));
 AND2x4_ASAP7_75t_SL \i54/i480  (.A(\i54/n35 ),
    .B(\i54/n4 ),
    .Y(\i54/n53 ));
 AND2x4_ASAP7_75t_SL \i54/i481  (.A(\i54/n3 ),
    .B(\i54/n39 ),
    .Y(\i54/n52 ));
 NAND2x1_ASAP7_75t_SL \i54/i482  (.A(\i54/n3 ),
    .B(\i54/n39 ),
    .Y(\i54/n51 ));
 AND2x4_ASAP7_75t_SL \i54/i483  (.A(\i54/n526 ),
    .B(\i54/n502 ),
    .Y(\i54/n50 ));
 AND2x4_ASAP7_75t_SL \i54/i484  (.A(\i54/n42 ),
    .B(\i54/n502 ),
    .Y(\i54/n48 ));
 OR2x6_ASAP7_75t_SL \i54/i485  (.A(\i54/n29 ),
    .B(\i54/n40 ),
    .Y(\i54/n46 ));
 INVx2_ASAP7_75t_SL \i54/i486  (.A(\i54/n43 ),
    .Y(\i54/n44 ));
 INVx2_ASAP7_75t_SL \i54/i487  (.A(\i54/n513 ),
    .Y(\i54/n42 ));
 NAND2xp5_ASAP7_75t_SL \i54/i488  (.A(\i54/n10 ),
    .B(\i54/n0 ),
    .Y(\i54/n40 ));
 AND2x2_ASAP7_75t_SL \i54/i489  (.A(\i54/n10 ),
    .B(\i54/n0 ),
    .Y(\i54/n43 ));
 NOR2xp33_ASAP7_75t_SL \i54/i49  (.A(\i54/n428 ),
    .B(\i54/n340 ),
    .Y(\i54/n465 ));
 AND2x2_ASAP7_75t_SL \i54/i490  (.A(\i54/n27 ),
    .B(\i54/n9 ),
    .Y(\i54/n41 ));
 INVx2_ASAP7_75t_SL \i54/i491  (.A(\i54/n7 ),
    .Y(\i54/n39 ));
 INVx1_ASAP7_75t_SL \i54/i492  (.A(\i54/n522 ),
    .Y(\i54/n37 ));
 INVx2_ASAP7_75t_SL \i54/i493  (.A(\i54/n34 ),
    .Y(\i54/n35 ));
 INVx2_ASAP7_75t_SL \i54/i494  (.A(\i54/n31 ),
    .Y(\i54/n30 ));
 NAND2xp5_ASAP7_75t_SL \i54/i495  (.A(\i54/n28 ),
    .B(\i54/n1 ),
    .Y(\i54/n29 ));
 AND2x2_ASAP7_75t_SL \i54/i496  (.A(n13[0]),
    .B(n13[1]),
    .Y(\i54/n38 ));
 AND2x4_ASAP7_75t_SL \i54/i497  (.A(n13[2]),
    .B(n13[3]),
    .Y(\i54/n36 ));
 NAND2xp5_ASAP7_75t_SL \i54/i498  (.A(\i54/n1 ),
    .B(n13[1]),
    .Y(\i54/n34 ));
 OR2x2_ASAP7_75t_SL \i54/i499  (.A(\i54/n0 ),
    .B(n13[3]),
    .Y(\i54/n33 ));
 INVx2_ASAP7_75t_SL \i54/i5  (.A(\i54/n515 ),
    .Y(\i54/n5 ));
 NAND2xp5_ASAP7_75t_SL \i54/i50  (.A(\i54/n435 ),
    .B(\i54/n431 ),
    .Y(\i54/n464 ));
 NAND2x1_ASAP7_75t_SL \i54/i500  (.A(n13[3]),
    .B(\i54/n0 ),
    .Y(\i54/n32 ));
 AND2x2_ASAP7_75t_SL \i54/i501  (.A(n13[7]),
    .B(n13[6]),
    .Y(\i54/n31 ));
 INVx1_ASAP7_75t_SL \i54/i502  (.A(n13[1]),
    .Y(\i54/n28 ));
 INVx3_ASAP7_75t_SL \i54/i503  (.A(n13[5]),
    .Y(\i54/n27 ));
 INVx2_ASAP7_75t_SL \i54/i504  (.A(n13[6]),
    .Y(\i54/n12 ));
 INVx2_ASAP7_75t_SL \i54/i505  (.A(n13[7]),
    .Y(\i54/n11 ));
 INVx2_ASAP7_75t_SL \i54/i506  (.A(n13[3]),
    .Y(\i54/n10 ));
 INVx2_ASAP7_75t_SL \i54/i507  (.A(n13[4]),
    .Y(\i54/n9 ));
 OR2x2_ASAP7_75t_SL \i54/i508  (.A(\i54/n138 ),
    .B(\i54/n541 ),
    .Y(\i54/n8 ));
 OR2x2_ASAP7_75t_SL \i54/i509  (.A(n13[0]),
    .B(n13[1]),
    .Y(\i54/n7 ));
 NOR2x1_ASAP7_75t_SL \i54/i51  (.A(\i54/n344 ),
    .B(\i54/n437 ),
    .Y(\i54/n463 ));
 AND2x4_ASAP7_75t_SL \i54/i510  (.A(n13[7]),
    .B(\i54/n12 ),
    .Y(\i54/n502 ));
 INVx3_ASAP7_75t_SL \i54/i511  (.A(\i54/n505 ),
    .Y(\i54/n503 ));
 OAI31xp33_ASAP7_75t_SL \i54/i512  (.A1(\i54/n60 ),
    .A2(\i54/n54 ),
    .A3(\i54/n90 ),
    .B(\i54/n505 ),
    .Y(\i54/n504 ));
 AOI21xp5_ASAP7_75t_SL \i54/i513  (.A1(\i54/n74 ),
    .A2(\i54/n505 ),
    .B(\i54/n262 ),
    .Y(\i54/n506 ));
 AOI22xp5_ASAP7_75t_SL \i54/i514  (.A1(\i54/n520 ),
    .A2(\i54/n52 ),
    .B1(\i54/n505 ),
    .B2(\i54/n72 ),
    .Y(\i54/n507 ));
 NAND2xp5_ASAP7_75t_SL \i54/i515  (.A(\i54/n505 ),
    .B(\i54/n70 ),
    .Y(\i54/n508 ));
 NAND2xp5_ASAP7_75t_SL \i54/i516  (.A(\i54/n505 ),
    .B(\i54/n57 ),
    .Y(\i54/n509 ));
 NOR2xp33_ASAP7_75t_SL \i54/i517  (.A(\i54/n505 ),
    .B(\i54/n85 ),
    .Y(\i54/n510 ));
 NAND2xp5_ASAP7_75t_SL \i54/i518  (.A(\i54/n505 ),
    .B(\i54/n80 ),
    .Y(\i54/n511 ));
 NOR2x1_ASAP7_75t_SL \i54/i519  (.A(\i54/n505 ),
    .B(\i54/n82 ),
    .Y(\i54/n512 ));
 NOR2x1_ASAP7_75t_SL \i54/i52  (.A(\i54/n411 ),
    .B(\i54/n422 ),
    .Y(\i54/n462 ));
 NAND2xp5_ASAP7_75t_SL \i54/i520  (.A(\i54/n9 ),
    .B(n13[5]),
    .Y(\i54/n513 ));
 OAI221xp5_ASAP7_75t_SL \i54/i521  (.A1(\i54/n122 ),
    .A2(\i54/n92 ),
    .B1(\i54/n122 ),
    .B2(\i54/n515 ),
    .C(\i54/n307 ),
    .Y(\i54/n516 ));
 OR2x2_ASAP7_75t_SL \i54/i522  (.A(\i54/n514 ),
    .B(\i54/n513 ),
    .Y(\i54/n515 ));
 NAND2xp5_ASAP7_75t_SL \i54/i523  (.A(\i54/n11 ),
    .B(n13[6]),
    .Y(\i54/n514 ));
 NAND2xp5_ASAP7_75t_SL \i54/i524  (.A(\i54/n66 ),
    .B(\i54/n515 ),
    .Y(\i54/n517 ));
 NAND2x1p5_ASAP7_75t_SL \i54/i525  (.A(n13[4]),
    .B(n13[5]),
    .Y(\i54/n518 ));
 AND2x4_ASAP7_75t_SL \i54/i526  (.A(\i54/n519 ),
    .B(\i54/n502 ),
    .Y(\i54/n505 ));
 AND2x4_ASAP7_75t_SL \i54/i527  (.A(\i54/n527 ),
    .B(\i54/n519 ),
    .Y(\i54/n520 ));
 OA21x2_ASAP7_75t_SL \i54/i528  (.A1(\i54/n542 ),
    .A2(\i54/n55 ),
    .B(\i54/n19 ),
    .Y(\i54/n521 ));
 AND2x4_ASAP7_75t_SL \i54/i529  (.A(n13[0]),
    .B(\i54/n28 ),
    .Y(\i54/n522 ));
 NAND2xp5_ASAP7_75t_SL \i54/i53  (.A(\i54/n553 ),
    .B(\i54/n416 ),
    .Y(\i54/n461 ));
 OAI21xp33_ASAP7_75t_SL \i54/i530  (.A1(\i54/n515 ),
    .A2(\i54/n523 ),
    .B(\i54/n131 ),
    .Y(\i54/n524 ));
 NAND2xp33_ASAP7_75t_SL \i54/i531  (.A(\i54/n61 ),
    .B(\i54/n523 ),
    .Y(\i54/n525 ));
 AND2x2_ASAP7_75t_SL \i54/i532  (.A(n13[4]),
    .B(\i54/n27 ),
    .Y(\i54/n526 ));
 AND2x2_ASAP7_75t_SL \i54/i533  (.A(\i54/n11 ),
    .B(\i54/n12 ),
    .Y(\i54/n527 ));
 INVx3_ASAP7_75t_SL \i54/i534  (.A(\i54/n528 ),
    .Y(\i54/n529 ));
 AND2x4_ASAP7_75t_SL \i54/i535  (.A(\i54/n526 ),
    .B(\i54/n527 ),
    .Y(\i54/n528 ));
 AOI21xp5_ASAP7_75t_SL \i54/i536  (.A1(\i54/n53 ),
    .A2(\i54/n528 ),
    .B(\i54/n273 ),
    .Y(\i54/n530 ));
 OAI21xp5_ASAP7_75t_SL \i54/i537  (.A1(\i54/n528 ),
    .A2(\i54/n165 ),
    .B(\i54/n72 ),
    .Y(\i54/n531 ));
 AOI22xp5_ASAP7_75t_SL \i54/i538  (.A1(\i54/n86 ),
    .A2(\i54/n161 ),
    .B1(\i54/n528 ),
    .B2(\i54/n89 ),
    .Y(\i54/n532 ));
 AOI222xp33_ASAP7_75t_SL \i54/i539  (.A1(\i54/n76 ),
    .A2(\i54/n62 ),
    .B1(\i54/n5 ),
    .B2(\i54/n45 ),
    .C1(\i54/n72 ),
    .C2(\i54/n528 ),
    .Y(\i54/n533 ));
 NOR5xp2_ASAP7_75t_SL \i54/i54  (.A(\i54/n302 ),
    .B(\i54/n547 ),
    .C(\i54/n315 ),
    .D(\i54/n25 ),
    .E(\i54/n280 ),
    .Y(\i54/n460 ));
 AOI22xp5_ASAP7_75t_SL \i54/i540  (.A1(\i54/n528 ),
    .A2(\i54/n60 ),
    .B1(\i54/n78 ),
    .B2(\i54/n57 ),
    .Y(\i54/n534 ));
 NAND2xp5_ASAP7_75t_SL \i54/i541  (.A(\i54/n57 ),
    .B(\i54/n528 ),
    .Y(\i54/n535 ));
 NAND2xp5_ASAP7_75t_SL \i54/i542  (.A(\i54/n528 ),
    .B(\i54/n70 ),
    .Y(\i54/n536 ));
 NAND2xp5_ASAP7_75t_SL \i54/i543  (.A(\i54/n60 ),
    .B(\i54/n528 ),
    .Y(\i54/n537 ));
 NOR2xp67_ASAP7_75t_SL \i54/i544  (.A(\i54/n542 ),
    .B(\i54/n87 ),
    .Y(\i54/n538 ));
 OAI22xp5_ASAP7_75t_SL \i54/i545  (.A1(\i54/n542 ),
    .A2(\i54/n51 ),
    .B1(\i54/n55 ),
    .B2(\i54/n49 ),
    .Y(\i54/n539 ));
 OAI22xp5_ASAP7_75t_SL \i54/i546  (.A1(\i54/n542 ),
    .A2(\i54/n61 ),
    .B1(\i54/n66 ),
    .B2(\i54/n73 ),
    .Y(\i54/n540 ));
 OAI22xp5_ASAP7_75t_SL \i54/i547  (.A1(\i54/n542 ),
    .A2(\i54/n79 ),
    .B1(\i54/n66 ),
    .B2(\i54/n55 ),
    .Y(\i54/n541 ));
 OAI22xp33_ASAP7_75t_SL \i54/i548  (.A1(\i54/n51 ),
    .A2(\i54/n529 ),
    .B1(\i54/n13 ),
    .B2(\i54/n542 ),
    .Y(\i54/n543 ));
 OAI22xp5_ASAP7_75t_SL \i54/i549  (.A1(\i54/n91 ),
    .A2(\i54/n542 ),
    .B1(\i54/n49 ),
    .B2(\i54/n13 ),
    .Y(\i54/n544 ));
 NOR2x1_ASAP7_75t_SL \i54/i55  (.A(\i54/n2 ),
    .B(\i54/n423 ),
    .Y(\i54/n459 ));
 AOI31xp33_ASAP7_75t_SL \i54/i550  (.A1(\i54/n542 ),
    .A2(\i54/n81 ),
    .A3(\i54/n67 ),
    .B(\i54/n55 ),
    .Y(\i54/n545 ));
 OAI222xp33_ASAP7_75t_SL \i54/i551  (.A1(\i54/n523 ),
    .A2(\i54/n542 ),
    .B1(\i54/n56 ),
    .B2(\i54/n66 ),
    .C1(\i54/n69 ),
    .C2(\i54/n77 ),
    .Y(\i54/n546 ));
 OAI221xp5_ASAP7_75t_SL \i54/i552  (.A1(\i54/n56 ),
    .A2(\i54/n63 ),
    .B1(\i54/n542 ),
    .B2(\i54/n55 ),
    .C(\i54/n19 ),
    .Y(\i54/n547 ));
 OAI21xp5_ASAP7_75t_SL \i54/i553  (.A1(\i54/n542 ),
    .A2(\i54/n145 ),
    .B(\i54/n192 ),
    .Y(\i54/n548 ));
 AOI31xp33_ASAP7_75t_SL \i54/i554  (.A1(\i54/n542 ),
    .A2(\i54/n14 ),
    .A3(\i54/n503 ),
    .B(\i54/n46 ),
    .Y(\i54/n549 ));
 INVx2_ASAP7_75t_SL \i54/i555  (.A(\i54/n518 ),
    .Y(\i54/n519 ));
 AND2x2_ASAP7_75t_SL \i54/i556  (.A(n13[6]),
    .B(\i54/n11 ),
    .Y(\i54/n550 ));
 INVx4_ASAP7_75t_SL \i54/i557  (.A(\i54/n551 ),
    .Y(\i54/n542 ));
 AND2x4_ASAP7_75t_SL \i54/i558  (.A(\i54/n519 ),
    .B(\i54/n550 ),
    .Y(\i54/n551 ));
 AO22x2_ASAP7_75t_SL \i54/i559  (.A1(\i54/n93 ),
    .A2(\i54/n90 ),
    .B1(\i54/n551 ),
    .B2(\i54/n83 ),
    .Y(\i54/n552 ));
 NAND2x1_ASAP7_75t_SL \i54/i56  (.A(\i54/n420 ),
    .B(\i54/n400 ),
    .Y(\i54/n472 ));
 AOI211xp5_ASAP7_75t_SL \i54/i560  (.A1(\i54/n124 ),
    .A2(\i54/n551 ),
    .B(\i54/n323 ),
    .C(\i54/n256 ),
    .Y(\i54/n553 ));
 NAND2xp5_ASAP7_75t_SL \i54/i561  (.A(\i54/n45 ),
    .B(\i54/n551 ),
    .Y(\i54/n554 ));
 NAND2xp5_ASAP7_75t_SL \i54/i562  (.A(\i54/n551 ),
    .B(\i54/n70 ),
    .Y(\i54/n555 ));
 AND2x2_ASAP7_75t_SL \i54/i563  (.A(\i54/n551 ),
    .B(\i54/n74 ),
    .Y(\i54/n556 ));
 NAND2xp5_ASAP7_75t_SL \i54/i564  (.A(\i54/n551 ),
    .B(\i54/n57 ),
    .Y(\i54/n557 ));
 NAND2x1p5_ASAP7_75t_SL \i54/i565  (.A(\i54/n3 ),
    .B(\i54/n522 ),
    .Y(\i54/n523 ));
 NAND2xp5_ASAP7_75t_SL \i54/i566  (.A(\i54/n6 ),
    .B(\i54/n528 ),
    .Y(\i54/n558 ));
 AND2x2_ASAP7_75t_SL \i54/i567  (.A(\i54/n62 ),
    .B(\i54/n6 ),
    .Y(\i54/n559 ));
 NAND2xp5_ASAP7_75t_SL \i54/i568  (.A(\i54/n65 ),
    .B(\i54/n6 ),
    .Y(\i54/n560 ));
 NAND2xp5_ASAP7_75t_SL \i54/i569  (.A(\i54/n64 ),
    .B(\i54/n6 ),
    .Y(\i54/n561 ));
 NOR2x1_ASAP7_75t_SL \i54/i57  (.A(\i54/n438 ),
    .B(\i54/n422 ),
    .Y(\i54/n458 ));
 NAND2xp5_ASAP7_75t_SL \i54/i570  (.A(\i54/n520 ),
    .B(\i54/n6 ),
    .Y(\i54/n562 ));
 OAI31xp33_ASAP7_75t_SL \i54/i571  (.A1(\i54/n72 ),
    .A2(\i54/n6 ),
    .A3(\i54/n53 ),
    .B(\i54/n50 ),
    .Y(\i54/n563 ));
 AOI22xp5_ASAP7_75t_SL \i54/i572  (.A1(\i54/n82 ),
    .A2(\i54/n60 ),
    .B1(\i54/n50 ),
    .B2(\i54/n6 ),
    .Y(\i54/n564 ));
 NOR2xp33_ASAP7_75t_SL \i54/i573  (.A(\i54/n89 ),
    .B(\i54/n6 ),
    .Y(\i54/n565 ));
 NAND2xp5_ASAP7_75t_SL \i54/i574  (.A(\i54/n85 ),
    .B(\i54/n6 ),
    .Y(\i54/n566 ));
 AOI22xp5_ASAP7_75t_SL \i54/i575  (.A1(\i54/n520 ),
    .A2(\i54/n80 ),
    .B1(\i54/n78 ),
    .B2(\i54/n6 ),
    .Y(\i54/n567 ));
 NAND2xp5_ASAP7_75t_SL \i54/i576  (.A(\i54/n6 ),
    .B(\i54/n59 ),
    .Y(\i54/n568 ));
 AO21x2_ASAP7_75t_SL \i54/i577  (.A1(\i54/n82 ),
    .A2(\i54/n6 ),
    .B(\i54/n213 ),
    .Y(\i54/n569 ));
 NAND2xp33_ASAP7_75t_L \i54/i578  (.A(\i54/n6 ),
    .B(\i54/n78 ),
    .Y(\i54/n570 ));
 AOI22xp33_ASAP7_75t_SL \i54/i579  (.A1(\i54/n93 ),
    .A2(\i54/n54 ),
    .B1(\i54/n64 ),
    .B2(\i54/n6 ),
    .Y(\i54/n571 ));
 NOR2x1_ASAP7_75t_SL \i54/i58  (.A(\i54/n358 ),
    .B(\i54/n421 ),
    .Y(\i54/n471 ));
 NAND2xp5_ASAP7_75t_SL \i54/i580  (.A(\i54/n48 ),
    .B(\i54/n6 ),
    .Y(\i54/n572 ));
 AND4x1_ASAP7_75t_SL \i54/i581  (.A(\i54/n533 ),
    .B(\i54/n342 ),
    .C(\i54/n575 ),
    .D(\i54/n275 ),
    .Y(\i54/n573 ));
 AND4x1_ASAP7_75t_SL \i54/i582  (.A(\i54/n291 ),
    .B(\i54/n506 ),
    .C(\i54/n532 ),
    .D(\i54/n533 ),
    .Y(\i54/n574 ));
 AOI21xp5_ASAP7_75t_SL \i54/i583  (.A1(\i54/n551 ),
    .A2(\i54/n72 ),
    .B(\i54/n539 ),
    .Y(\i54/n575 ));
 AND2x2_ASAP7_75t_SL \i54/i584  (.A(\i54/n576 ),
    .B(\i54/n434 ),
    .Y(\i54/n577 ));
 AOI21xp33_ASAP7_75t_SL \i54/i585  (.A1(\i54/n45 ),
    .A2(\i54/n68 ),
    .B(\i54/n125 ),
    .Y(\i54/n576 ));
 NAND3xp33_ASAP7_75t_SL \i54/i586  (.A(\i54/n578 ),
    .B(\i54/n268 ),
    .C(\i54/n334 ),
    .Y(\i54/n579 ));
 AO21x1_ASAP7_75t_SL \i54/i587  (.A1(\i54/n63 ),
    .A2(\i54/n542 ),
    .B(\i54/n88 ),
    .Y(\i54/n578 ));
 NOR3xp33_ASAP7_75t_SL \i54/i588  (.A(\i54/n580 ),
    .B(\i54/n548 ),
    .C(\i54/n213 ),
    .Y(\i54/n581 ));
 OAI21xp5_ASAP7_75t_SL \i54/i589  (.A1(\i54/n66 ),
    .A2(\i54/n15 ),
    .B(\i54/n568 ),
    .Y(\i54/n580 ));
 INVxp67_ASAP7_75t_SL \i54/i59  (.A(\i54/n456 ),
    .Y(\i54/n457 ));
 INVx2_ASAP7_75t_SL \i54/i6  (.A(\i54/n523 ),
    .Y(\i54/n6 ));
 INVxp67_ASAP7_75t_SL \i54/i60  (.A(\i54/n452 ),
    .Y(\i54/n453 ));
 AND5x1_ASAP7_75t_SL \i54/i61  (.A(\i54/n372 ),
    .B(\i54/n575 ),
    .C(\i54/n364 ),
    .D(\i54/n289 ),
    .E(\i54/n261 ),
    .Y(\i54/n451 ));
 NOR3xp33_ASAP7_75t_SL \i54/i62  (.A(\i54/n382 ),
    .B(\i54/n363 ),
    .C(\i54/n345 ),
    .Y(\i54/n450 ));
 NOR3xp33_ASAP7_75t_SL \i54/i63  (.A(\i54/n408 ),
    .B(\i54/n346 ),
    .C(\i54/n300 ),
    .Y(\i54/n449 ));
 AND5x1_ASAP7_75t_SL \i54/i64  (.A(\i54/n336 ),
    .B(\i54/n349 ),
    .C(\i54/n331 ),
    .D(\i54/n339 ),
    .E(\i54/n270 ),
    .Y(\i54/n448 ));
 NOR2xp33_ASAP7_75t_SL \i54/i65  (.A(\i54/n409 ),
    .B(\i54/n414 ),
    .Y(\i54/n447 ));
 NAND4xp25_ASAP7_75t_SL \i54/i66  (.A(\i54/n391 ),
    .B(\i54/n399 ),
    .C(\i54/n404 ),
    .D(\i54/n387 ),
    .Y(\i54/n446 ));
 NAND5xp2_ASAP7_75t_SL \i54/i67  (.A(\i54/n371 ),
    .B(\i54/n330 ),
    .C(\i54/n230 ),
    .D(\i54/n216 ),
    .E(\i54/n311 ),
    .Y(\i54/n445 ));
 NOR4xp25_ASAP7_75t_SL \i54/i68  (.A(\i54/n361 ),
    .B(\i54/n547 ),
    .C(\i54/n316 ),
    .D(\i54/n293 ),
    .Y(\i54/n444 ));
 NAND4xp25_ASAP7_75t_SL \i54/i69  (.A(\i54/n379 ),
    .B(\i54/n393 ),
    .C(\i54/n396 ),
    .D(\i54/n398 ),
    .Y(\i54/n443 ));
 NOR2x1p5_ASAP7_75t_SL \i54/i7  (.A(\i54/n497 ),
    .B(\i54/n496 ),
    .Y(n12[4]));
 NAND4xp25_ASAP7_75t_SL \i54/i70  (.A(\i54/n406 ),
    .B(\i54/n404 ),
    .C(\i54/n521 ),
    .D(\i54/n260 ),
    .Y(\i54/n442 ));
 NAND3xp33_ASAP7_75t_SL \i54/i71  (.A(\i54/n398 ),
    .B(\i54/n370 ),
    .C(\i54/n18 ),
    .Y(\i54/n456 ));
 NAND4xp75_ASAP7_75t_SL \i54/i72  (.A(\i54/n307 ),
    .B(\i54/n279 ),
    .C(\i54/n357 ),
    .D(\i54/n21 ),
    .Y(\i54/n455 ));
 NAND2xp33_ASAP7_75t_L \i54/i73  (.A(\i54/n378 ),
    .B(\i54/n439 ),
    .Y(\i54/n441 ));
 AND2x2_ASAP7_75t_SL \i54/i74  (.A(\i54/n381 ),
    .B(\i54/n429 ),
    .Y(\i54/n454 ));
 NAND2x1p5_ASAP7_75t_SL \i54/i75  (.A(\i54/n436 ),
    .B(\i54/n392 ),
    .Y(\i54/n452 ));
 INVx1_ASAP7_75t_L \i54/i76  (.A(\i54/n439 ),
    .Y(\i54/n440 ));
 NOR5xp2_ASAP7_75t_SL \i54/i77  (.A(\i54/n325 ),
    .B(\i54/n299 ),
    .C(\i54/n222 ),
    .D(\i54/n188 ),
    .E(\i54/n99 ),
    .Y(\i54/n432 ));
 NOR3xp33_ASAP7_75t_SL \i54/i78  (.A(\i54/n403 ),
    .B(\i54/n320 ),
    .C(\i54/n314 ),
    .Y(\i54/n431 ));
 NOR2xp33_ASAP7_75t_SL \i54/i79  (.A(\i54/n360 ),
    .B(\i54/n380 ),
    .Y(\i54/n430 ));
 NOR2x2_ASAP7_75t_SL \i54/i8  (.A(\i54/n492 ),
    .B(\i54/n498 ),
    .Y(n12[3]));
 NOR2xp33_ASAP7_75t_SL \i54/i80  (.A(\i54/n401 ),
    .B(\i54/n351 ),
    .Y(\i54/n429 ));
 NOR2x1_ASAP7_75t_SL \i54/i81  (.A(\i54/n365 ),
    .B(\i54/n337 ),
    .Y(\i54/n439 ));
 NAND3xp33_ASAP7_75t_SL \i54/i82  (.A(\i54/n310 ),
    .B(\i54/n563 ),
    .C(\i54/n224 ),
    .Y(\i54/n428 ));
 NAND2xp5_ASAP7_75t_L \i54/i83  (.A(\i54/n400 ),
    .B(\i54/n369 ),
    .Y(\i54/n427 ));
 NAND2xp5_ASAP7_75t_SL \i54/i84  (.A(\i54/n350 ),
    .B(\i54/n390 ),
    .Y(\i54/n426 ));
 NAND3xp33_ASAP7_75t_SL \i54/i85  (.A(\i54/n575 ),
    .B(\i54/n294 ),
    .C(\i54/n275 ),
    .Y(\i54/n438 ));
 NOR3xp33_ASAP7_75t_SL \i54/i86  (.A(\i54/n516 ),
    .B(\i54/n8 ),
    .C(\i54/n277 ),
    .Y(\i54/n425 ));
 NAND2xp5_ASAP7_75t_SL \i54/i87  (.A(\i54/n511 ),
    .B(\i54/n379 ),
    .Y(\i54/n437 ));
 OR3x1_ASAP7_75t_SL \i54/i88  (.A(\i54/n302 ),
    .B(\i54/n315 ),
    .C(\i54/n25 ),
    .Y(\i54/n424 ));
 NOR2x1_ASAP7_75t_SL \i54/i89  (.A(\i54/n314 ),
    .B(\i54/n403 ),
    .Y(\i54/n436 ));
 AND5x2_ASAP7_75t_SL \i54/i9  (.A(\i54/n490 ),
    .B(\i54/n481 ),
    .C(\i54/n483 ),
    .D(\i54/n468 ),
    .E(\i54/n460 ),
    .Y(n12[6]));
 NOR2xp33_ASAP7_75t_SL \i54/i90  (.A(\i54/n362 ),
    .B(\i54/n348 ),
    .Y(\i54/n435 ));
 NOR2xp67_ASAP7_75t_L \i54/i91  (.A(\i54/n303 ),
    .B(\i54/n389 ),
    .Y(\i54/n434 ));
 NOR3x1_ASAP7_75t_SL \i54/i92  (.A(\i54/n309 ),
    .B(\i54/n200 ),
    .C(\i54/n354 ),
    .Y(\i54/n433 ));
 NOR3xp33_ASAP7_75t_SL \i54/i93  (.A(\i54/n317 ),
    .B(\i54/n229 ),
    .C(\i54/n306 ),
    .Y(\i54/n420 ));
 NOR2xp33_ASAP7_75t_SL \i54/i94  (.A(\i54/n579 ),
    .B(\i54/n375 ),
    .Y(\i54/n419 ));
 NAND3xp33_ASAP7_75t_SL \i54/i95  (.A(\i54/n533 ),
    .B(\i54/n367 ),
    .C(\i54/n532 ),
    .Y(\i54/n418 ));
 NAND4xp25_ASAP7_75t_SL \i54/i96  (.A(\i54/n284 ),
    .B(\i54/n298 ),
    .C(\i54/n326 ),
    .D(\i54/n504 ),
    .Y(\i54/n417 ));
 NAND2x1_ASAP7_75t_SL \i54/i97  (.A(\i54/n388 ),
    .B(\i54/n402 ),
    .Y(\i54/n423 ));
 NOR5xp2_ASAP7_75t_SL \i54/i98  (.A(\i54/n397 ),
    .B(\i54/n318 ),
    .C(\i54/n137 ),
    .D(\i54/n244 ),
    .E(\i54/n171 ),
    .Y(\i54/n416 ));
 NAND3xp33_ASAP7_75t_SL \i54/i99  (.A(\i54/n353 ),
    .B(\i54/n373 ),
    .C(\i54/n232 ),
    .Y(\i54/n415 ));
 OAI22xp5_ASAP7_75t_SL i540 (.A1(n277),
    .A2(n477),
    .B1(n1152),
    .B2(n478),
    .Y(n932));
 OAI22xp5_ASAP7_75t_SL i541 (.A1(n564),
    .A2(n483),
    .B1(n563),
    .B2(n482),
    .Y(n931));
 AOI22xp5_ASAP7_75t_SL i542 (.A1(n499),
    .A2(n575),
    .B1(n576),
    .B2(n500),
    .Y(n930));
 OAI22xp5_ASAP7_75t_SL i543 (.A1(n235),
    .A2(n481),
    .B1(n1151),
    .B2(n480),
    .Y(n929));
 OAI22xp5_ASAP7_75t_SL i544 (.A1(n574),
    .A2(n789),
    .B1(n573),
    .B2(n1176),
    .Y(n928));
 OAI22xp5_ASAP7_75t_SL i545 (.A1(n577),
    .A2(n491),
    .B1(n490),
    .B2(n1230),
    .Y(n927));
 XNOR2xp5_ASAP7_75t_SL i546 (.A(n348),
    .B(n503),
    .Y(n926));
 OAI22xp5_ASAP7_75t_SL i547 (.A1(n1231),
    .A2(n510),
    .B1(n511),
    .B2(n581),
    .Y(n925));
 AOI22xp5_ASAP7_75t_SL i548 (.A1(n488),
    .A2(n765),
    .B1(n489),
    .B2(n764),
    .Y(n924));
 AOI22xp5_ASAP7_75t_SL i549 (.A1(n783),
    .A2(n757),
    .B1(n784),
    .B2(n756),
    .Y(n923));
 INVx2_ASAP7_75t_SL \i55/i0  (.A(n11[7]),
    .Y(\i55/n0 ));
 INVx2_ASAP7_75t_SL \i55/i1  (.A(n11[2]),
    .Y(\i55/n1 ));
 NOR2x1p5_ASAP7_75t_SL \i55/i10  (.A(\i55/n487 ),
    .B(\i55/n478 ),
    .Y(n10[5]));
 NAND5xp2_ASAP7_75t_SL \i55/i100  (.A(\i55/n267 ),
    .B(\i55/n340 ),
    .C(\i55/n199 ),
    .D(\i55/n554 ),
    .E(\i55/n251 ),
    .Y(\i55/n400 ));
 NAND3xp33_ASAP7_75t_L \i55/i101  (.A(\i55/n260 ),
    .B(\i55/n294 ),
    .C(\i55/n364 ),
    .Y(\i55/n399 ));
 NOR5xp2_ASAP7_75t_SL \i55/i102  (.A(\i55/n258 ),
    .B(\i55/n106 ),
    .C(\i55/n249 ),
    .D(\i55/n273 ),
    .E(\i55/n90 ),
    .Y(\i55/n398 ));
 NAND4xp25_ASAP7_75t_SL \i55/i103  (.A(\i55/n202 ),
    .B(\i55/n215 ),
    .C(\i55/n314 ),
    .D(\i55/n17 ),
    .Y(\i55/n397 ));
 NOR5xp2_ASAP7_75t_SL \i55/i104  (.A(\i55/n221 ),
    .B(\i55/n263 ),
    .C(\i55/n207 ),
    .D(\i55/n173 ),
    .E(\i55/n171 ),
    .Y(\i55/n396 ));
 NOR2xp33_ASAP7_75t_SL \i55/i105  (.A(\i55/n355 ),
    .B(\i55/n390 ),
    .Y(\i55/n395 ));
 NOR2xp33_ASAP7_75t_SL \i55/i106  (.A(\i55/n345 ),
    .B(\i55/n374 ),
    .Y(\i55/n394 ));
 NAND3x1_ASAP7_75t_SL \i55/i107  (.A(\i55/n219 ),
    .B(\i55/n372 ),
    .C(\i55/n340 ),
    .Y(\i55/n410 ));
 NAND3x1_ASAP7_75t_SL \i55/i108  (.A(\i55/n335 ),
    .B(\i55/n315 ),
    .C(\i55/n282 ),
    .Y(\i55/n409 ));
 AOI21xp5_ASAP7_75t_L \i55/i109  (.A1(\i55/n499 ),
    .A2(\i55/n558 ),
    .B(\i55/n151 ),
    .Y(\i55/n386 ));
 AND2x4_ASAP7_75t_SL \i55/i11  (.A(\i55/n488 ),
    .B(\i55/n471 ),
    .Y(n10[0]));
 NOR2xp33_ASAP7_75t_SL \i55/i110  (.A(\i55/n286 ),
    .B(\i55/n325 ),
    .Y(\i55/n385 ));
 NAND2xp5_ASAP7_75t_SL \i55/i111  (.A(\i55/n313 ),
    .B(\i55/n344 ),
    .Y(\i55/n384 ));
 NOR2xp33_ASAP7_75t_SL \i55/i112  (.A(\i55/n343 ),
    .B(\i55/n530 ),
    .Y(\i55/n383 ));
 NOR2xp33_ASAP7_75t_SL \i55/i113  (.A(\i55/n320 ),
    .B(\i55/n330 ),
    .Y(\i55/n382 ));
 NOR2xp67_ASAP7_75t_SL \i55/i114  (.A(\i55/n159 ),
    .B(\i55/n327 ),
    .Y(\i55/n381 ));
 NOR2xp33_ASAP7_75t_SL \i55/i115  (.A(\i55/n22 ),
    .B(\i55/n325 ),
    .Y(\i55/n380 ));
 NOR4xp25_ASAP7_75t_SL \i55/i116  (.A(\i55/n298 ),
    .B(\i55/n24 ),
    .C(\i55/n22 ),
    .D(\i55/n168 ),
    .Y(\i55/n379 ));
 NAND2xp5_ASAP7_75t_SL \i55/i117  (.A(\i55/n245 ),
    .B(\i55/n306 ),
    .Y(\i55/n378 ));
 NOR4xp25_ASAP7_75t_SL \i55/i118  (.A(\i55/n103 ),
    .B(\i55/n237 ),
    .C(\i55/n209 ),
    .D(\i55/n223 ),
    .Y(\i55/n377 ));
 NOR3xp33_ASAP7_75t_SL \i55/i119  (.A(\i55/n242 ),
    .B(\i55/n201 ),
    .C(\i55/n241 ),
    .Y(\i55/n376 ));
 NOR3xp33_ASAP7_75t_SL \i55/i12  (.A(\i55/n460 ),
    .B(\i55/n456 ),
    .C(\i55/n463 ),
    .Y(\i55/n488 ));
 NAND2xp5_ASAP7_75t_SL \i55/i120  (.A(\i55/n277 ),
    .B(\i55/n332 ),
    .Y(\i55/n375 ));
 NAND2xp5_ASAP7_75t_SL \i55/i121  (.A(\i55/n293 ),
    .B(\i55/n23 ),
    .Y(\i55/n374 ));
 NOR2xp33_ASAP7_75t_SL \i55/i122  (.A(\i55/n286 ),
    .B(\i55/n288 ),
    .Y(\i55/n373 ));
 NOR2x1p5_ASAP7_75t_SL \i55/i123  (.A(\i55/n268 ),
    .B(\i55/n502 ),
    .Y(\i55/n372 ));
 NAND2xp33_ASAP7_75t_SL \i55/i124  (.A(\i55/n342 ),
    .B(\i55/n323 ),
    .Y(\i55/n371 ));
 NAND3xp33_ASAP7_75t_SL \i55/i125  (.A(\i55/n25 ),
    .B(\i55/n540 ),
    .C(\i55/n496 ),
    .Y(\i55/n370 ));
 NOR3xp33_ASAP7_75t_SL \i55/i126  (.A(\i55/n203 ),
    .B(\i55/n216 ),
    .C(\i55/n186 ),
    .Y(\i55/n393 ));
 NAND2xp5_ASAP7_75t_SL \i55/i127  (.A(\i55/n297 ),
    .B(\i55/n202 ),
    .Y(\i55/n392 ));
 NOR2x1_ASAP7_75t_SL \i55/i128  (.A(\i55/n266 ),
    .B(\i55/n291 ),
    .Y(\i55/n391 ));
 NAND2xp67_ASAP7_75t_SL \i55/i129  (.A(\i55/n199 ),
    .B(\i55/n299 ),
    .Y(\i55/n390 ));
 NOR2x2_ASAP7_75t_SL \i55/i13  (.A(\i55/n480 ),
    .B(\i55/n481 ),
    .Y(n10[2]));
 NOR2x1_ASAP7_75t_SL \i55/i130  (.A(\i55/n269 ),
    .B(\i55/n328 ),
    .Y(\i55/n389 ));
 NAND2xp33_ASAP7_75t_SL \i55/i131  (.A(\i55/n556 ),
    .B(\i55/n287 ),
    .Y(\i55/n369 ));
 NOR2x1_ASAP7_75t_SL \i55/i132  (.A(\i55/n24 ),
    .B(\i55/n286 ),
    .Y(\i55/n388 ));
 NOR3x1_ASAP7_75t_SL \i55/i133  (.A(\i55/n207 ),
    .B(\i55/n196 ),
    .C(\i55/n170 ),
    .Y(\i55/n387 ));
 INVx1_ASAP7_75t_SL \i55/i134  (.A(\i55/n366 ),
    .Y(\i55/n367 ));
 INVx1_ASAP7_75t_SL \i55/i135  (.A(\i55/n27 ),
    .Y(\i55/n365 ));
 NOR4xp25_ASAP7_75t_SL \i55/i136  (.A(\i55/n190 ),
    .B(\i55/n226 ),
    .C(\i55/n214 ),
    .D(\i55/n182 ),
    .Y(\i55/n364 ));
 AOI211xp5_ASAP7_75t_SL \i55/i137  (.A1(\i55/n109 ),
    .A2(\i55/n53 ),
    .B(\i55/n309 ),
    .C(\i55/n240 ),
    .Y(\i55/n363 ));
 NAND2xp33_ASAP7_75t_SL \i55/i138  (.A(\i55/n283 ),
    .B(\i55/n308 ),
    .Y(\i55/n362 ));
 NAND5xp2_ASAP7_75t_SL \i55/i139  (.A(\i55/n224 ),
    .B(\i55/n236 ),
    .C(\i55/n247 ),
    .D(\i55/n166 ),
    .E(\i55/n104 ),
    .Y(\i55/n361 ));
 NAND4xp75_ASAP7_75t_SL \i55/i14  (.A(\i55/n446 ),
    .B(\i55/n466 ),
    .C(\i55/n444 ),
    .D(\i55/n572 ),
    .Y(\i55/n487 ));
 OAI221xp5_ASAP7_75t_SL \i55/i140  (.A1(\i55/n107 ),
    .A2(\i55/n83 ),
    .B1(\i55/n107 ),
    .B2(\i55/n14 ),
    .C(\i55/n293 ),
    .Y(\i55/n360 ));
 NOR2xp33_ASAP7_75t_SL \i55/i141  (.A(\i55/n274 ),
    .B(\i55/n278 ),
    .Y(\i55/n359 ));
 AOI211xp5_ASAP7_75t_SL \i55/i142  (.A1(\i55/n155 ),
    .A2(\i55/n529 ),
    .B(\i55/n257 ),
    .C(\i55/n174 ),
    .Y(\i55/n358 ));
 OA21x2_ASAP7_75t_SL \i55/i143  (.A1(\i55/n537 ),
    .A2(\i55/n499 ),
    .B(\i55/n341 ),
    .Y(\i55/n357 ));
 NOR4xp25_ASAP7_75t_SL \i55/i144  (.A(\i55/n250 ),
    .B(\i55/n163 ),
    .C(\i55/n195 ),
    .D(\i55/n170 ),
    .Y(\i55/n356 ));
 NAND5xp2_ASAP7_75t_SL \i55/i145  (.A(\i55/n137 ),
    .B(\i55/n94 ),
    .C(\i55/n145 ),
    .D(\i55/n561 ),
    .E(\i55/n88 ),
    .Y(\i55/n355 ));
 NOR3xp33_ASAP7_75t_SL \i55/i146  (.A(\i55/n292 ),
    .B(\i55/n165 ),
    .C(\i55/n87 ),
    .Y(\i55/n354 ));
 NAND5xp2_ASAP7_75t_SL \i55/i147  (.A(\i55/n197 ),
    .B(\i55/n99 ),
    .C(\i55/n539 ),
    .D(\i55/n181 ),
    .E(\i55/n180 ),
    .Y(\i55/n353 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i55/i148  (.A1(\i55/n72 ),
    .A2(\i55/n91 ),
    .B(\i55/n507 ),
    .C(\i55/n262 ),
    .Y(\i55/n352 ));
 NAND4xp25_ASAP7_75t_SL \i55/i149  (.A(\i55/n304 ),
    .B(\i55/n516 ),
    .C(\i55/n105 ),
    .D(\i55/n167 ),
    .Y(\i55/n351 ));
 NOR3xp33_ASAP7_75t_SL \i55/i15  (.A(\i55/n464 ),
    .B(\i55/n429 ),
    .C(\i55/n474 ),
    .Y(\i55/n486 ));
 NAND5xp2_ASAP7_75t_SL \i55/i150  (.A(\i55/n156 ),
    .B(\i55/n138 ),
    .C(\i55/n228 ),
    .D(\i55/n101 ),
    .E(\i55/n97 ),
    .Y(\i55/n350 ));
 NAND2xp5_ASAP7_75t_SL \i55/i151  (.A(\i55/n271 ),
    .B(\i55/n296 ),
    .Y(\i55/n349 ));
 NAND2xp5_ASAP7_75t_SL \i55/i152  (.A(\i55/n219 ),
    .B(\i55/n340 ),
    .Y(\i55/n348 ));
 NOR2xp33_ASAP7_75t_L \i55/i153  (.A(\i55/n318 ),
    .B(\i55/n330 ),
    .Y(\i55/n368 ));
 NAND2xp5_ASAP7_75t_SL \i55/i154  (.A(\i55/n220 ),
    .B(\i55/n342 ),
    .Y(\i55/n347 ));
 NOR2x1_ASAP7_75t_SL \i55/i155  (.A(\i55/n276 ),
    .B(\i55/n322 ),
    .Y(\i55/n366 ));
 NAND3x1_ASAP7_75t_SL \i55/i156  (.A(\i55/n254 ),
    .B(\i55/n130 ),
    .C(\i55/n140 ),
    .Y(\i55/n27 ));
 INVxp67_ASAP7_75t_SL \i55/i157  (.A(\i55/n345 ),
    .Y(\i55/n346 ));
 INVxp67_ASAP7_75t_SL \i55/i158  (.A(\i55/n7 ),
    .Y(\i55/n344 ));
 INVxp67_ASAP7_75t_SL \i55/i159  (.A(\i55/n338 ),
    .Y(\i55/n339 ));
 NAND4xp75_ASAP7_75t_SL \i55/i16  (.A(\i55/n476 ),
    .B(\i55/n445 ),
    .C(\i55/n450 ),
    .D(\i55/n440 ),
    .Y(\i55/n485 ));
 INVxp67_ASAP7_75t_SL \i55/i160  (.A(\i55/n336 ),
    .Y(\i55/n337 ));
 INVx2_ASAP7_75t_SL \i55/i161  (.A(\i55/n334 ),
    .Y(\i55/n335 ));
 INVxp67_ASAP7_75t_SL \i55/i162  (.A(\i55/n332 ),
    .Y(\i55/n333 ));
 INVxp67_ASAP7_75t_SL \i55/i163  (.A(\i55/n328 ),
    .Y(\i55/n329 ));
 INVxp67_ASAP7_75t_SL \i55/i164  (.A(\i55/n26 ),
    .Y(\i55/n326 ));
 INVx1_ASAP7_75t_SL \i55/i165  (.A(\i55/n323 ),
    .Y(\i55/n324 ));
 NAND2xp5_ASAP7_75t_SL \i55/i166  (.A(\i55/n213 ),
    .B(\i55/n211 ),
    .Y(\i55/n322 ));
 NOR2xp33_ASAP7_75t_SL \i55/i167  (.A(\i55/n248 ),
    .B(\i55/n242 ),
    .Y(\i55/n321 ));
 NAND2xp33_ASAP7_75t_SL \i55/i168  (.A(\i55/n540 ),
    .B(\i55/n199 ),
    .Y(\i55/n320 ));
 OAI21xp5_ASAP7_75t_SL \i55/i169  (.A1(\i55/n52 ),
    .A2(\i55/n564 ),
    .B(\i55/n179 ),
    .Y(\i55/n319 ));
 AND3x4_ASAP7_75t_SL \i55/i17  (.A(\i55/n467 ),
    .B(\i55/n482 ),
    .C(\i55/n472 ),
    .Y(n10[7]));
 NAND2xp5_ASAP7_75t_SL \i55/i170  (.A(\i55/n169 ),
    .B(\i55/n540 ),
    .Y(\i55/n318 ));
 AOI31xp33_ASAP7_75t_SL \i55/i171  (.A1(\i55/n52 ),
    .A2(\i55/n15 ),
    .A3(\i55/n63 ),
    .B(\i55/n45 ),
    .Y(\i55/n317 ));
 NOR3xp33_ASAP7_75t_SL \i55/i172  (.A(\i55/n201 ),
    .B(\i55/n129 ),
    .C(\i55/n115 ),
    .Y(\i55/n316 ));
 NOR3xp33_ASAP7_75t_SL \i55/i173  (.A(\i55/n108 ),
    .B(\i55/n123 ),
    .C(\i55/n248 ),
    .Y(\i55/n315 ));
 OAI31xp33_ASAP7_75t_SL \i55/i174  (.A1(\i55/n47 ),
    .A2(\i55/n49 ),
    .A3(\i55/n70 ),
    .B(\i55/n81 ),
    .Y(\i55/n314 ));
 AOI221xp5_ASAP7_75t_SL \i55/i175  (.A1(\i55/n72 ),
    .A2(\i55/n84 ),
    .B1(\i55/n55 ),
    .B2(\i55/n65 ),
    .C(\i55/n183 ),
    .Y(\i55/n313 ));
 OAI31xp33_ASAP7_75t_R \i55/i176  (.A1(\i55/n529 ),
    .A2(\i55/n71 ),
    .A3(\i55/n72 ),
    .B(\i55/n70 ),
    .Y(\i55/n312 ));
 AOI21xp5_ASAP7_75t_SL \i55/i177  (.A1(\i55/n151 ),
    .A2(\i55/n63 ),
    .B(\i55/n552 ),
    .Y(\i55/n345 ));
 AOI21xp5_ASAP7_75t_L \i55/i178  (.A1(\i55/n63 ),
    .A2(\i55/n160 ),
    .B(\i55/n80 ),
    .Y(\i55/n311 ));
 OAI221xp5_ASAP7_75t_SL \i55/i179  (.A1(\i55/n16 ),
    .A2(\i55/n83 ),
    .B1(\i55/n48 ),
    .B2(\i55/n57 ),
    .C(\i55/n559 ),
    .Y(\i55/n310 ));
 NAND4xp75_ASAP7_75t_SL \i55/i18  (.A(\i55/n475 ),
    .B(\i55/n449 ),
    .C(\i55/n458 ),
    .D(\i55/n571 ),
    .Y(\i55/n484 ));
 AOI21xp33_ASAP7_75t_SL \i55/i180  (.A1(\i55/n160 ),
    .A2(\i55/n46 ),
    .B(\i55/n497 ),
    .Y(\i55/n309 ));
 NOR3xp33_ASAP7_75t_SL \i55/i181  (.A(\i55/n222 ),
    .B(\i55/n108 ),
    .C(\i55/n134 ),
    .Y(\i55/n308 ));
 NAND3xp33_ASAP7_75t_SL \i55/i182  (.A(\i55/n19 ),
    .B(\i55/n21 ),
    .C(\i55/n158 ),
    .Y(\i55/n307 ));
 AOI22xp5_ASAP7_75t_SL \i55/i183  (.A1(\i55/n59 ),
    .A2(\i55/n147 ),
    .B1(\i55/n65 ),
    .B2(\i55/n54 ),
    .Y(\i55/n306 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i55/i184  (.A1(\i55/n80 ),
    .A2(\i55/n50 ),
    .B(\i55/n69 ),
    .C(\i55/n111 ),
    .Y(\i55/n305 ));
 OAI21xp5_ASAP7_75t_SL \i55/i185  (.A1(\i55/n61 ),
    .A2(\i55/n153 ),
    .B(\i55/n529 ),
    .Y(\i55/n304 ));
 NAND4xp25_ASAP7_75t_SL \i55/i186  (.A(\i55/n172 ),
    .B(\i55/n167 ),
    .C(\i55/n521 ),
    .D(\i55/n141 ),
    .Y(\i55/n303 ));
 NAND2xp33_ASAP7_75t_SL \i55/i187  (.A(\i55/n231 ),
    .B(\i55/n133 ),
    .Y(\i55/n302 ));
 OAI211xp5_ASAP7_75t_SL \i55/i188  (.A1(\i55/n68 ),
    .A2(\i55/n497 ),
    .B(\i55/n560 ),
    .C(\i55/n146 ),
    .Y(\i55/n343 ));
 NOR2xp67_ASAP7_75t_SL \i55/i189  (.A(\i55/n198 ),
    .B(\i55/n249 ),
    .Y(\i55/n342 ));
 NAND2x1_ASAP7_75t_SL \i55/i19  (.A(\i55/n437 ),
    .B(\i55/n468 ),
    .Y(\i55/n483 ));
 AO21x1_ASAP7_75t_SL \i55/i190  (.A1(\i55/n56 ),
    .A2(\i55/n150 ),
    .B(\i55/n135 ),
    .Y(\i55/n341 ));
 AOI21x1_ASAP7_75t_SL \i55/i191  (.A1(\i55/n54 ),
    .A2(\i55/n61 ),
    .B(\i55/n257 ),
    .Y(\i55/n340 ));
 NOR2xp33_ASAP7_75t_SL \i55/i192  (.A(\i55/n234 ),
    .B(\i55/n250 ),
    .Y(\i55/n338 ));
 OAI211xp5_ASAP7_75t_SL \i55/i193  (.A1(\i55/n63 ),
    .A2(\i55/n497 ),
    .B(\i55/n179 ),
    .C(\i55/n520 ),
    .Y(\i55/n336 ));
 OR2x2_ASAP7_75t_SL \i55/i194  (.A(\i55/n192 ),
    .B(\i55/n212 ),
    .Y(\i55/n334 ));
 AOI21xp5_ASAP7_75t_SL \i55/i195  (.A1(\i55/n71 ),
    .A2(\i55/n64 ),
    .B(\i55/n246 ),
    .Y(\i55/n332 ));
 OAI211xp5_ASAP7_75t_SL \i55/i196  (.A1(\i55/n83 ),
    .A2(\i55/n74 ),
    .B(\i55/n176 ),
    .C(\i55/n125 ),
    .Y(\i55/n331 ));
 NAND2xp5_ASAP7_75t_SL \i55/i197  (.A(\i55/n251 ),
    .B(\i55/n252 ),
    .Y(\i55/n330 ));
 NAND2xp5_ASAP7_75t_SL \i55/i198  (.A(\i55/n25 ),
    .B(\i55/n187 ),
    .Y(\i55/n328 ));
 NAND2xp5_ASAP7_75t_SL \i55/i199  (.A(\i55/n230 ),
    .B(\i55/n494 ),
    .Y(\i55/n327 ));
 INVx2_ASAP7_75t_SL \i55/i2  (.A(n11[0]),
    .Y(\i55/n2 ));
 NOR2xp67_ASAP7_75t_SL \i55/i20  (.A(\i55/n469 ),
    .B(\i55/n430 ),
    .Y(\i55/n482 ));
 OAI221xp5_ASAP7_75t_SL \i55/i200  (.A1(\i55/n57 ),
    .A2(\i55/n500 ),
    .B1(\i55/n52 ),
    .B2(\i55/n56 ),
    .C(\i55/n541 ),
    .Y(\i55/n26 ));
 NAND2xp5_ASAP7_75t_SL \i55/i201  (.A(\i55/n562 ),
    .B(\i55/n492 ),
    .Y(\i55/n325 ));
 NOR2x1_ASAP7_75t_SL \i55/i202  (.A(\i55/n232 ),
    .B(\i55/n208 ),
    .Y(\i55/n323 ));
 INVx1_ASAP7_75t_SL \i55/i203  (.A(\i55/n298 ),
    .Y(\i55/n299 ));
 INVx1_ASAP7_75t_SL \i55/i204  (.A(\i55/n294 ),
    .Y(\i55/n295 ));
 INVx1_ASAP7_75t_SL \i55/i205  (.A(\i55/n290 ),
    .Y(\i55/n291 ));
 NAND4xp25_ASAP7_75t_SL \i55/i206  (.A(\i55/n543 ),
    .B(\i55/n126 ),
    .C(\i55/n111 ),
    .D(\i55/n536 ),
    .Y(\i55/n285 ));
 AOI31xp33_ASAP7_75t_SL \i55/i207  (.A1(\i55/n525 ),
    .A2(\i55/n499 ),
    .A3(\i55/n45 ),
    .B(\i55/n46 ),
    .Y(\i55/n284 ));
 NOR4xp25_ASAP7_75t_SL \i55/i208  (.A(\i55/n103 ),
    .B(\i55/n118 ),
    .C(\i55/n178 ),
    .D(\i55/n86 ),
    .Y(\i55/n283 ));
 AOI211xp5_ASAP7_75t_SL \i55/i209  (.A1(\i55/n127 ),
    .A2(\i55/n528 ),
    .B(\i55/n165 ),
    .C(\i55/n92 ),
    .Y(\i55/n282 ));
 NAND4xp75_ASAP7_75t_SL \i55/i21  (.A(\i55/n441 ),
    .B(\i55/n453 ),
    .C(\i55/n435 ),
    .D(\i55/n438 ),
    .Y(\i55/n481 ));
 NOR2xp33_ASAP7_75t_L \i55/i210  (.A(\i55/n185 ),
    .B(\i55/n243 ),
    .Y(\i55/n281 ));
 OAI31xp33_ASAP7_75t_SL \i55/i211  (.A1(\i55/n59 ),
    .A2(\i55/n55 ),
    .A3(\i55/n81 ),
    .B(\i55/n64 ),
    .Y(\i55/n280 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i55/i212  (.A1(\i55/n497 ),
    .A2(\i55/n50 ),
    .B(\i55/n78 ),
    .C(\i55/n519 ),
    .Y(\i55/n279 ));
 OAI22xp33_ASAP7_75t_SL \i55/i213  (.A1(\i55/n74 ),
    .A2(\i55/n154 ),
    .B1(\i55/n68 ),
    .B2(\i55/n526 ),
    .Y(\i55/n278 ));
 NOR2xp33_ASAP7_75t_SL \i55/i214  (.A(\i55/n205 ),
    .B(\i55/n188 ),
    .Y(\i55/n277 ));
 OAI222xp33_ASAP7_75t_SL \i55/i215  (.A1(\i55/n80 ),
    .A2(\i55/n46 ),
    .B1(\i55/n50 ),
    .B2(\i55/n15 ),
    .C1(\i55/n499 ),
    .C2(\i55/n68 ),
    .Y(\i55/n276 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i55/i216  (.A1(\i55/n59 ),
    .A2(\i55/n58 ),
    .B(\i55/n62 ),
    .C(\i55/n161 ),
    .Y(\i55/n275 ));
 NAND2xp33_ASAP7_75t_L \i55/i217  (.A(\i55/n545 ),
    .B(\i55/n538 ),
    .Y(\i55/n274 ));
 NAND2xp33_ASAP7_75t_SL \i55/i218  (.A(\i55/n239 ),
    .B(\i55/n124 ),
    .Y(\i55/n273 ));
 AOI22xp5_ASAP7_75t_SL \i55/i219  (.A1(\i55/n71 ),
    .A2(\i55/n100 ),
    .B1(\i55/n528 ),
    .B2(\i55/n72 ),
    .Y(\i55/n272 ));
 OR3x1_ASAP7_75t_SL \i55/i22  (.A(\i55/n461 ),
    .B(\i55/n459 ),
    .C(\i55/n442 ),
    .Y(\i55/n480 ));
 OAI21xp33_ASAP7_75t_SL \i55/i220  (.A1(\i55/n109 ),
    .A2(\i55/n71 ),
    .B(\i55/n528 ),
    .Y(\i55/n271 ));
 OA21x2_ASAP7_75t_SL \i55/i221  (.A1(\i55/n46 ),
    .A2(\i55/n564 ),
    .B(\i55/n120 ),
    .Y(\i55/n270 ));
 NAND2xp5_ASAP7_75t_SL \i55/i222  (.A(\i55/n193 ),
    .B(\i55/n256 ),
    .Y(\i55/n269 ));
 NAND4xp25_ASAP7_75t_SL \i55/i223  (.A(\i55/n565 ),
    .B(\i55/n142 ),
    .C(\i55/n98 ),
    .D(\i55/n524 ),
    .Y(\i55/n268 ));
 AOI221xp5_ASAP7_75t_SL \i55/i224  (.A1(\i55/n65 ),
    .A2(\i55/n44 ),
    .B1(\i55/n51 ),
    .B2(\i55/n67 ),
    .C(\i55/n200 ),
    .Y(\i55/n267 ));
 OAI221xp5_ASAP7_75t_SL \i55/i225  (.A1(\i55/n82 ),
    .A2(\i55/n78 ),
    .B1(\i55/n515 ),
    .B2(\i55/n14 ),
    .C(\i55/n102 ),
    .Y(\i55/n301 ));
 OAI222xp33_ASAP7_75t_SL \i55/i226  (.A1(\i55/n489 ),
    .A2(\i55/n52 ),
    .B1(\i55/n57 ),
    .B2(\i55/n68 ),
    .C1(\i55/n515 ),
    .C2(\i55/n73 ),
    .Y(\i55/n266 ));
 OAI221xp5_ASAP7_75t_SL \i55/i227  (.A1(\i55/n80 ),
    .A2(\i55/n73 ),
    .B1(\i55/n515 ),
    .B2(\i55/n69 ),
    .C(\i55/n206 ),
    .Y(\i55/n265 ));
 AND3x1_ASAP7_75t_SL \i55/i228  (.A(\i55/n119 ),
    .B(\i55/n126 ),
    .C(\i55/n518 ),
    .Y(\i55/n264 ));
 AOI31xp33_ASAP7_75t_SL \i55/i229  (.A1(\i55/n52 ),
    .A2(\i55/n76 ),
    .A3(\i55/n69 ),
    .B(\i55/n56 ),
    .Y(\i55/n263 ));
 OR3x1_ASAP7_75t_SL \i55/i23  (.A(\i55/n462 ),
    .B(\i55/n428 ),
    .C(\i55/n403 ),
    .Y(\i55/n479 ));
 NAND2xp33_ASAP7_75t_SL \i55/i230  (.A(\i55/n194 ),
    .B(\i55/n227 ),
    .Y(\i55/n262 ));
 OAI221xp5_ASAP7_75t_SL \i55/i231  (.A1(\i55/n80 ),
    .A2(\i55/n76 ),
    .B1(\i55/n16 ),
    .B2(\i55/n15 ),
    .C(\i55/n238 ),
    .Y(\i55/n261 ));
 OAI222xp33_ASAP7_75t_SL \i55/i232  (.A1(\i55/n74 ),
    .A2(\i55/n76 ),
    .B1(\i55/n82 ),
    .B2(\i55/n73 ),
    .C1(\i55/n16 ),
    .C2(\i55/n63 ),
    .Y(\i55/n300 ));
 NAND3x1_ASAP7_75t_SL \i55/i233  (.A(\i55/n535 ),
    .B(\i55/n144 ),
    .C(\i55/n139 ),
    .Y(\i55/n298 ));
 AOI22xp5_ASAP7_75t_SL \i55/i234  (.A1(\i55/n143 ),
    .A2(\i55/n81 ),
    .B1(\i55/n70 ),
    .B2(\i55/n55 ),
    .Y(\i55/n297 ));
 AOI22xp5_ASAP7_75t_SL \i55/i235  (.A1(\i55/n84 ),
    .A2(\i55/n95 ),
    .B1(\i55/n47 ),
    .B2(\i55/n529 ),
    .Y(\i55/n296 ));
 AOI221x1_ASAP7_75t_SL \i55/i236  (.A1(\i55/n81 ),
    .A2(\i55/n70 ),
    .B1(\i55/n72 ),
    .B2(\i55/n507 ),
    .C(\i55/n557 ),
    .Y(\i55/n294 ));
 AOI211x1_ASAP7_75t_SL \i55/i237  (.A1(\i55/n96 ),
    .A2(\i55/n66 ),
    .B(\i55/n522 ),
    .C(\i55/n178 ),
    .Y(\i55/n293 ));
 OAI21xp5_ASAP7_75t_SL \i55/i238  (.A1(\i55/n45 ),
    .A2(\i55/n78 ),
    .B(\i55/n235 ),
    .Y(\i55/n292 ));
 NOR2x1_ASAP7_75t_SL \i55/i239  (.A(\i55/n121 ),
    .B(\i55/n191 ),
    .Y(\i55/n290 ));
 NAND3xp33_ASAP7_75t_SL \i55/i24  (.A(\i55/n473 ),
    .B(\i55/n458 ),
    .C(\i55/n441 ),
    .Y(\i55/n478 ));
 OAI221xp5_ASAP7_75t_SL \i55/i240  (.A1(\i55/n20 ),
    .A2(\i55/n82 ),
    .B1(\i55/n60 ),
    .B2(\i55/n69 ),
    .C(\i55/n563 ),
    .Y(\i55/n289 ));
 OAI211xp5_ASAP7_75t_SL \i55/i241  (.A1(\i55/n69 ),
    .A2(\i55/n551 ),
    .B(\i55/n105 ),
    .C(\i55/n490 ),
    .Y(\i55/n288 ));
 NOR2xp33_ASAP7_75t_SL \i55/i242  (.A(\i55/n131 ),
    .B(\i55/n253 ),
    .Y(\i55/n260 ));
 AOI222xp33_ASAP7_75t_SL \i55/i243  (.A1(\i55/n72 ),
    .A2(\i55/n65 ),
    .B1(\i55/n62 ),
    .B2(\i55/n44 ),
    .C1(\i55/n529 ),
    .C2(\i55/n61 ),
    .Y(\i55/n287 ));
 OAI221xp5_ASAP7_75t_SL \i55/i244  (.A1(\i55/n537 ),
    .A2(\i55/n50 ),
    .B1(\i55/n46 ),
    .B2(\i55/n56 ),
    .C(\i55/n114 ),
    .Y(\i55/n286 ));
 INVxp67_ASAP7_75t_SL \i55/i245  (.A(\i55/n494 ),
    .Y(\i55/n258 ));
 INVx1_ASAP7_75t_SL \i55/i246  (.A(\i55/n255 ),
    .Y(\i55/n256 ));
 INVx1_ASAP7_75t_SL \i55/i247  (.A(\i55/n253 ),
    .Y(\i55/n254 ));
 INVxp67_ASAP7_75t_SL \i55/i248  (.A(\i55/n246 ),
    .Y(\i55/n247 ));
 INVx1_ASAP7_75t_SL \i55/i249  (.A(\i55/n243 ),
    .Y(\i55/n244 ));
 NOR2x1_ASAP7_75t_SL \i55/i25  (.A(\i55/n384 ),
    .B(\i55/n459 ),
    .Y(\i55/n476 ));
 OAI21xp33_ASAP7_75t_SL \i55/i250  (.A1(\i55/n510 ),
    .A2(\i55/n498 ),
    .B(\i55/n523 ),
    .Y(\i55/n241 ));
 NAND2xp5_ASAP7_75t_SL \i55/i251  (.A(\i55/n495 ),
    .B(\i55/n125 ),
    .Y(\i55/n240 ));
 OAI21xp5_ASAP7_75t_SL \i55/i252  (.A1(\i55/n55 ),
    .A2(\i55/n54 ),
    .B(\i55/n505 ),
    .Y(\i55/n239 ));
 NOR2xp33_ASAP7_75t_SL \i55/i253  (.A(\i55/n132 ),
    .B(\i55/n164 ),
    .Y(\i55/n238 ));
 NAND2xp33_ASAP7_75t_L \i55/i254  (.A(\i55/n493 ),
    .B(\i55/n93 ),
    .Y(\i55/n237 ));
 NOR2xp33_ASAP7_75t_SL \i55/i255  (.A(\i55/n18 ),
    .B(\i55/n112 ),
    .Y(\i55/n236 ));
 OAI21xp33_ASAP7_75t_SL \i55/i256  (.A1(\i55/n71 ),
    .A2(\i55/n77 ),
    .B(\i55/n65 ),
    .Y(\i55/n235 ));
 OAI21xp5_ASAP7_75t_SL \i55/i257  (.A1(\i55/n537 ),
    .A2(\i55/n552 ),
    .B(\i55/n162 ),
    .Y(\i55/n234 ));
 AOI22xp5_ASAP7_75t_SL \i55/i258  (.A1(\i55/n505 ),
    .A2(\i55/n58 ),
    .B1(\i55/n507 ),
    .B2(\i55/n529 ),
    .Y(\i55/n233 ));
 OAI21xp5_ASAP7_75t_SL \i55/i259  (.A1(\i55/n15 ),
    .A2(\i55/n515 ),
    .B(\i55/n128 ),
    .Y(\i55/n232 ));
 NOR2x1_ASAP7_75t_SL \i55/i26  (.A(\i55/n443 ),
    .B(\i55/n439 ),
    .Y(\i55/n475 ));
 OAI21xp5_ASAP7_75t_SL \i55/i260  (.A1(\i55/n71 ),
    .A2(\i55/n54 ),
    .B(\i55/n67 ),
    .Y(\i55/n231 ));
 AOI22xp5_ASAP7_75t_SL \i55/i261  (.A1(\i55/n44 ),
    .A2(\i55/n84 ),
    .B1(\i55/n47 ),
    .B2(\i55/n71 ),
    .Y(\i55/n230 ));
 OA21x2_ASAP7_75t_SL \i55/i262  (.A1(\i55/n500 ),
    .A2(\i55/n13 ),
    .B(\i55/n166 ),
    .Y(\i55/n259 ));
 AOI21xp33_ASAP7_75t_SL \i55/i263  (.A1(\i55/n68 ),
    .A2(\i55/n500 ),
    .B(\i55/n45 ),
    .Y(\i55/n229 ));
 OAI21xp5_ASAP7_75t_SL \i55/i264  (.A1(\i55/n507 ),
    .A2(\i55/n84 ),
    .B(\i55/n79 ),
    .Y(\i55/n228 ));
 OAI21xp5_ASAP7_75t_SL \i55/i265  (.A1(\i55/n67 ),
    .A2(\i55/n47 ),
    .B(\i55/n79 ),
    .Y(\i55/n227 ));
 AOI21xp33_ASAP7_75t_SL \i55/i266  (.A1(\i55/n63 ),
    .A2(\i55/n78 ),
    .B(\i55/n45 ),
    .Y(\i55/n226 ));
 OAI21xp5_ASAP7_75t_SL \i55/i267  (.A1(\i55/n537 ),
    .A2(\i55/n515 ),
    .B(\i55/n23 ),
    .Y(\i55/n225 ));
 AOI22xp5_ASAP7_75t_SL \i55/i268  (.A1(\i55/n61 ),
    .A2(\i55/n59 ),
    .B1(\i55/n507 ),
    .B2(\i55/n58 ),
    .Y(\i55/n224 ));
 AOI21xp33_ASAP7_75t_SL \i55/i269  (.A1(\i55/n497 ),
    .A2(\i55/n45 ),
    .B(\i55/n69 ),
    .Y(\i55/n223 ));
 NAND3xp33_ASAP7_75t_SL \i55/i27  (.A(\i55/n423 ),
    .B(\i55/n580 ),
    .C(\i55/n547 ),
    .Y(\i55/n474 ));
 NAND2xp5_ASAP7_75t_SL \i55/i270  (.A(\i55/n79 ),
    .B(\i55/n152 ),
    .Y(\i55/n25 ));
 NAND2xp5_ASAP7_75t_L \i55/i271  (.A(\i55/n179 ),
    .B(\i55/n520 ),
    .Y(\i55/n222 ));
 OAI22xp5_ASAP7_75t_SL \i55/i272  (.A1(\i55/n498 ),
    .A2(\i55/n80 ),
    .B1(\i55/n85 ),
    .B2(\i55/n13 ),
    .Y(\i55/n257 ));
 OAI22xp5_ASAP7_75t_SL \i55/i273  (.A1(\i55/n85 ),
    .A2(\i55/n515 ),
    .B1(\i55/n16 ),
    .B2(\i55/n68 ),
    .Y(\i55/n255 ));
 OAI22xp5_ASAP7_75t_SL \i55/i274  (.A1(\i55/n83 ),
    .A2(\i55/n57 ),
    .B1(\i55/n537 ),
    .B2(\i55/n74 ),
    .Y(\i55/n253 ));
 AOI22xp5_ASAP7_75t_SL \i55/i275  (.A1(\i55/n66 ),
    .A2(\i55/n81 ),
    .B1(\i55/n62 ),
    .B2(\i55/n77 ),
    .Y(\i55/n252 ));
 AOI22xp5_ASAP7_75t_SL \i55/i276  (.A1(\i55/n66 ),
    .A2(\i55/n59 ),
    .B1(\i55/n527 ),
    .B2(\i55/n58 ),
    .Y(\i55/n251 ));
 OAI22xp5_ASAP7_75t_SL \i55/i277  (.A1(\i55/n69 ),
    .A2(\i55/n74 ),
    .B1(\i55/n515 ),
    .B2(\i55/n48 ),
    .Y(\i55/n250 ));
 OAI22xp33_ASAP7_75t_SL \i55/i278  (.A1(\i55/n85 ),
    .A2(\i55/n82 ),
    .B1(\i55/n46 ),
    .B2(\i55/n489 ),
    .Y(\i55/n249 ));
 NAND2xp5_ASAP7_75t_L \i55/i279  (.A(\i55/n17 ),
    .B(\i55/n148 ),
    .Y(\i55/n248 ));
 NOR2x1_ASAP7_75t_SL \i55/i28  (.A(\i55/n448 ),
    .B(\i55/n412 ),
    .Y(\i55/n473 ));
 OAI22xp5_ASAP7_75t_SL \i55/i280  (.A1(\i55/n537 ),
    .A2(\i55/n82 ),
    .B1(\i55/n68 ),
    .B2(\i55/n552 ),
    .Y(\i55/n246 ));
 OAI21xp5_ASAP7_75t_SL \i55/i281  (.A1(\i55/n71 ),
    .A2(\i55/n51 ),
    .B(\i55/n505 ),
    .Y(\i55/n245 ));
 NOR2xp33_ASAP7_75t_L \i55/i282  (.A(\i55/n13 ),
    .B(\i55/n20 ),
    .Y(\i55/n243 ));
 NAND2xp33_ASAP7_75t_L \i55/i283  (.A(\i55/n105 ),
    .B(\i55/n490 ),
    .Y(\i55/n221 ));
 OAI21xp5_ASAP7_75t_SL \i55/i284  (.A1(\i55/n69 ),
    .A2(\i55/n57 ),
    .B(\i55/n104 ),
    .Y(\i55/n242 ));
 INVxp67_ASAP7_75t_SL \i55/i285  (.A(\i55/n217 ),
    .Y(\i55/n218 ));
 INVxp67_ASAP7_75t_SL \i55/i286  (.A(\i55/n215 ),
    .Y(\i55/n216 ));
 INVx1_ASAP7_75t_SL \i55/i287  (.A(\i55/n213 ),
    .Y(\i55/n214 ));
 INVx1_ASAP7_75t_SL \i55/i288  (.A(\i55/n210 ),
    .Y(\i55/n211 ));
 INVxp67_ASAP7_75t_SL \i55/i289  (.A(\i55/n559 ),
    .Y(\i55/n209 ));
 NOR5xp2_ASAP7_75t_SL \i55/i29  (.A(\i55/n414 ),
    .B(\i55/n361 ),
    .C(\i55/n405 ),
    .D(\i55/n327 ),
    .E(\i55/n331 ),
    .Y(\i55/n472 ));
 INVxp67_ASAP7_75t_SL \i55/i290  (.A(\i55/n205 ),
    .Y(\i55/n206 ));
 INVxp67_ASAP7_75t_SL \i55/i291  (.A(\i55/n203 ),
    .Y(\i55/n204 ));
 OAI22xp33_ASAP7_75t_SL \i55/i292  (.A1(\i55/n48 ),
    .A2(\i55/n82 ),
    .B1(\i55/n56 ),
    .B2(\i55/n498 ),
    .Y(\i55/n198 ));
 OAI21xp33_ASAP7_75t_SL \i55/i293  (.A1(\i55/n58 ),
    .A2(\i55/n75 ),
    .B(\i55/n507 ),
    .Y(\i55/n197 ));
 OAI21xp5_ASAP7_75t_SL \i55/i294  (.A1(\i55/n14 ),
    .A2(\i55/n489 ),
    .B(\i55/n116 ),
    .Y(\i55/n196 ));
 AOI21xp33_ASAP7_75t_SL \i55/i295  (.A1(\i55/n515 ),
    .A2(\i55/n74 ),
    .B(\i55/n76 ),
    .Y(\i55/n195 ));
 OAI21xp5_ASAP7_75t_SL \i55/i296  (.A1(\i55/n44 ),
    .A2(\i55/n51 ),
    .B(\i55/n49 ),
    .Y(\i55/n194 ));
 AOI22xp33_ASAP7_75t_SL \i55/i297  (.A1(\i55/n66 ),
    .A2(\i55/n71 ),
    .B1(\i55/n62 ),
    .B2(\i55/n55 ),
    .Y(\i55/n193 ));
 OAI22xp33_ASAP7_75t_SL \i55/i298  (.A1(\i55/n498 ),
    .A2(\i55/n45 ),
    .B1(\i55/n80 ),
    .B2(\i55/n63 ),
    .Y(\i55/n192 ));
 AOI22xp5_ASAP7_75t_SL \i55/i299  (.A1(\i55/n527 ),
    .A2(\i55/n79 ),
    .B1(\i55/n505 ),
    .B2(\i55/n54 ),
    .Y(\i55/n220 ));
 INVx2_ASAP7_75t_SL \i55/i3  (.A(\i55/n32 ),
    .Y(\i55/n3 ));
 NOR3xp33_ASAP7_75t_SL \i55/i30  (.A(\i55/n410 ),
    .B(\i55/n425 ),
    .C(\i55/n457 ),
    .Y(\i55/n471 ));
 OAI22xp33_ASAP7_75t_SL \i55/i300  (.A1(\i55/n16 ),
    .A2(\i55/n498 ),
    .B1(\i55/n74 ),
    .B2(\i55/n78 ),
    .Y(\i55/n191 ));
 OAI22xp5_ASAP7_75t_SL \i55/i301  (.A1(\i55/n83 ),
    .A2(\i55/n489 ),
    .B1(\i55/n14 ),
    .B2(\i55/n80 ),
    .Y(\i55/n190 ));
 OAI22xp5_ASAP7_75t_SL \i55/i302  (.A1(\i55/n63 ),
    .A2(\i55/n489 ),
    .B1(\i55/n78 ),
    .B2(\i55/n497 ),
    .Y(\i55/n189 ));
 AOI22xp33_ASAP7_75t_SL \i55/i303  (.A1(\i55/n44 ),
    .A2(\i55/n47 ),
    .B1(\i55/n527 ),
    .B2(\i55/n71 ),
    .Y(\i55/n219 ));
 OAI22xp33_ASAP7_75t_SL \i55/i304  (.A1(\i55/n50 ),
    .A2(\i55/n498 ),
    .B1(\i55/n13 ),
    .B2(\i55/n52 ),
    .Y(\i55/n188 ));
 AOI22xp5_ASAP7_75t_SL \i55/i305  (.A1(\i55/n65 ),
    .A2(\i55/n75 ),
    .B1(\i55/n47 ),
    .B2(\i55/n77 ),
    .Y(\i55/n187 ));
 OAI22xp5_ASAP7_75t_SL \i55/i306  (.A1(\i55/n498 ),
    .A2(\i55/n82 ),
    .B1(\i55/n68 ),
    .B2(\i55/n13 ),
    .Y(\i55/n186 ));
 OAI21xp5_ASAP7_75t_SL \i55/i307  (.A1(\i55/n73 ),
    .A2(\i55/n56 ),
    .B(\i55/n124 ),
    .Y(\i55/n185 ));
 OAI21xp5_ASAP7_75t_SL \i55/i308  (.A1(\i55/n46 ),
    .A2(\i55/n57 ),
    .B(\i55/n113 ),
    .Y(\i55/n217 ));
 AOI22xp5_ASAP7_75t_SL \i55/i309  (.A1(\i55/n44 ),
    .A2(\i55/n67 ),
    .B1(\i55/n47 ),
    .B2(\i55/n54 ),
    .Y(\i55/n215 ));
 NOR2x1_ASAP7_75t_SL \i55/i31  (.A(\i55/n454 ),
    .B(\i55/n415 ),
    .Y(\i55/n470 ));
 AOI22xp5_ASAP7_75t_SL \i55/i310  (.A1(\i55/n49 ),
    .A2(\i55/n51 ),
    .B1(\i55/n59 ),
    .B2(\i55/n65 ),
    .Y(\i55/n213 ));
 OA21x2_ASAP7_75t_SL \i55/i311  (.A1(\i55/n52 ),
    .A2(\i55/n56 ),
    .B(\i55/n541 ),
    .Y(\i55/n184 ));
 OAI22xp5_ASAP7_75t_SL \i55/i312  (.A1(\i55/n52 ),
    .A2(\i55/n74 ),
    .B1(\i55/n68 ),
    .B2(\i55/n56 ),
    .Y(\i55/n212 ));
 OAI22xp5_ASAP7_75t_SL \i55/i313  (.A1(\i55/n45 ),
    .A2(\i55/n14 ),
    .B1(\i55/n498 ),
    .B2(\i55/n499 ),
    .Y(\i55/n183 ));
 NAND2xp33_ASAP7_75t_SL \i55/i314  (.A(\i55/n180 ),
    .B(\i55/n181 ),
    .Y(\i55/n182 ));
 OAI22x1_ASAP7_75t_SL \i55/i315  (.A1(\i55/n15 ),
    .A2(\i55/n82 ),
    .B1(\i55/n48 ),
    .B2(\i55/n510 ),
    .Y(\i55/n210 ));
 AO22x2_ASAP7_75t_SL \i55/i316  (.A1(\i55/n84 ),
    .A2(\i55/n81 ),
    .B1(\i55/n53 ),
    .B2(\i55/n77 ),
    .Y(\i55/n208 ));
 OAI21xp5_ASAP7_75t_SL \i55/i317  (.A1(\i55/n73 ),
    .A2(\i55/n50 ),
    .B(\i55/n542 ),
    .Y(\i55/n207 ));
 OAI22xp5_ASAP7_75t_L \i55/i318  (.A1(\i55/n76 ),
    .A2(\i55/n45 ),
    .B1(\i55/n46 ),
    .B2(\i55/n74 ),
    .Y(\i55/n205 ));
 OAI22xp5_ASAP7_75t_SL \i55/i319  (.A1(\i55/n63 ),
    .A2(\i55/n50 ),
    .B1(\i55/n68 ),
    .B2(\i55/n74 ),
    .Y(\i55/n203 ));
 NAND2xp5_ASAP7_75t_SL \i55/i32  (.A(\i55/n413 ),
    .B(\i55/n431 ),
    .Y(\i55/n469 ));
 AOI22xp5_ASAP7_75t_SL \i55/i320  (.A1(\i55/n44 ),
    .A2(\i55/n49 ),
    .B1(\i55/n70 ),
    .B2(\i55/n77 ),
    .Y(\i55/n202 ));
 OAI22xp5_ASAP7_75t_R \i55/i321  (.A1(\i55/n52 ),
    .A2(\i55/n60 ),
    .B1(\i55/n68 ),
    .B2(\i55/n510 ),
    .Y(\i55/n201 ));
 OAI22xp5_ASAP7_75t_SL \i55/i322  (.A1(\i55/n500 ),
    .A2(\i55/n74 ),
    .B1(\i55/n69 ),
    .B2(\i55/n80 ),
    .Y(\i55/n24 ));
 OAI22xp5_ASAP7_75t_SL \i55/i323  (.A1(\i55/n52 ),
    .A2(\i55/n50 ),
    .B1(\i55/n56 ),
    .B2(\i55/n48 ),
    .Y(\i55/n200 ));
 AOI22xp5_ASAP7_75t_SL \i55/i324  (.A1(\i55/n527 ),
    .A2(\i55/n51 ),
    .B1(\i55/n64 ),
    .B2(\i55/n529 ),
    .Y(\i55/n199 ));
 INVxp67_ASAP7_75t_SL \i55/i325  (.A(\i55/n522 ),
    .Y(\i55/n177 ));
 INVx1_ASAP7_75t_SL \i55/i326  (.A(\i55/n175 ),
    .Y(\i55/n176 ));
 INVxp67_ASAP7_75t_SL \i55/i327  (.A(\i55/n562 ),
    .Y(\i55/n174 ));
 INVxp67_ASAP7_75t_SL \i55/i328  (.A(\i55/n172 ),
    .Y(\i55/n173 ));
 INVxp67_ASAP7_75t_SL \i55/i329  (.A(\i55/n523 ),
    .Y(\i55/n171 ));
 NOR3x1_ASAP7_75t_SL \i55/i33  (.A(\i55/n27 ),
    .B(\i55/n427 ),
    .C(\i55/n569 ),
    .Y(\i55/n477 ));
 INVxp67_ASAP7_75t_SL \i55/i330  (.A(\i55/n168 ),
    .Y(\i55/n169 ));
 INVxp67_ASAP7_75t_SL \i55/i331  (.A(\i55/n162 ),
    .Y(\i55/n163 ));
 INVxp67_ASAP7_75t_SL \i55/i332  (.A(\i55/n493 ),
    .Y(\i55/n161 ));
 INVxp67_ASAP7_75t_SL \i55/i333  (.A(\i55/n158 ),
    .Y(\i55/n159 ));
 INVxp67_ASAP7_75t_SL \i55/i334  (.A(\i55/n563 ),
    .Y(\i55/n157 ));
 INVxp67_ASAP7_75t_SL \i55/i335  (.A(\i55/n154 ),
    .Y(\i55/n155 ));
 INVxp67_ASAP7_75t_SL \i55/i336  (.A(\i55/n20 ),
    .Y(\i55/n153 ));
 INVx1_ASAP7_75t_SL \i55/i337  (.A(\i55/n152 ),
    .Y(\i55/n151 ));
 NAND2xp5_ASAP7_75t_SL \i55/i338  (.A(\i55/n67 ),
    .B(\i55/n79 ),
    .Y(\i55/n181 ));
 NAND2xp5_ASAP7_75t_SL \i55/i339  (.A(\i55/n505 ),
    .B(\i55/n77 ),
    .Y(\i55/n150 ));
 NOR3xp33_ASAP7_75t_SL \i55/i34  (.A(\i55/n371 ),
    .B(\i55/n27 ),
    .C(\i55/n451 ),
    .Y(\i55/n467 ));
 NAND2xp5_ASAP7_75t_SL \i55/i340  (.A(\i55/n78 ),
    .B(\i55/n76 ),
    .Y(\i55/n149 ));
 NAND2xp5_ASAP7_75t_SL \i55/i341  (.A(\i55/n47 ),
    .B(\i55/n81 ),
    .Y(\i55/n148 ));
 NAND2xp33_ASAP7_75t_SL \i55/i342  (.A(\i55/n63 ),
    .B(\i55/n537 ),
    .Y(\i55/n147 ));
 NAND2xp5_ASAP7_75t_SL \i55/i343  (.A(\i55/n58 ),
    .B(\i55/n61 ),
    .Y(\i55/n146 ));
 NAND2xp5_ASAP7_75t_SL \i55/i344  (.A(\i55/n58 ),
    .B(\i55/n65 ),
    .Y(\i55/n180 ));
 NAND2xp5_ASAP7_75t_SL \i55/i345  (.A(\i55/n65 ),
    .B(\i55/n79 ),
    .Y(\i55/n145 ));
 NAND2xp5_ASAP7_75t_SL \i55/i346  (.A(\i55/n4 ),
    .B(\i55/n61 ),
    .Y(\i55/n144 ));
 NAND2xp5_ASAP7_75t_SL \i55/i347  (.A(\i55/n68 ),
    .B(\i55/n14 ),
    .Y(\i55/n143 ));
 NAND2xp5_ASAP7_75t_SL \i55/i348  (.A(\i55/n67 ),
    .B(\i55/n4 ),
    .Y(\i55/n142 ));
 NAND2xp5_ASAP7_75t_SL \i55/i349  (.A(\i55/n529 ),
    .B(\i55/n70 ),
    .Y(\i55/n141 ));
 NOR2xp67_ASAP7_75t_SL \i55/i35  (.A(\i55/n432 ),
    .B(\i55/n27 ),
    .Y(\i55/n466 ));
 NAND2xp5_ASAP7_75t_SL \i55/i350  (.A(\i55/n65 ),
    .B(\i55/n529 ),
    .Y(\i55/n140 ));
 NAND2xp5_ASAP7_75t_SL \i55/i351  (.A(\i55/n44 ),
    .B(\i55/n53 ),
    .Y(\i55/n139 ));
 NAND2xp5_ASAP7_75t_SL \i55/i352  (.A(\i55/n44 ),
    .B(\i55/n507 ),
    .Y(\i55/n179 ));
 AND2x2_ASAP7_75t_SL \i55/i353  (.A(\i55/n53 ),
    .B(\i55/n71 ),
    .Y(\i55/n178 ));
 AND2x2_ASAP7_75t_SL \i55/i354  (.A(\i55/n527 ),
    .B(\i55/n529 ),
    .Y(\i55/n175 ));
 NAND2xp5_ASAP7_75t_SL \i55/i355  (.A(\i55/n529 ),
    .B(\i55/n62 ),
    .Y(\i55/n23 ));
 NAND2xp5_ASAP7_75t_SL \i55/i356  (.A(\i55/n84 ),
    .B(\i55/n51 ),
    .Y(\i55/n172 ));
 AND2x2_ASAP7_75t_SL \i55/i357  (.A(\i55/n67 ),
    .B(\i55/n59 ),
    .Y(\i55/n170 ));
 NOR2xp33_ASAP7_75t_SL \i55/i358  (.A(\i55/n500 ),
    .B(\i55/n515 ),
    .Y(\i55/n22 ));
 NOR2xp33_ASAP7_75t_SL \i55/i359  (.A(\i55/n56 ),
    .B(\i55/n500 ),
    .Y(\i55/n168 ));
 NOR3xp33_ASAP7_75t_SL \i55/i36  (.A(\i55/n411 ),
    .B(\i55/n8 ),
    .C(\i55/n406 ),
    .Y(\i55/n465 ));
 NAND2xp5_ASAP7_75t_SL \i55/i360  (.A(\i55/n66 ),
    .B(\i55/n4 ),
    .Y(\i55/n138 ));
 NAND2xp5_ASAP7_75t_SL \i55/i361  (.A(\i55/n72 ),
    .B(\i55/n66 ),
    .Y(\i55/n167 ));
 NAND2xp5_ASAP7_75t_SL \i55/i362  (.A(\i55/n64 ),
    .B(\i55/n58 ),
    .Y(\i55/n166 ));
 NAND2xp5_ASAP7_75t_SL \i55/i363  (.A(\i55/n59 ),
    .B(\i55/n61 ),
    .Y(\i55/n137 ));
 NOR2xp33_ASAP7_75t_SL \i55/i364  (.A(\i55/n498 ),
    .B(\i55/n74 ),
    .Y(\i55/n165 ));
 AND2x2_ASAP7_75t_SL \i55/i365  (.A(\i55/n65 ),
    .B(\i55/n4 ),
    .Y(\i55/n164 ));
 NOR2xp33_ASAP7_75t_SL \i55/i366  (.A(\i55/n15 ),
    .B(\i55/n13 ),
    .Y(\i55/n136 ));
 NAND2xp5_ASAP7_75t_SL \i55/i367  (.A(\i55/n66 ),
    .B(\i55/n51 ),
    .Y(\i55/n162 ));
 NOR2xp33_ASAP7_75t_SL \i55/i368  (.A(\i55/n64 ),
    .B(\i55/n505 ),
    .Y(\i55/n135 ));
 NOR2xp33_ASAP7_75t_SL \i55/i369  (.A(\i55/n498 ),
    .B(\i55/n552 ),
    .Y(\i55/n134 ));
 NAND4xp25_ASAP7_75t_SL \i55/i37  (.A(\i55/n394 ),
    .B(\i55/n388 ),
    .C(\i55/n387 ),
    .D(\i55/n419 ),
    .Y(\i55/n464 ));
 NOR2xp33_ASAP7_75t_L \i55/i370  (.A(\i55/n84 ),
    .B(\i55/n49 ),
    .Y(\i55/n160 ));
 NAND2xp5_ASAP7_75t_SL \i55/i371  (.A(\i55/n64 ),
    .B(\i55/n75 ),
    .Y(\i55/n21 ));
 NAND2xp5_ASAP7_75t_SL \i55/i372  (.A(\i55/n84 ),
    .B(\i55/n54 ),
    .Y(\i55/n158 ));
 NAND2xp5_ASAP7_75t_SL \i55/i373  (.A(\i55/n84 ),
    .B(\i55/n529 ),
    .Y(\i55/n156 ));
 NAND2xp5_ASAP7_75t_SL \i55/i374  (.A(\i55/n67 ),
    .B(\i55/n72 ),
    .Y(\i55/n133 ));
 NOR2xp67_ASAP7_75t_SL \i55/i375  (.A(\i55/n505 ),
    .B(\i55/n67 ),
    .Y(\i55/n154 ));
 NOR2xp33_ASAP7_75t_SL \i55/i376  (.A(\i55/n57 ),
    .B(\i55/n78 ),
    .Y(\i55/n132 ));
 NOR2x1_ASAP7_75t_SL \i55/i377  (.A(\i55/n64 ),
    .B(\i55/n528 ),
    .Y(\i55/n20 ));
 OR2x2_ASAP7_75t_SL \i55/i378  (.A(\i55/n49 ),
    .B(\i55/n66 ),
    .Y(\i55/n152 ));
 INVxp67_ASAP7_75t_SL \i55/i379  (.A(\i55/n130 ),
    .Y(\i55/n131 ));
 NAND3xp33_ASAP7_75t_L \i55/i38  (.A(\i55/n368 ),
    .B(\i55/n388 ),
    .C(\i55/n436 ),
    .Y(\i55/n463 ));
 INVxp67_ASAP7_75t_SL \i55/i380  (.A(\i55/n128 ),
    .Y(\i55/n129 ));
 INVx1_ASAP7_75t_SL \i55/i381  (.A(\i55/n525 ),
    .Y(\i55/n127 ));
 INVxp67_ASAP7_75t_SL \i55/i382  (.A(\i55/n565 ),
    .Y(\i55/n122 ));
 INVxp67_ASAP7_75t_SL \i55/i383  (.A(\i55/n120 ),
    .Y(\i55/n121 ));
 INVxp67_ASAP7_75t_SL \i55/i384  (.A(\i55/n118 ),
    .Y(\i55/n119 ));
 INVxp67_ASAP7_75t_SL \i55/i385  (.A(\i55/n116 ),
    .Y(\i55/n117 ));
 INVxp67_ASAP7_75t_SL \i55/i386  (.A(\i55/n114 ),
    .Y(\i55/n115 ));
 INVxp67_ASAP7_75t_SL \i55/i387  (.A(\i55/n112 ),
    .Y(\i55/n113 ));
 INVxp67_ASAP7_75t_SL \i55/i388  (.A(\i55/n543 ),
    .Y(\i55/n106 ));
 INVx1_ASAP7_75t_SL \i55/i389  (.A(\i55/n545 ),
    .Y(\i55/n103 ));
 NAND3xp33_ASAP7_75t_SL \i55/i39  (.A(\i55/n373 ),
    .B(\i55/n421 ),
    .C(\i55/n407 ),
    .Y(\i55/n462 ));
 INVx1_ASAP7_75t_SL \i55/i390  (.A(\i55/n17 ),
    .Y(\i55/n18 ));
 NAND2xp5_ASAP7_75t_SL \i55/i391  (.A(\i55/n528 ),
    .B(\i55/n71 ),
    .Y(\i55/n102 ));
 NAND2xp5_ASAP7_75t_SL \i55/i392  (.A(\i55/n49 ),
    .B(\i55/n72 ),
    .Y(\i55/n101 ));
 NAND2xp5_ASAP7_75t_SL \i55/i393  (.A(\i55/n73 ),
    .B(\i55/n69 ),
    .Y(\i55/n100 ));
 NAND2xp33_ASAP7_75t_SL \i55/i394  (.A(\i55/n72 ),
    .B(\i55/n47 ),
    .Y(\i55/n99 ));
 NAND2xp5_ASAP7_75t_SL \i55/i395  (.A(\i55/n507 ),
    .B(\i55/n59 ),
    .Y(\i55/n98 ));
 NAND2xp5_ASAP7_75t_SL \i55/i396  (.A(\i55/n70 ),
    .B(\i55/n54 ),
    .Y(\i55/n97 ));
 NAND2xp5_ASAP7_75t_L \i55/i397  (.A(\i55/n16 ),
    .B(\i55/n45 ),
    .Y(\i55/n96 ));
 NAND2xp33_ASAP7_75t_SL \i55/i398  (.A(\i55/n60 ),
    .B(\i55/n489 ),
    .Y(\i55/n95 ));
 NAND2xp5_ASAP7_75t_SL \i55/i399  (.A(\i55/n62 ),
    .B(\i55/n58 ),
    .Y(\i55/n94 ));
 INVx2_ASAP7_75t_SL \i55/i4  (.A(\i55/n489 ),
    .Y(\i55/n4 ));
 NAND2xp5_ASAP7_75t_L \i55/i40  (.A(\i55/n420 ),
    .B(\i55/n452 ),
    .Y(\i55/n461 ));
 NAND2xp5_ASAP7_75t_SL \i55/i400  (.A(\i55/n527 ),
    .B(\i55/n55 ),
    .Y(\i55/n130 ));
 NAND2xp5_ASAP7_75t_SL \i55/i401  (.A(\i55/n528 ),
    .B(\i55/n58 ),
    .Y(\i55/n93 ));
 NOR2xp33_ASAP7_75t_SL \i55/i402  (.A(\i55/n57 ),
    .B(\i55/n537 ),
    .Y(\i55/n92 ));
 NAND2xp5_ASAP7_75t_SL \i55/i403  (.A(\i55/n505 ),
    .B(\i55/n59 ),
    .Y(\i55/n128 ));
 NAND2xp5_ASAP7_75t_SL \i55/i404  (.A(\i55/n62 ),
    .B(\i55/n75 ),
    .Y(\i55/n126 ));
 NAND2xp5_ASAP7_75t_SL \i55/i405  (.A(\i55/n507 ),
    .B(\i55/n54 ),
    .Y(\i55/n125 ));
 NAND2xp5_ASAP7_75t_SL \i55/i406  (.A(\i55/n53 ),
    .B(\i55/n58 ),
    .Y(\i55/n124 ));
 AND2x2_ASAP7_75t_SL \i55/i407  (.A(\i55/n62 ),
    .B(\i55/n51 ),
    .Y(\i55/n123 ));
 NAND2xp5_ASAP7_75t_SL \i55/i408  (.A(\i55/n528 ),
    .B(\i55/n51 ),
    .Y(\i55/n120 ));
 NOR2xp67_ASAP7_75t_SL \i55/i409  (.A(\i55/n52 ),
    .B(\i55/n80 ),
    .Y(\i55/n118 ));
 NAND2xp33_ASAP7_75t_SL \i55/i41  (.A(\i55/n417 ),
    .B(\i55/n434 ),
    .Y(\i55/n460 ));
 NAND2xp5_ASAP7_75t_SL \i55/i410  (.A(\i55/n47 ),
    .B(\i55/n51 ),
    .Y(\i55/n116 ));
 NAND2xp33_ASAP7_75t_L \i55/i411  (.A(\i55/n50 ),
    .B(\i55/n510 ),
    .Y(\i55/n91 ));
 NAND2x1_ASAP7_75t_SL \i55/i412  (.A(\i55/n44 ),
    .B(\i55/n527 ),
    .Y(\i55/n114 ));
 NOR2xp33_ASAP7_75t_SL \i55/i413  (.A(\i55/n45 ),
    .B(\i55/n537 ),
    .Y(\i55/n112 ));
 NAND2xp5_ASAP7_75t_SL \i55/i414  (.A(\i55/n49 ),
    .B(\i55/n75 ),
    .Y(\i55/n19 ));
 NAND2xp5_ASAP7_75t_SL \i55/i415  (.A(\i55/n49 ),
    .B(\i55/n77 ),
    .Y(\i55/n111 ));
 AND2x2_ASAP7_75t_SL \i55/i416  (.A(\i55/n527 ),
    .B(\i55/n77 ),
    .Y(\i55/n110 ));
 NAND2xp5_ASAP7_75t_L \i55/i417  (.A(\i55/n13 ),
    .B(\i55/n16 ),
    .Y(\i55/n109 ));
 AND2x2_ASAP7_75t_SL \i55/i418  (.A(\i55/n527 ),
    .B(\i55/n59 ),
    .Y(\i55/n108 ));
 NOR2xp33_ASAP7_75t_SL \i55/i419  (.A(\i55/n60 ),
    .B(\i55/n46 ),
    .Y(\i55/n90 ));
 NOR2x1_ASAP7_75t_SL \i55/i42  (.A(\i55/n433 ),
    .B(\i55/n442 ),
    .Y(\i55/n468 ));
 NOR2xp33_ASAP7_75t_SL \i55/i420  (.A(\i55/n56 ),
    .B(\i55/n48 ),
    .Y(\i55/n89 ));
 NOR2xp67_ASAP7_75t_SL \i55/i421  (.A(\i55/n55 ),
    .B(\i55/n71 ),
    .Y(\i55/n107 ));
 NAND2xp5_ASAP7_75t_SL \i55/i422  (.A(\i55/n62 ),
    .B(\i55/n77 ),
    .Y(\i55/n88 ));
 NAND2xp5_ASAP7_75t_SL \i55/i423  (.A(\i55/n507 ),
    .B(\i55/n77 ),
    .Y(\i55/n105 ));
 NAND2xp5_ASAP7_75t_SL \i55/i424  (.A(\i55/n527 ),
    .B(\i55/n72 ),
    .Y(\i55/n104 ));
 NOR2xp33_ASAP7_75t_SL \i55/i425  (.A(\i55/n85 ),
    .B(\i55/n13 ),
    .Y(\i55/n87 ));
 NOR2xp33_ASAP7_75t_SL \i55/i426  (.A(\i55/n85 ),
    .B(\i55/n57 ),
    .Y(\i55/n86 ));
 NAND2xp5_ASAP7_75t_SL \i55/i427  (.A(\i55/n62 ),
    .B(\i55/n54 ),
    .Y(\i55/n17 ));
 INVx2_ASAP7_75t_SL \i55/i428  (.A(\i55/n527 ),
    .Y(\i55/n85 ));
 INVx1_ASAP7_75t_SL \i55/i429  (.A(\i55/n84 ),
    .Y(\i55/n83 ));
 NAND2xp33_ASAP7_75t_L \i55/i43  (.A(\i55/n422 ),
    .B(\i55/n396 ),
    .Y(\i55/n457 ));
 INVx3_ASAP7_75t_SL \i55/i430  (.A(\i55/n82 ),
    .Y(\i55/n81 ));
 INVx5_ASAP7_75t_SL \i55/i431  (.A(\i55/n80 ),
    .Y(\i55/n79 ));
 INVx2_ASAP7_75t_SL \i55/i432  (.A(\i55/n505 ),
    .Y(\i55/n78 ));
 INVx2_ASAP7_75t_SL \i55/i433  (.A(\i55/n528 ),
    .Y(\i55/n76 ));
 INVx4_ASAP7_75t_SL \i55/i434  (.A(\i55/n75 ),
    .Y(\i55/n74 ));
 INVx2_ASAP7_75t_SL \i55/i435  (.A(\i55/n507 ),
    .Y(\i55/n73 ));
 INVx3_ASAP7_75t_SL \i55/i436  (.A(\i55/n70 ),
    .Y(\i55/n69 ));
 INVx3_ASAP7_75t_SL \i55/i437  (.A(\i55/n68 ),
    .Y(\i55/n67 ));
 AND2x4_ASAP7_75t_SL \i55/i438  (.A(\i55/n40 ),
    .B(\i55/n38 ),
    .Y(\i55/n84 ));
 OR2x2_ASAP7_75t_SL \i55/i439  (.A(\i55/n31 ),
    .B(\i55/n6 ),
    .Y(\i55/n82 ));
 NAND2xp33_ASAP7_75t_L \i55/i44  (.A(\i55/n420 ),
    .B(\i55/n401 ),
    .Y(\i55/n456 ));
 OR2x6_ASAP7_75t_SL \i55/i440  (.A(\i55/n34 ),
    .B(\i55/n43 ),
    .Y(\i55/n80 ));
 AND2x4_ASAP7_75t_SL \i55/i441  (.A(\i55/n512 ),
    .B(\i55/n36 ),
    .Y(\i55/n77 ));
 NAND2x1_ASAP7_75t_SL \i55/i442  (.A(\i55/n512 ),
    .B(\i55/n36 ),
    .Y(\i55/n16 ));
 AND2x4_ASAP7_75t_SL \i55/i443  (.A(\i55/n42 ),
    .B(\i55/n513 ),
    .Y(\i55/n75 ));
 AND2x4_ASAP7_75t_SL \i55/i444  (.A(\i55/n512 ),
    .B(\i55/n35 ),
    .Y(\i55/n72 ));
 AND2x4_ASAP7_75t_SL \i55/i445  (.A(\i55/n548 ),
    .B(\i55/n511 ),
    .Y(\i55/n71 ));
 AND2x4_ASAP7_75t_SL \i55/i446  (.A(\i55/n40 ),
    .B(\i55/n39 ),
    .Y(\i55/n70 ));
 OR2x6_ASAP7_75t_SL \i55/i447  (.A(\i55/n41 ),
    .B(\i55/n504 ),
    .Y(\i55/n68 ));
 INVx3_ASAP7_75t_SL \i55/i448  (.A(\i55/n65 ),
    .Y(\i55/n15 ));
 INVx3_ASAP7_75t_SL \i55/i449  (.A(\i55/n64 ),
    .Y(\i55/n63 ));
 NOR2xp33_ASAP7_75t_SL \i55/i45  (.A(\i55/n400 ),
    .B(\i55/n424 ),
    .Y(\i55/n455 ));
 INVx4_ASAP7_75t_SL \i55/i450  (.A(\i55/n14 ),
    .Y(\i55/n62 ));
 INVx4_ASAP7_75t_SL \i55/i451  (.A(\i55/n60 ),
    .Y(\i55/n59 ));
 INVx3_ASAP7_75t_SL \i55/i452  (.A(\i55/n58 ),
    .Y(\i55/n57 ));
 INVx4_ASAP7_75t_SL \i55/i453  (.A(\i55/n56 ),
    .Y(\i55/n55 ));
 INVx3_ASAP7_75t_SL \i55/i454  (.A(\i55/n54 ),
    .Y(\i55/n13 ));
 INVx4_ASAP7_75t_SL \i55/i455  (.A(\i55/n53 ),
    .Y(\i55/n52 ));
 INVx3_ASAP7_75t_SL \i55/i456  (.A(\i55/n49 ),
    .Y(\i55/n48 ));
 INVx3_ASAP7_75t_SL \i55/i457  (.A(\i55/n47 ),
    .Y(\i55/n46 ));
 INVx3_ASAP7_75t_SL \i55/i458  (.A(\i55/n45 ),
    .Y(\i55/n44 ));
 AND2x4_ASAP7_75t_SL \i55/i459  (.A(\i55/n40 ),
    .B(\i55/n533 ),
    .Y(\i55/n66 ));
 NAND3xp33_ASAP7_75t_SL \i55/i46  (.A(\i55/n391 ),
    .B(\i55/n398 ),
    .C(\i55/n517 ),
    .Y(\i55/n454 ));
 AND2x4_ASAP7_75t_SL \i55/i460  (.A(\i55/n38 ),
    .B(\i55/n508 ),
    .Y(\i55/n65 ));
 AND2x4_ASAP7_75t_SL \i55/i461  (.A(\i55/n5 ),
    .B(\i55/n39 ),
    .Y(\i55/n64 ));
 OR2x2_ASAP7_75t_SL \i55/i462  (.A(\i55/n10 ),
    .B(\i55/n509 ),
    .Y(\i55/n14 ));
 AND2x4_ASAP7_75t_SL \i55/i463  (.A(\i55/n532 ),
    .B(\i55/n38 ),
    .Y(\i55/n61 ));
 NAND2x1p5_ASAP7_75t_SL \i55/i464  (.A(\i55/n548 ),
    .B(\i55/n42 ),
    .Y(\i55/n60 ));
 AND2x4_ASAP7_75t_SL \i55/i465  (.A(\i55/n35 ),
    .B(\i55/n511 ),
    .Y(\i55/n58 ));
 OR2x2_ASAP7_75t_SL \i55/i466  (.A(\i55/n32 ),
    .B(\i55/n33 ),
    .Y(\i55/n56 ));
 AND2x4_ASAP7_75t_SL \i55/i467  (.A(\i55/n513 ),
    .B(\i55/n511 ),
    .Y(\i55/n54 ));
 AND2x4_ASAP7_75t_SL \i55/i468  (.A(\i55/n5 ),
    .B(\i55/n533 ),
    .Y(\i55/n53 ));
 AND2x4_ASAP7_75t_SL \i55/i469  (.A(\i55/n3 ),
    .B(\i55/n36 ),
    .Y(\i55/n51 ));
 NOR2x1_ASAP7_75t_SL \i55/i47  (.A(\i55/n348 ),
    .B(\i55/n409 ),
    .Y(\i55/n453 ));
 NAND2x1_ASAP7_75t_SL \i55/i470  (.A(\i55/n3 ),
    .B(\i55/n36 ),
    .Y(\i55/n50 ));
 AND2x4_ASAP7_75t_SL \i55/i471  (.A(\i55/n532 ),
    .B(\i55/n39 ),
    .Y(\i55/n49 ));
 AND2x4_ASAP7_75t_SL \i55/i472  (.A(\i55/n508 ),
    .B(\i55/n39 ),
    .Y(\i55/n47 ));
 OR2x6_ASAP7_75t_SL \i55/i473  (.A(\i55/n30 ),
    .B(\i55/n37 ),
    .Y(\i55/n45 ));
 INVx2_ASAP7_75t_SL \i55/i474  (.A(\i55/n42 ),
    .Y(\i55/n43 ));
 NAND2xp5_ASAP7_75t_SL \i55/i475  (.A(\i55/n11 ),
    .B(\i55/n1 ),
    .Y(\i55/n37 ));
 AND2x2_ASAP7_75t_SL \i55/i476  (.A(\i55/n11 ),
    .B(\i55/n1 ),
    .Y(\i55/n42 ));
 NAND2x1p5_ASAP7_75t_SL \i55/i477  (.A(n11[4]),
    .B(n11[5]),
    .Y(\i55/n41 ));
 AND2x2_ASAP7_75t_SL \i55/i478  (.A(\i55/n28 ),
    .B(\i55/n9 ),
    .Y(\i55/n40 ));
 AND2x2_ASAP7_75t_SL \i55/i479  (.A(n11[7]),
    .B(\i55/n12 ),
    .Y(\i55/n39 ));
 NOR2xp33_ASAP7_75t_SL \i55/i48  (.A(\i55/n531 ),
    .B(\i55/n327 ),
    .Y(\i55/n452 ));
 AND2x2_ASAP7_75t_SL \i55/i480  (.A(\i55/n0 ),
    .B(\i55/n12 ),
    .Y(\i55/n38 ));
 INVx2_ASAP7_75t_SL \i55/i481  (.A(\i55/n6 ),
    .Y(\i55/n36 ));
 INVx1_ASAP7_75t_SL \i55/i482  (.A(\i55/n35 ),
    .Y(\i55/n34 ));
 NAND2xp5_ASAP7_75t_SL \i55/i483  (.A(\i55/n29 ),
    .B(\i55/n2 ),
    .Y(\i55/n30 ));
 AND2x4_ASAP7_75t_SL \i55/i484  (.A(n11[0]),
    .B(\i55/n29 ),
    .Y(\i55/n35 ));
 NAND2xp5_ASAP7_75t_SL \i55/i485  (.A(\i55/n2 ),
    .B(n11[1]),
    .Y(\i55/n33 ));
 OR2x2_ASAP7_75t_SL \i55/i486  (.A(\i55/n1 ),
    .B(n11[3]),
    .Y(\i55/n32 ));
 NAND2x1_ASAP7_75t_SL \i55/i487  (.A(n11[3]),
    .B(\i55/n1 ),
    .Y(\i55/n31 ));
 INVx1_ASAP7_75t_SL \i55/i488  (.A(n11[1]),
    .Y(\i55/n29 ));
 INVx3_ASAP7_75t_SL \i55/i489  (.A(n11[5]),
    .Y(\i55/n28 ));
 NAND2xp5_ASAP7_75t_SL \i55/i49  (.A(\i55/n422 ),
    .B(\i55/n418 ),
    .Y(\i55/n451 ));
 INVx2_ASAP7_75t_SL \i55/i490  (.A(n11[6]),
    .Y(\i55/n12 ));
 INVx2_ASAP7_75t_SL \i55/i491  (.A(n11[3]),
    .Y(\i55/n11 ));
 INVx1_ASAP7_75t_SL \i55/i492  (.A(\i55/n421 ),
    .Y(\i55/n8 ));
 NAND2xp33_ASAP7_75t_SL \i55/i493  (.A(\i55/n0 ),
    .B(n11[6]),
    .Y(\i55/n10 ));
 INVx2_ASAP7_75t_SL \i55/i494  (.A(n11[4]),
    .Y(\i55/n9 ));
 OR2x2_ASAP7_75t_SL \i55/i495  (.A(\i55/n123 ),
    .B(\i55/n212 ),
    .Y(\i55/n7 ));
 OR2x2_ASAP7_75t_SL \i55/i496  (.A(n11[0]),
    .B(n11[1]),
    .Y(\i55/n6 ));
 NAND2x1p5_ASAP7_75t_SL \i55/i497  (.A(\i55/n3 ),
    .B(\i55/n35 ),
    .Y(\i55/n489 ));
 NAND2xp5_ASAP7_75t_SL \i55/i498  (.A(\i55/n4 ),
    .B(\i55/n527 ),
    .Y(\i55/n490 ));
 OAI31xp33_ASAP7_75t_SL \i55/i499  (.A1(\i55/n529 ),
    .A2(\i55/n4 ),
    .A3(\i55/n54 ),
    .B(\i55/n49 ),
    .Y(\i55/n491 ));
 INVx2_ASAP7_75t_SL \i55/i5  (.A(\i55/n41 ),
    .Y(\i55/n5 ));
 NOR2x1_ASAP7_75t_SL \i55/i50  (.A(\i55/n331 ),
    .B(\i55/n424 ),
    .Y(\i55/n450 ));
 AOI22xp5_ASAP7_75t_SL \i55/i500  (.A1(\i55/n528 ),
    .A2(\i55/n59 ),
    .B1(\i55/n49 ),
    .B2(\i55/n4 ),
    .Y(\i55/n492 ));
 NAND2xp5_ASAP7_75t_SL \i55/i501  (.A(\i55/n505 ),
    .B(\i55/n4 ),
    .Y(\i55/n493 ));
 AOI22xp5_ASAP7_75t_SL \i55/i502  (.A1(\i55/n527 ),
    .A2(\i55/n75 ),
    .B1(\i55/n507 ),
    .B2(\i55/n4 ),
    .Y(\i55/n494 ));
 NAND2xp33_ASAP7_75t_L \i55/i503  (.A(\i55/n4 ),
    .B(\i55/n507 ),
    .Y(\i55/n495 ));
 AOI22xp33_ASAP7_75t_SL \i55/i504  (.A1(\i55/n84 ),
    .A2(\i55/n55 ),
    .B1(\i55/n66 ),
    .B2(\i55/n4 ),
    .Y(\i55/n496 ));
 INVx3_ASAP7_75t_SL \i55/i505  (.A(\i55/n72 ),
    .Y(\i55/n497 ));
 INVx3_ASAP7_75t_SL \i55/i506  (.A(\i55/n61 ),
    .Y(\i55/n498 ));
 INVx2_ASAP7_75t_SL \i55/i507  (.A(\i55/n529 ),
    .Y(\i55/n499 ));
 INVx2_ASAP7_75t_SL \i55/i508  (.A(\i55/n66 ),
    .Y(\i55/n500 ));
 AO21x2_ASAP7_75t_SL \i55/i509  (.A1(\i55/n528 ),
    .A2(\i55/n4 ),
    .B(\i55/n501 ),
    .Y(\i55/n502 ));
 NOR2x1_ASAP7_75t_SL \i55/i51  (.A(\i55/n399 ),
    .B(\i55/n410 ),
    .Y(\i55/n449 ));
 OAI22xp5_ASAP7_75t_SL \i55/i510  (.A1(\i55/n497 ),
    .A2(\i55/n498 ),
    .B1(\i55/n499 ),
    .B2(\i55/n500 ),
    .Y(\i55/n501 ));
 INVx2_ASAP7_75t_SL \i55/i511  (.A(\i55/n503 ),
    .Y(\i55/n504 ));
 AND2x2_ASAP7_75t_SL \i55/i512  (.A(n11[7]),
    .B(n11[6]),
    .Y(\i55/n503 ));
 AND2x4_ASAP7_75t_SL \i55/i513  (.A(\i55/n503 ),
    .B(\i55/n508 ),
    .Y(\i55/n505 ));
 AOI211xp5_ASAP7_75t_SL \i55/i514  (.A1(\i55/n81 ),
    .A2(\i55/n503 ),
    .B(\i55/n110 ),
    .C(\i55/n117 ),
    .Y(\i55/n506 ));
 AND2x4_ASAP7_75t_SL \i55/i515  (.A(\i55/n503 ),
    .B(\i55/n532 ),
    .Y(\i55/n507 ));
 AND2x2_ASAP7_75t_SL \i55/i516  (.A(n11[5]),
    .B(\i55/n9 ),
    .Y(\i55/n508 ));
 NAND2xp5_ASAP7_75t_SL \i55/i517  (.A(n11[5]),
    .B(\i55/n9 ),
    .Y(\i55/n509 ));
 INVx3_ASAP7_75t_SL \i55/i518  (.A(\i55/n71 ),
    .Y(\i55/n510 ));
 INVx2_ASAP7_75t_SL \i55/i519  (.A(\i55/n31 ),
    .Y(\i55/n511 ));
 NAND2xp5_ASAP7_75t_SL \i55/i52  (.A(\i55/n363 ),
    .B(\i55/n404 ),
    .Y(\i55/n448 ));
 AND2x4_ASAP7_75t_SL \i55/i520  (.A(n11[3]),
    .B(n11[2]),
    .Y(\i55/n512 ));
 INVx2_ASAP7_75t_SL \i55/i521  (.A(\i55/n33 ),
    .Y(\i55/n513 ));
 INVx3_ASAP7_75t_SL \i55/i522  (.A(\i55/n514 ),
    .Y(\i55/n515 ));
 AND2x4_ASAP7_75t_SL \i55/i523  (.A(\i55/n512 ),
    .B(\i55/n513 ),
    .Y(\i55/n514 ));
 OAI21xp5_ASAP7_75t_SL \i55/i524  (.A1(\i55/n514 ),
    .A2(\i55/n58 ),
    .B(\i55/n49 ),
    .Y(\i55/n516 ));
 AOI211xp5_ASAP7_75t_SL \i55/i525  (.A1(\i55/n514 ),
    .A2(\i55/n67 ),
    .B(\i55/n164 ),
    .C(\i55/n502 ),
    .Y(\i55/n517 ));
 OAI21xp5_ASAP7_75t_SL \i55/i526  (.A1(\i55/n71 ),
    .A2(\i55/n514 ),
    .B(\i55/n84 ),
    .Y(\i55/n518 ));
 OAI21xp5_ASAP7_75t_SL \i55/i527  (.A1(\i55/n514 ),
    .A2(\i55/n59 ),
    .B(\i55/n507 ),
    .Y(\i55/n519 ));
 NAND2xp5_ASAP7_75t_SL \i55/i528  (.A(\i55/n61 ),
    .B(\i55/n514 ),
    .Y(\i55/n520 ));
 NAND2xp5_ASAP7_75t_SL \i55/i529  (.A(\i55/n53 ),
    .B(\i55/n514 ),
    .Y(\i55/n521 ));
 NOR5xp2_ASAP7_75t_SL \i55/i53  (.A(\i55/n288 ),
    .B(\i55/n26 ),
    .C(\i55/n301 ),
    .D(\i55/n530 ),
    .E(\i55/n265 ),
    .Y(\i55/n447 ));
 AND2x2_ASAP7_75t_SL \i55/i530  (.A(\i55/n505 ),
    .B(\i55/n514 ),
    .Y(\i55/n522 ));
 NAND2xp5_ASAP7_75t_SL \i55/i531  (.A(\i55/n64 ),
    .B(\i55/n514 ),
    .Y(\i55/n523 ));
 NAND2xp5_ASAP7_75t_SL \i55/i532  (.A(\i55/n47 ),
    .B(\i55/n514 ),
    .Y(\i55/n524 ));
 NOR2xp33_ASAP7_75t_SL \i55/i533  (.A(\i55/n514 ),
    .B(\i55/n77 ),
    .Y(\i55/n525 ));
 NOR2xp33_ASAP7_75t_SL \i55/i534  (.A(\i55/n514 ),
    .B(\i55/n58 ),
    .Y(\i55/n526 ));
 AND2x4_ASAP7_75t_SL \i55/i535  (.A(\i55/n38 ),
    .B(\i55/n5 ),
    .Y(\i55/n527 ));
 AND2x4_ASAP7_75t_SL \i55/i536  (.A(\i55/n503 ),
    .B(\i55/n40 ),
    .Y(\i55/n528 ));
 AND2x4_ASAP7_75t_SL \i55/i537  (.A(\i55/n548 ),
    .B(\i55/n512 ),
    .Y(\i55/n529 ));
 NAND2xp5_ASAP7_75t_SL \i55/i538  (.A(\i55/n233 ),
    .B(\i55/n550 ),
    .Y(\i55/n530 ));
 NAND3xp33_ASAP7_75t_SL \i55/i539  (.A(\i55/n296 ),
    .B(\i55/n491 ),
    .C(\i55/n550 ),
    .Y(\i55/n531 ));
 NOR2x1_ASAP7_75t_SL \i55/i54  (.A(\i55/n8 ),
    .B(\i55/n411 ),
    .Y(\i55/n446 ));
 AND2x2_ASAP7_75t_SL \i55/i540  (.A(n11[4]),
    .B(\i55/n28 ),
    .Y(\i55/n532 ));
 AND2x2_ASAP7_75t_SL \i55/i541  (.A(\i55/n0 ),
    .B(n11[6]),
    .Y(\i55/n533 ));
 OAI21xp5_ASAP7_75t_SL \i55/i542  (.A1(\i55/n534 ),
    .A2(\i55/n70 ),
    .B(\i55/n514 ),
    .Y(\i55/n535 ));
 AND2x4_ASAP7_75t_SL \i55/i543  (.A(\i55/n532 ),
    .B(\i55/n533 ),
    .Y(\i55/n534 ));
 NAND2xp5_ASAP7_75t_SL \i55/i544  (.A(\i55/n4 ),
    .B(\i55/n534 ),
    .Y(\i55/n536 ));
 INVx4_ASAP7_75t_SL \i55/i545  (.A(\i55/n534 ),
    .Y(\i55/n537 ));
 OAI21xp5_ASAP7_75t_SL \i55/i546  (.A1(\i55/n55 ),
    .A2(\i55/n51 ),
    .B(\i55/n534 ),
    .Y(\i55/n538 ));
 OAI21xp5_ASAP7_75t_SL \i55/i547  (.A1(\i55/n528 ),
    .A2(\i55/n534 ),
    .B(\i55/n55 ),
    .Y(\i55/n539 ));
 AOI22xp5_ASAP7_75t_SL \i55/i548  (.A1(\i55/n534 ),
    .A2(\i55/n77 ),
    .B1(\i55/n47 ),
    .B2(\i55/n59 ),
    .Y(\i55/n540 ));
 NAND2xp5_ASAP7_75t_SL \i55/i549  (.A(\i55/n534 ),
    .B(\i55/n71 ),
    .Y(\i55/n541 ));
 NAND2x1_ASAP7_75t_SL \i55/i55  (.A(\i55/n408 ),
    .B(\i55/n389 ),
    .Y(\i55/n459 ));
 NAND2xp5_ASAP7_75t_SL \i55/i550  (.A(\i55/n534 ),
    .B(\i55/n72 ),
    .Y(\i55/n542 ));
 NAND2xp5_ASAP7_75t_SL \i55/i551  (.A(\i55/n534 ),
    .B(\i55/n54 ),
    .Y(\i55/n543 ));
 NAND2xp5_ASAP7_75t_SL \i55/i552  (.A(\i55/n534 ),
    .B(\i55/n75 ),
    .Y(\i55/n544 ));
 NAND2x1_ASAP7_75t_SL \i55/i553  (.A(\i55/n534 ),
    .B(\i55/n79 ),
    .Y(\i55/n545 ));
 OR2x2_ASAP7_75t_SL \i55/i554  (.A(\i55/n289 ),
    .B(\i55/n378 ),
    .Y(\i55/n546 ));
 NOR2xp33_ASAP7_75t_SL \i55/i555  (.A(\i55/n289 ),
    .B(\i55/n378 ),
    .Y(\i55/n547 ));
 AND2x2_ASAP7_75t_SL \i55/i556  (.A(n11[0]),
    .B(n11[1]),
    .Y(\i55/n548 ));
 AOI22xp5_ASAP7_75t_SL \i55/i557  (.A1(\i55/n549 ),
    .A2(\i55/n527 ),
    .B1(\i55/n528 ),
    .B2(\i55/n529 ),
    .Y(\i55/n550 ));
 AND2x4_ASAP7_75t_SL \i55/i558  (.A(\i55/n548 ),
    .B(\i55/n3 ),
    .Y(\i55/n549 ));
 NOR2xp33_ASAP7_75t_SL \i55/i559  (.A(\i55/n549 ),
    .B(\i55/n4 ),
    .Y(\i55/n551 ));
 NOR2x1_ASAP7_75t_SL \i55/i56  (.A(\i55/n425 ),
    .B(\i55/n410 ),
    .Y(\i55/n445 ));
 INVx3_ASAP7_75t_SL \i55/i560  (.A(\i55/n549 ),
    .Y(\i55/n552 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i55/i561  (.A1(\i55/n549 ),
    .A2(\i55/n51 ),
    .B(\i55/n70 ),
    .C(\i55/n566 ),
    .Y(\i55/n553 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i55/i562  (.A1(\i55/n505 ),
    .A2(\i55/n62 ),
    .B(\i55/n549 ),
    .C(\i55/n18 ),
    .Y(\i55/n554 ));
 AOI21xp5_ASAP7_75t_SL \i55/i563  (.A1(\i55/n152 ),
    .A2(\i55/n549 ),
    .B(\i55/n225 ),
    .Y(\i55/n555 ));
 AOI22xp5_ASAP7_75t_SL \i55/i564  (.A1(\i55/n79 ),
    .A2(\i55/n149 ),
    .B1(\i55/n61 ),
    .B2(\i55/n549 ),
    .Y(\i55/n556 ));
 OA21x2_ASAP7_75t_SL \i55/i565  (.A1(\i55/n62 ),
    .A2(\i55/n84 ),
    .B(\i55/n549 ),
    .Y(\i55/n557 ));
 OAI21xp5_ASAP7_75t_SL \i55/i566  (.A1(\i55/n549 ),
    .A2(\i55/n71 ),
    .B(\i55/n49 ),
    .Y(\i55/n558 ));
 AOI22xp5_ASAP7_75t_SL \i55/i567  (.A1(\i55/n49 ),
    .A2(\i55/n59 ),
    .B1(\i55/n47 ),
    .B2(\i55/n549 ),
    .Y(\i55/n559 ));
 NAND2xp5_ASAP7_75t_SL \i55/i568  (.A(\i55/n505 ),
    .B(\i55/n549 ),
    .Y(\i55/n560 ));
 NAND2xp5_ASAP7_75t_SL \i55/i569  (.A(\i55/n67 ),
    .B(\i55/n549 ),
    .Y(\i55/n561 ));
 NOR2x1_ASAP7_75t_SL \i55/i57  (.A(\i55/n347 ),
    .B(\i55/n409 ),
    .Y(\i55/n458 ));
 NAND2xp5_ASAP7_75t_SL \i55/i570  (.A(\i55/n507 ),
    .B(\i55/n549 ),
    .Y(\i55/n562 ));
 NAND2xp5_ASAP7_75t_SL \i55/i571  (.A(\i55/n549 ),
    .B(\i55/n65 ),
    .Y(\i55/n563 ));
 NOR2xp33_ASAP7_75t_SL \i55/i572  (.A(\i55/n549 ),
    .B(\i55/n75 ),
    .Y(\i55/n564 ));
 NAND2xp5_ASAP7_75t_SL \i55/i573  (.A(\i55/n528 ),
    .B(\i55/n549 ),
    .Y(\i55/n565 ));
 AND2x2_ASAP7_75t_SL \i55/i574  (.A(\i55/n62 ),
    .B(\i55/n72 ),
    .Y(\i55/n566 ));
 NAND2xp5_ASAP7_75t_SL \i55/i575  (.A(\i55/n272 ),
    .B(\i55/n568 ),
    .Y(\i55/n569 ));
 NOR2xp67_ASAP7_75t_SL \i55/i576  (.A(\i55/n566 ),
    .B(\i55/n567 ),
    .Y(\i55/n568 ));
 OAI22xp33_ASAP7_75t_SL \i55/i577  (.A1(\i55/n82 ),
    .A2(\i55/n52 ),
    .B1(\i55/n48 ),
    .B2(\i55/n13 ),
    .Y(\i55/n567 ));
 NAND5xp2_ASAP7_75t_SL \i55/i578  (.A(\i55/n568 ),
    .B(\i55/n341 ),
    .C(\i55/n199 ),
    .D(\i55/n544 ),
    .E(\i55/n177 ),
    .Y(\i55/n570 ));
 AOI211x1_ASAP7_75t_SL \i55/i579  (.A1(\i55/n44 ),
    .A2(\i55/n70 ),
    .B(\i55/n110 ),
    .C(\i55/n546 ),
    .Y(\i55/n571 ));
 INVxp67_ASAP7_75t_SL \i55/i58  (.A(\i55/n443 ),
    .Y(\i55/n444 ));
 AND4x1_ASAP7_75t_SL \i55/i580  (.A(\i55/n287 ),
    .B(\i55/n329 ),
    .C(\i55/n581 ),
    .D(\i55/n259 ),
    .Y(\i55/n572 ));
 NOR3xp33_ASAP7_75t_SL \i55/i581  (.A(\i55/n573 ),
    .B(\i55/n317 ),
    .C(\i55/n136 ),
    .Y(\i55/n574 ));
 OAI21xp5_ASAP7_75t_SL \i55/i582  (.A1(\i55/n69 ),
    .A2(\i55/n74 ),
    .B(\i55/n156 ),
    .Y(\i55/n573 ));
 NAND3xp33_ASAP7_75t_SL \i55/i583  (.A(\i55/n575 ),
    .B(\i55/n252 ),
    .C(\i55/n321 ),
    .Y(\i55/n576 ));
 AO21x1_ASAP7_75t_SL \i55/i584  (.A1(\i55/n500 ),
    .A2(\i55/n52 ),
    .B(\i55/n552 ),
    .Y(\i55/n575 ));
 NAND2xp33_ASAP7_75t_SL \i55/i585  (.A(\i55/n577 ),
    .B(\i55/n290 ),
    .Y(\i55/n578 ));
 OAI21xp5_ASAP7_75t_SL \i55/i586  (.A1(\i55/n4 ),
    .A2(\i55/n71 ),
    .B(\i55/n47 ),
    .Y(\i55/n577 ));
 NOR3xp33_ASAP7_75t_SL \i55/i587  (.A(\i55/n579 ),
    .B(\i55/n319 ),
    .C(\i55/n501 ),
    .Y(\i55/n580 ));
 OAI21xp5_ASAP7_75t_SL \i55/i588  (.A1(\i55/n68 ),
    .A2(\i55/n16 ),
    .B(\i55/n536 ),
    .Y(\i55/n579 ));
 AOI21xp5_ASAP7_75t_SL \i55/i589  (.A1(\i55/n53 ),
    .A2(\i55/n529 ),
    .B(\i55/n200 ),
    .Y(\i55/n581 ));
 INVxp67_ASAP7_75t_SL \i55/i59  (.A(\i55/n439 ),
    .Y(\i55/n440 ));
 NOR2x1p5_ASAP7_75t_SL \i55/i6  (.A(\i55/n484 ),
    .B(\i55/n483 ),
    .Y(n10[4]));
 AND5x1_ASAP7_75t_SL \i55/i60  (.A(\i55/n359 ),
    .B(\i55/n581 ),
    .C(\i55/n352 ),
    .D(\i55/n275 ),
    .E(\i55/n245 ),
    .Y(\i55/n438 ));
 NOR3xp33_ASAP7_75t_SL \i55/i61  (.A(\i55/n370 ),
    .B(\i55/n351 ),
    .C(\i55/n333 ),
    .Y(\i55/n437 ));
 NOR3xp33_ASAP7_75t_SL \i55/i62  (.A(\i55/n397 ),
    .B(\i55/n334 ),
    .C(\i55/n285 ),
    .Y(\i55/n436 ));
 AND5x1_ASAP7_75t_SL \i55/i63  (.A(\i55/n323 ),
    .B(\i55/n337 ),
    .C(\i55/n506 ),
    .D(\i55/n326 ),
    .E(\i55/n254 ),
    .Y(\i55/n435 ));
 NOR2xp33_ASAP7_75t_SL \i55/i64  (.A(\i55/n570 ),
    .B(\i55/n402 ),
    .Y(\i55/n434 ));
 NAND4xp25_ASAP7_75t_SL \i55/i65  (.A(\i55/n380 ),
    .B(\i55/n388 ),
    .C(\i55/n393 ),
    .D(\i55/n376 ),
    .Y(\i55/n433 ));
 NAND5xp2_ASAP7_75t_SL \i55/i66  (.A(\i55/n358 ),
    .B(\i55/n316 ),
    .C(\i55/n218 ),
    .D(\i55/n204 ),
    .E(\i55/n297 ),
    .Y(\i55/n432 ));
 NOR4xp25_ASAP7_75t_SL \i55/i67  (.A(\i55/n349 ),
    .B(\i55/n26 ),
    .C(\i55/n302 ),
    .D(\i55/n279 ),
    .Y(\i55/n431 ));
 NAND4xp25_ASAP7_75t_SL \i55/i68  (.A(\i55/n366 ),
    .B(\i55/n382 ),
    .C(\i55/n385 ),
    .D(\i55/n387 ),
    .Y(\i55/n430 ));
 NAND4xp25_ASAP7_75t_SL \i55/i69  (.A(\i55/n395 ),
    .B(\i55/n393 ),
    .C(\i55/n184 ),
    .D(\i55/n244 ),
    .Y(\i55/n429 ));
 NOR2x2_ASAP7_75t_SL \i55/i7  (.A(\i55/n479 ),
    .B(\i55/n485 ),
    .Y(n10[3]));
 NAND3xp33_ASAP7_75t_SL \i55/i70  (.A(\i55/n387 ),
    .B(\i55/n357 ),
    .C(\i55/n19 ),
    .Y(\i55/n443 ));
 NAND4xp75_ASAP7_75t_SL \i55/i71  (.A(\i55/n293 ),
    .B(\i55/n264 ),
    .C(\i55/n346 ),
    .D(\i55/n23 ),
    .Y(\i55/n442 ));
 NAND2xp33_ASAP7_75t_L \i55/i72  (.A(\i55/n365 ),
    .B(\i55/n426 ),
    .Y(\i55/n428 ));
 AND2x2_ASAP7_75t_SL \i55/i73  (.A(\i55/n368 ),
    .B(\i55/n416 ),
    .Y(\i55/n441 ));
 NAND2x1p5_ASAP7_75t_SL \i55/i74  (.A(\i55/n423 ),
    .B(\i55/n381 ),
    .Y(\i55/n439 ));
 INVxp67_ASAP7_75t_SL \i55/i75  (.A(\i55/n426 ),
    .Y(\i55/n427 ));
 NOR5xp2_ASAP7_75t_SL \i55/i76  (.A(\i55/n311 ),
    .B(\i55/n284 ),
    .C(\i55/n210 ),
    .D(\i55/n175 ),
    .E(\i55/n89 ),
    .Y(\i55/n419 ));
 NOR3xp33_ASAP7_75t_SL \i55/i77  (.A(\i55/n392 ),
    .B(\i55/n307 ),
    .C(\i55/n300 ),
    .Y(\i55/n418 ));
 NOR2xp33_ASAP7_75t_SL \i55/i78  (.A(\i55/n578 ),
    .B(\i55/n367 ),
    .Y(\i55/n417 ));
 NOR2xp33_ASAP7_75t_SL \i55/i79  (.A(\i55/n390 ),
    .B(\i55/n339 ),
    .Y(\i55/n416 ));
 AND5x2_ASAP7_75t_SL \i55/i8  (.A(\i55/n477 ),
    .B(\i55/n468 ),
    .C(\i55/n470 ),
    .D(\i55/n455 ),
    .E(\i55/n447 ),
    .Y(n10[6]));
 NOR2x1_ASAP7_75t_SL \i55/i80  (.A(\i55/n353 ),
    .B(\i55/n324 ),
    .Y(\i55/n426 ));
 NAND2xp5_ASAP7_75t_SL \i55/i81  (.A(\i55/n389 ),
    .B(\i55/n356 ),
    .Y(\i55/n415 ));
 NAND2xp5_ASAP7_75t_SL \i55/i82  (.A(\i55/n379 ),
    .B(\i55/n338 ),
    .Y(\i55/n414 ));
 NAND3xp33_ASAP7_75t_SL \i55/i83  (.A(\i55/n581 ),
    .B(\i55/n281 ),
    .C(\i55/n259 ),
    .Y(\i55/n425 ));
 NOR3xp33_ASAP7_75t_SL \i55/i84  (.A(\i55/n360 ),
    .B(\i55/n7 ),
    .C(\i55/n261 ),
    .Y(\i55/n413 ));
 NAND2xp5_ASAP7_75t_SL \i55/i85  (.A(\i55/n21 ),
    .B(\i55/n366 ),
    .Y(\i55/n424 ));
 OR3x1_ASAP7_75t_SL \i55/i86  (.A(\i55/n288 ),
    .B(\i55/n301 ),
    .C(\i55/n530 ),
    .Y(\i55/n412 ));
 NOR2x1_ASAP7_75t_SL \i55/i87  (.A(\i55/n300 ),
    .B(\i55/n392 ),
    .Y(\i55/n423 ));
 NOR2xp33_ASAP7_75t_L \i55/i88  (.A(\i55/n350 ),
    .B(\i55/n336 ),
    .Y(\i55/n422 ));
 NOR3x1_ASAP7_75t_SL \i55/i89  (.A(\i55/n295 ),
    .B(\i55/n189 ),
    .C(\i55/n343 ),
    .Y(\i55/n421 ));
 AND3x4_ASAP7_75t_SL \i55/i9  (.A(\i55/n477 ),
    .B(\i55/n486 ),
    .C(\i55/n465 ),
    .Y(n10[1]));
 NOR2xp67_ASAP7_75t_SL \i55/i90  (.A(\i55/n375 ),
    .B(\i55/n369 ),
    .Y(\i55/n420 ));
 NOR3xp33_ASAP7_75t_SL \i55/i91  (.A(\i55/n303 ),
    .B(\i55/n217 ),
    .C(\i55/n292 ),
    .Y(\i55/n408 ));
 NOR2xp33_ASAP7_75t_SL \i55/i92  (.A(\i55/n576 ),
    .B(\i55/n362 ),
    .Y(\i55/n407 ));
 NAND3xp33_ASAP7_75t_SL \i55/i93  (.A(\i55/n287 ),
    .B(\i55/n354 ),
    .C(\i55/n556 ),
    .Y(\i55/n406 ));
 NAND4xp25_ASAP7_75t_SL \i55/i94  (.A(\i55/n270 ),
    .B(\i55/n553 ),
    .C(\i55/n312 ),
    .D(\i55/n280 ),
    .Y(\i55/n405 ));
 NAND2x1_ASAP7_75t_SL \i55/i95  (.A(\i55/n377 ),
    .B(\i55/n391 ),
    .Y(\i55/n411 ));
 NOR5xp2_ASAP7_75t_SL \i55/i96  (.A(\i55/n386 ),
    .B(\i55/n305 ),
    .C(\i55/n122 ),
    .D(\i55/n229 ),
    .E(\i55/n157 ),
    .Y(\i55/n404 ));
 NAND3xp33_ASAP7_75t_SL \i55/i97  (.A(\i55/n342 ),
    .B(\i55/n574 ),
    .C(\i55/n220 ),
    .Y(\i55/n403 ));
 NAND2xp33_ASAP7_75t_SL \i55/i98  (.A(\i55/n555 ),
    .B(\i55/n383 ),
    .Y(\i55/n402 ));
 NOR5xp2_ASAP7_75t_SL \i55/i99  (.A(\i55/n325 ),
    .B(\i55/n289 ),
    .C(\i55/n310 ),
    .D(\i55/n255 ),
    .E(\i55/n208 ),
    .Y(\i55/n401 ));
 OAI22xp5_ASAP7_75t_SL i550 (.A1(n583),
    .A2(n487),
    .B1(n582),
    .B2(n486),
    .Y(n922));
 AOI22xp5_ASAP7_75t_SL i551 (.A1(n579),
    .A2(n783),
    .B1(n580),
    .B2(n784),
    .Y(n921));
 OAI22xp5_ASAP7_75t_SL i552 (.A1(n562),
    .A2(n791),
    .B1(n561),
    .B2(n790),
    .Y(n920));
 AOI22xp5_ASAP7_75t_SL i553 (.A1(n483),
    .A2(n217),
    .B1(n482),
    .B2(n533),
    .Y(n919));
 AOI22xp5_ASAP7_75t_SL i554 (.A1(n786),
    .A2(n523),
    .B1(n785),
    .B2(n524),
    .Y(n918));
 AOI22xp5_ASAP7_75t_SL i555 (.A1(n548),
    .A2(n488),
    .B1(n549),
    .B2(n489),
    .Y(n917));
 OAI22xp5_ASAP7_75t_SL i556 (.A1(n556),
    .A2(n809),
    .B1(n810),
    .B2(n555),
    .Y(n916));
 AOI22xp5_ASAP7_75t_SL i557 (.A1(n807),
    .A2(n125),
    .B1(n808),
    .B2(n475),
    .Y(n915));
 AOI22xp33_ASAP7_75t_SL i558 (.A1(n477),
    .A2(n223),
    .B1(n778),
    .B2(n478),
    .Y(n914));
 OAI22xp5_ASAP7_75t_SL i559 (.A1(n500),
    .A2(n764),
    .B1(n499),
    .B2(n765),
    .Y(n913));
 INVx1_ASAP7_75t_SL \i56/i0  (.A(n9[5]),
    .Y(\i56/n0 ));
 INVx2_ASAP7_75t_SL \i56/i1  (.A(\i56/n62 ),
    .Y(\i56/n1 ));
 NAND4xp25_ASAP7_75t_SL \i56/i10  (.A(\i56/n457 ),
    .B(\i56/n393 ),
    .C(\i56/n382 ),
    .D(\i56/n398 ),
    .Y(\i56/n481 ));
 NOR2xp33_ASAP7_75t_SL \i56/i100  (.A(\i56/n332 ),
    .B(\i56/n364 ),
    .Y(\i56/n391 ));
 NAND2xp5_ASAP7_75t_SL \i56/i101  (.A(\i56/n350 ),
    .B(\i56/n386 ),
    .Y(\i56/n400 ));
 INVxp33_ASAP7_75t_SL \i56/i102  (.A(\i56/n388 ),
    .Y(\i56/n389 ));
 INVxp67_ASAP7_75t_SL \i56/i103  (.A(\i56/n384 ),
    .Y(\i56/n385 ));
 NOR3xp33_ASAP7_75t_SL \i56/i104  (.A(\i56/n251 ),
    .B(\i56/n212 ),
    .C(\i56/n91 ),
    .Y(\i56/n380 ));
 OAI211xp5_ASAP7_75t_SL \i56/i105  (.A1(\i56/n66 ),
    .A2(\i56/n177 ),
    .B(\i56/n498 ),
    .C(\i56/n291 ),
    .Y(\i56/n379 ));
 NOR2xp33_ASAP7_75t_SL \i56/i106  (.A(\i56/n331 ),
    .B(\i56/n14 ),
    .Y(\i56/n378 ));
 OAI21xp5_ASAP7_75t_SL \i56/i107  (.A1(\i56/n57 ),
    .A2(\i56/n79 ),
    .B(\i56/n334 ),
    .Y(\i56/n377 ));
 NOR4xp25_ASAP7_75t_SL \i56/i108  (.A(\i56/n235 ),
    .B(\i56/n236 ),
    .C(\i56/n203 ),
    .D(\i56/n227 ),
    .Y(\i56/n376 ));
 NAND2xp33_ASAP7_75t_SL \i56/i109  (.A(\i56/n554 ),
    .B(\i56/n336 ),
    .Y(\i56/n375 ));
 NOR3xp33_ASAP7_75t_SL \i56/i11  (.A(\i56/n440 ),
    .B(\i56/n470 ),
    .C(\i56/n453 ),
    .Y(\i56/n480 ));
 NOR3xp33_ASAP7_75t_SL \i56/i110  (.A(\i56/n511 ),
    .B(\i56/n131 ),
    .C(\i56/n187 ),
    .Y(\i56/n374 ));
 NAND2xp5_ASAP7_75t_SL \i56/i111  (.A(\i56/n222 ),
    .B(\i56/n500 ),
    .Y(\i56/n373 ));
 NOR2xp33_ASAP7_75t_L \i56/i112  (.A(\i56/n276 ),
    .B(\i56/n299 ),
    .Y(\i56/n390 ));
 OAI211xp5_ASAP7_75t_SL \i56/i113  (.A1(\i56/n45 ),
    .A2(\i56/n57 ),
    .B(\i56/n225 ),
    .C(\i56/n216 ),
    .Y(\i56/n372 ));
 NAND3xp33_ASAP7_75t_L \i56/i114  (.A(\i56/n253 ),
    .B(\i56/n522 ),
    .C(\i56/n301 ),
    .Y(\i56/n371 ));
 NAND2xp5_ASAP7_75t_SL \i56/i115  (.A(\i56/n499 ),
    .B(\i56/n225 ),
    .Y(\i56/n370 ));
 NAND2xp5_ASAP7_75t_L \i56/i116  (.A(\i56/n245 ),
    .B(\i56/n263 ),
    .Y(\i56/n369 ));
 NOR3xp33_ASAP7_75t_SL \i56/i117  (.A(\i56/n296 ),
    .B(\i56/n204 ),
    .C(\i56/n220 ),
    .Y(\i56/n368 ));
 NOR3xp33_ASAP7_75t_SL \i56/i118  (.A(\i56/n13 ),
    .B(\i56/n195 ),
    .C(\i56/n182 ),
    .Y(\i56/n367 ));
 NOR4xp25_ASAP7_75t_SL \i56/i119  (.A(\i56/n13 ),
    .B(\i56/n205 ),
    .C(\i56/n198 ),
    .D(\i56/n94 ),
    .Y(\i56/n366 ));
 AND2x2_ASAP7_75t_SL \i56/i12  (.A(\i56/n475 ),
    .B(\i56/n476 ),
    .Y(n8[2]));
 AOI211x1_ASAP7_75t_SL \i56/i120  (.A1(\i56/n111 ),
    .A2(\i56/n75 ),
    .B(\i56/n232 ),
    .C(\i56/n223 ),
    .Y(\i56/n388 ));
 NOR3xp33_ASAP7_75t_SL \i56/i121  (.A(\i56/n258 ),
    .B(\i56/n131 ),
    .C(\i56/n239 ),
    .Y(\i56/n387 ));
 NOR2xp33_ASAP7_75t_L \i56/i122  (.A(\i56/n220 ),
    .B(\i56/n340 ),
    .Y(\i56/n365 ));
 NOR2x1_ASAP7_75t_SL \i56/i123  (.A(\i56/n264 ),
    .B(\i56/n328 ),
    .Y(\i56/n386 ));
 NOR2xp33_ASAP7_75t_SL \i56/i124  (.A(\i56/n269 ),
    .B(\i56/n335 ),
    .Y(\i56/n384 ));
 NAND2xp5_ASAP7_75t_SL \i56/i125  (.A(\i56/n216 ),
    .B(\i56/n539 ),
    .Y(\i56/n383 ));
 NOR2xp67_ASAP7_75t_SL \i56/i126  (.A(\i56/n314 ),
    .B(\i56/n337 ),
    .Y(\i56/n382 ));
 NOR3x1_ASAP7_75t_SL \i56/i127  (.A(\i56/n512 ),
    .B(\i56/n251 ),
    .C(\i56/n509 ),
    .Y(\i56/n381 ));
 INVx1_ASAP7_75t_SL \i56/i128  (.A(\i56/n360 ),
    .Y(\i56/n361 ));
 NOR2xp33_ASAP7_75t_SL \i56/i129  (.A(\i56/n502 ),
    .B(\i56/n309 ),
    .Y(\i56/n358 ));
 NOR3xp33_ASAP7_75t_SL \i56/i13  (.A(\i56/n454 ),
    .B(\i56/n400 ),
    .C(\i56/n458 ),
    .Y(\i56/n479 ));
 NAND5xp2_ASAP7_75t_SL \i56/i130  (.A(\i56/n92 ),
    .B(\i56/n199 ),
    .C(\i56/n166 ),
    .D(\i56/n168 ),
    .E(\i56/n193 ),
    .Y(\i56/n357 ));
 NOR2xp33_ASAP7_75t_SL \i56/i131  (.A(\i56/n310 ),
    .B(\i56/n323 ),
    .Y(\i56/n356 ));
 OAI211xp5_ASAP7_75t_SL \i56/i132  (.A1(\i56/n45 ),
    .A2(\i56/n180 ),
    .B(\i56/n538 ),
    .C(\i56/n257 ),
    .Y(\i56/n355 ));
 A2O1A1Ixp33_ASAP7_75t_R \i56/i133  (.A1(\i56/n76 ),
    .A2(\i56/n194 ),
    .B(\i56/n4 ),
    .C(\i56/n249 ),
    .Y(\i56/n354 ));
 NAND3xp33_ASAP7_75t_SL \i56/i134  (.A(\i56/n520 ),
    .B(\i56/n240 ),
    .C(\i56/n233 ),
    .Y(\i56/n353 ));
 OAI21xp5_ASAP7_75t_SL \i56/i135  (.A1(\i56/n55 ),
    .A2(\i56/n501 ),
    .B(\i56/n551 ),
    .Y(\i56/n364 ));
 NOR3xp33_ASAP7_75t_SL \i56/i136  (.A(\i56/n266 ),
    .B(\i56/n219 ),
    .C(\i56/n224 ),
    .Y(\i56/n352 ));
 NAND3xp33_ASAP7_75t_L \i56/i137  (.A(\i56/n218 ),
    .B(\i56/n216 ),
    .C(\i56/n303 ),
    .Y(\i56/n351 ));
 NOR3xp33_ASAP7_75t_SL \i56/i138  (.A(\i56/n279 ),
    .B(\i56/n255 ),
    .C(\i56/n219 ),
    .Y(\i56/n350 ));
 AOI211xp5_ASAP7_75t_SL \i56/i139  (.A1(\i56/n71 ),
    .A2(\i56/n82 ),
    .B(\i56/n321 ),
    .C(\i56/n132 ),
    .Y(\i56/n349 ));
 NOR3xp33_ASAP7_75t_SL \i56/i14  (.A(\i56/n432 ),
    .B(\i56/n437 ),
    .C(\i56/n415 ),
    .Y(\i56/n478 ));
 OAI221xp5_ASAP7_75t_SL \i56/i140  (.A1(\i56/n177 ),
    .A2(\i56/n45 ),
    .B1(\i56/n118 ),
    .B2(\i56/n61 ),
    .C(\i56/n186 ),
    .Y(\i56/n348 ));
 AOI211xp5_ASAP7_75t_SL \i56/i141  (.A1(\i56/n84 ),
    .A2(\i56/n44 ),
    .B(\i56/n252 ),
    .C(\i56/n259 ),
    .Y(\i56/n347 ));
 NAND2xp33_ASAP7_75t_SL \i56/i142  (.A(\i56/n277 ),
    .B(\i56/n274 ),
    .Y(\i56/n346 ));
 NOR2xp33_ASAP7_75t_SL \i56/i143  (.A(\i56/n320 ),
    .B(\i56/n285 ),
    .Y(\i56/n345 ));
 NAND4xp25_ASAP7_75t_SL \i56/i144  (.A(\i56/n11 ),
    .B(\i56/n114 ),
    .C(\i56/n529 ),
    .D(\i56/n150 ),
    .Y(\i56/n344 ));
 OAI221xp5_ASAP7_75t_SL \i56/i145  (.A1(\i56/n241 ),
    .A2(\i56/n88 ),
    .B1(\i56/n8 ),
    .B2(\i56/n549 ),
    .C(\i56/n535 ),
    .Y(\i56/n343 ));
 NAND4xp25_ASAP7_75t_SL \i56/i146  (.A(\i56/n524 ),
    .B(\i56/n211 ),
    .C(\i56/n188 ),
    .D(\i56/n494 ),
    .Y(\i56/n342 ));
 NOR2xp33_ASAP7_75t_SL \i56/i147  (.A(\i56/n287 ),
    .B(\i56/n297 ),
    .Y(\i56/n363 ));
 NAND2xp33_ASAP7_75t_L \i56/i148  (.A(\i56/n327 ),
    .B(\i56/n228 ),
    .Y(\i56/n341 ));
 NOR2xp33_ASAP7_75t_SL \i56/i149  (.A(\i56/n306 ),
    .B(\i56/n324 ),
    .Y(\i56/n362 ));
 NOR3xp33_ASAP7_75t_SL \i56/i15  (.A(\i56/n443 ),
    .B(\i56/n445 ),
    .C(\i56/n427 ),
    .Y(\i56/n477 ));
 NAND2x1_ASAP7_75t_SL \i56/i150  (.A(\i56/n268 ),
    .B(\i56/n217 ),
    .Y(\i56/n360 ));
 NOR3xp33_ASAP7_75t_SL \i56/i151  (.A(\i56/n227 ),
    .B(\i56/n209 ),
    .C(\i56/n544 ),
    .Y(\i56/n359 ));
 NOR2xp67_ASAP7_75t_SL \i56/i152  (.A(\i56/n267 ),
    .B(\i56/n275 ),
    .Y(\i56/n15 ));
 INVxp67_ASAP7_75t_SL \i56/i153  (.A(\i56/n337 ),
    .Y(\i56/n338 ));
 INVxp33_ASAP7_75t_SL \i56/i154  (.A(\i56/n335 ),
    .Y(\i56/n336 ));
 INVx1_ASAP7_75t_SL \i56/i155  (.A(\i56/n332 ),
    .Y(\i56/n333 ));
 INVxp67_ASAP7_75t_SL \i56/i156  (.A(\i56/n328 ),
    .Y(\i56/n329 ));
 INVxp67_ASAP7_75t_SL \i56/i157  (.A(\i56/n14 ),
    .Y(\i56/n327 ));
 INVxp67_ASAP7_75t_SL \i56/i158  (.A(\i56/n325 ),
    .Y(\i56/n326 ));
 NAND2xp5_ASAP7_75t_SL \i56/i159  (.A(\i56/n522 ),
    .B(\i56/n523 ),
    .Y(\i56/n324 ));
 NOR4xp25_ASAP7_75t_SL \i56/i16  (.A(\i56/n424 ),
    .B(\i56/n412 ),
    .C(\i56/n416 ),
    .D(\i56/n426 ),
    .Y(\i56/n476 ));
 NAND2xp33_ASAP7_75t_SL \i56/i160  (.A(\i56/n486 ),
    .B(\i56/n243 ),
    .Y(\i56/n323 ));
 AOI21xp5_ASAP7_75t_SL \i56/i161  (.A1(\i56/n184 ),
    .A2(\i56/n89 ),
    .B(\i56/n255 ),
    .Y(\i56/n322 ));
 OAI22xp5_ASAP7_75t_SL \i56/i162  (.A1(\i56/n109 ),
    .A2(\i56/n146 ),
    .B1(\i56/n86 ),
    .B2(\i56/n129 ),
    .Y(\i56/n321 ));
 NAND4xp25_ASAP7_75t_SL \i56/i163  (.A(\i56/n190 ),
    .B(\i56/n141 ),
    .C(\i56/n140 ),
    .D(\i56/n115 ),
    .Y(\i56/n320 ));
 NAND3xp33_ASAP7_75t_SL \i56/i164  (.A(\i56/n137 ),
    .B(\i56/n149 ),
    .C(\i56/n5 ),
    .Y(\i56/n319 ));
 NAND3xp33_ASAP7_75t_SL \i56/i165  (.A(\i56/n176 ),
    .B(\i56/n189 ),
    .C(\i56/n548 ),
    .Y(\i56/n318 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i56/i166  (.A1(\i56/n47 ),
    .A2(\i56/n42 ),
    .B(\i56/n84 ),
    .C(\i56/n223 ),
    .Y(\i56/n317 ));
 NOR2xp33_ASAP7_75t_SL \i56/i167  (.A(\i56/n509 ),
    .B(\i56/n234 ),
    .Y(\i56/n316 ));
 OAI21xp5_ASAP7_75t_SL \i56/i168  (.A1(\i56/n86 ),
    .A2(\i56/n157 ),
    .B(\i56/n99 ),
    .Y(\i56/n315 ));
 NAND4xp25_ASAP7_75t_SL \i56/i169  (.A(\i56/n201 ),
    .B(\i56/n151 ),
    .C(\i56/n138 ),
    .D(\i56/n525 ),
    .Y(\i56/n314 ));
 NOR5xp2_ASAP7_75t_SL \i56/i17  (.A(\i56/n452 ),
    .B(\i56/n421 ),
    .C(\i56/n454 ),
    .D(\i56/n404 ),
    .E(\i56/n385 ),
    .Y(\i56/n475 ));
 AOI211xp5_ASAP7_75t_SL \i56/i170  (.A1(\i56/n42 ),
    .A2(\i56/n1 ),
    .B(\i56/n148 ),
    .C(\i56/n143 ),
    .Y(\i56/n313 ));
 NOR2xp33_ASAP7_75t_L \i56/i171  (.A(\i56/n208 ),
    .B(\i56/n247 ),
    .Y(\i56/n312 ));
 NOR2xp33_ASAP7_75t_L \i56/i172  (.A(\i56/n207 ),
    .B(\i56/n226 ),
    .Y(\i56/n311 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i56/i173  (.A1(\i56/n66 ),
    .A2(\i56/n41 ),
    .B(\i56/n50 ),
    .C(\i56/n250 ),
    .Y(\i56/n310 ));
 NAND3xp33_ASAP7_75t_SL \i56/i174  (.A(\i56/n245 ),
    .B(\i56/n188 ),
    .C(\i56/n90 ),
    .Y(\i56/n309 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i56/i175  (.A1(\i56/n65 ),
    .A2(\i56/n69 ),
    .B(\i56/n56 ),
    .C(\i56/n130 ),
    .Y(\i56/n308 ));
 NAND4xp25_ASAP7_75t_SL \i56/i176  (.A(\i56/n547 ),
    .B(\i56/n125 ),
    .C(\i56/n10 ),
    .D(\i56/n12 ),
    .Y(\i56/n307 ));
 OAI211xp5_ASAP7_75t_SL \i56/i177  (.A1(\i56/n58 ),
    .A2(\i56/n519 ),
    .B(\i56/n102 ),
    .C(\i56/n123 ),
    .Y(\i56/n306 ));
 OAI31xp33_ASAP7_75t_SL \i56/i178  (.A1(\i56/n40 ),
    .A2(\i56/n51 ),
    .A3(\i56/n84 ),
    .B(\i56/n73 ),
    .Y(\i56/n305 ));
 AOI221xp5_ASAP7_75t_SL \i56/i179  (.A1(\i56/n169 ),
    .A2(\i56/n59 ),
    .B1(\i56/n53 ),
    .B2(\i56/n89 ),
    .C(\i56/n153 ),
    .Y(\i56/n304 ));
 NOR3xp33_ASAP7_75t_SL \i56/i18  (.A(\i56/n392 ),
    .B(\i56/n455 ),
    .C(\i56/n468 ),
    .Y(\i56/n474 ));
 NOR2xp33_ASAP7_75t_SL \i56/i180  (.A(\i56/n136 ),
    .B(\i56/n510 ),
    .Y(\i56/n303 ));
 OAI221xp5_ASAP7_75t_SL \i56/i181  (.A1(\i56/n41 ),
    .A2(\i56/n39 ),
    .B1(\i56/n52 ),
    .B2(\i56/n68 ),
    .C(\i56/n158 ),
    .Y(\i56/n340 ));
 AOI222xp33_ASAP7_75t_SL \i56/i182  (.A1(\i56/n60 ),
    .A2(\i56/n56 ),
    .B1(\i56/n78 ),
    .B2(\i56/n75 ),
    .C1(\i56/n65 ),
    .C2(\i56/n82 ),
    .Y(\i56/n339 ));
 NAND2xp5_ASAP7_75t_SL \i56/i183  (.A(\i56/n244 ),
    .B(\i56/n206 ),
    .Y(\i56/n337 ));
 OAI221xp5_ASAP7_75t_SL \i56/i184  (.A1(\i56/n519 ),
    .A2(\i56/n55 ),
    .B1(\i56/n483 ),
    .B2(\i56/n57 ),
    .C(\i56/n5 ),
    .Y(\i56/n335 ));
 OAI21xp5_ASAP7_75t_SL \i56/i185  (.A1(\i56/n59 ),
    .A2(\i56/n128 ),
    .B(\i56/n178 ),
    .Y(\i56/n334 ));
 NOR2xp33_ASAP7_75t_SL \i56/i186  (.A(\i56/n131 ),
    .B(\i56/n258 ),
    .Y(\i56/n302 ));
 NAND2xp5_ASAP7_75t_SL \i56/i187  (.A(\i56/n210 ),
    .B(\i56/n243 ),
    .Y(\i56/n332 ));
 NOR2xp33_ASAP7_75t_SL \i56/i188  (.A(\i56/n544 ),
    .B(\i56/n227 ),
    .Y(\i56/n301 ));
 NAND2xp5_ASAP7_75t_SL \i56/i189  (.A(\i56/n213 ),
    .B(\i56/n215 ),
    .Y(\i56/n331 ));
 NOR3xp33_ASAP7_75t_SL \i56/i19  (.A(\i56/n434 ),
    .B(\i56/n421 ),
    .C(\i56/n459 ),
    .Y(\i56/n473 ));
 NAND2xp5_ASAP7_75t_SL \i56/i190  (.A(\i56/n497 ),
    .B(\i56/n250 ),
    .Y(\i56/n330 ));
 OAI221xp5_ASAP7_75t_SL \i56/i191  (.A1(\i56/n548 ),
    .A2(\i56/n536 ),
    .B1(\i56/n70 ),
    .B2(\i56/n86 ),
    .C(\i56/n145 ),
    .Y(\i56/n328 ));
 NAND2x1_ASAP7_75t_SL \i56/i192  (.A(\i56/n541 ),
    .B(\i56/n218 ),
    .Y(\i56/n14 ));
 NAND3xp33_ASAP7_75t_SL \i56/i193  (.A(\i56/n144 ),
    .B(\i56/n139 ),
    .C(\i56/n135 ),
    .Y(\i56/n13 ));
 NOR2xp33_ASAP7_75t_SL \i56/i194  (.A(\i56/n259 ),
    .B(\i56/n252 ),
    .Y(\i56/n300 ));
 OAI211xp5_ASAP7_75t_SL \i56/i195  (.A1(\i56/n81 ),
    .A2(\i56/n72 ),
    .B(\i56/n545 ),
    .C(\i56/n495 ),
    .Y(\i56/n325 ));
 INVxp67_ASAP7_75t_SL \i56/i196  (.A(\i56/n297 ),
    .Y(\i56/n298 ));
 INVxp67_ASAP7_75t_SL \i56/i197  (.A(\i56/n295 ),
    .Y(\i56/n296 ));
 INVxp67_ASAP7_75t_SL \i56/i198  (.A(\i56/n293 ),
    .Y(\i56/n294 ));
 INVx1_ASAP7_75t_SL \i56/i199  (.A(\i56/n291 ),
    .Y(\i56/n292 ));
 AND3x2_ASAP7_75t_SL \i56/i2  (.A(\i56/n469 ),
    .B(\i56/n482 ),
    .C(\i56/n465 ),
    .Y(n8[6]));
 AND4x1_ASAP7_75t_SL \i56/i20  (.A(\i56/n450 ),
    .B(\i56/n456 ),
    .C(\i56/n438 ),
    .D(\i56/n423 ),
    .Y(\i56/n472 ));
 INVx1_ASAP7_75t_SL \i56/i200  (.A(\i56/n289 ),
    .Y(\i56/n290 ));
 OAI22xp5_ASAP7_75t_SL \i56/i201  (.A1(\i56/n483 ),
    .A2(\i56/n492 ),
    .B1(\i56/n76 ),
    .B2(\i56/n72 ),
    .Y(\i56/n287 ));
 AOI21xp5_ASAP7_75t_SL \i56/i202  (.A1(\i56/n107 ),
    .A2(\i56/n77 ),
    .B(\i56/n132 ),
    .Y(\i56/n286 ));
 OAI22xp5_ASAP7_75t_SL \i56/i203  (.A1(\i56/n57 ),
    .A2(\i56/n104 ),
    .B1(\i56/n55 ),
    .B2(\i56/n192 ),
    .Y(\i56/n285 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i56/i204  (.A1(\i56/n71 ),
    .A2(\i56/n67 ),
    .B(\i56/n75 ),
    .C(\i56/n96 ),
    .Y(\i56/n284 ));
 AOI21xp5_ASAP7_75t_SL \i56/i205  (.A1(\i56/n179 ),
    .A2(\i56/n71 ),
    .B(\i56/n237 ),
    .Y(\i56/n283 ));
 AOI22xp5_ASAP7_75t_SL \i56/i206  (.A1(\i56/n51 ),
    .A2(\i56/n108 ),
    .B1(\i56/n80 ),
    .B2(\i56/n172 ),
    .Y(\i56/n282 ));
 AOI211xp5_ASAP7_75t_SL \i56/i207  (.A1(\i56/n51 ),
    .A2(\i56/n54 ),
    .B(\i56/n132 ),
    .C(\i56/n98 ),
    .Y(\i56/n281 ));
 OAI22xp5_ASAP7_75t_SL \i56/i208  (.A1(\i56/n66 ),
    .A2(\i56/n167 ),
    .B1(\i56/n4 ),
    .B2(\i56/n527 ),
    .Y(\i56/n280 ));
 OAI22xp5_ASAP7_75t_SL \i56/i209  (.A1(\i56/n62 ),
    .A2(\i56/n160 ),
    .B1(\i56/n55 ),
    .B2(\i56/n76 ),
    .Y(\i56/n279 ));
 NAND3xp33_ASAP7_75t_SL \i56/i21  (.A(\i56/n408 ),
    .B(\i56/n382 ),
    .C(\i56/n405 ),
    .Y(\i56/n470 ));
 AOI221xp5_ASAP7_75t_SL \i56/i210  (.A1(\i56/n46 ),
    .A2(\i56/n84 ),
    .B1(\i56/n42 ),
    .B2(\i56/n40 ),
    .C(\i56/n238 ),
    .Y(\i56/n278 ));
 AND4x1_ASAP7_75t_SL \i56/i211  (.A(\i56/n138 ),
    .B(\i56/n7 ),
    .C(\i56/n9 ),
    .D(\i56/n145 ),
    .Y(\i56/n277 ));
 NAND4xp25_ASAP7_75t_SL \i56/i212  (.A(\i56/n133 ),
    .B(\i56/n155 ),
    .C(\i56/n121 ),
    .D(\i56/n491 ),
    .Y(\i56/n276 ));
 NAND4xp25_ASAP7_75t_SL \i56/i213  (.A(\i56/n144 ),
    .B(\i56/n141 ),
    .C(\i56/n493 ),
    .D(\i56/n139 ),
    .Y(\i56/n275 ));
 AOI22xp5_ASAP7_75t_SL \i56/i214  (.A1(\i56/n514 ),
    .A2(\i56/n103 ),
    .B1(\i56/n82 ),
    .B2(\i56/n122 ),
    .Y(\i56/n274 ));
 AOI22xp5_ASAP7_75t_SL \i56/i215  (.A1(\i56/n49 ),
    .A2(\i56/n127 ),
    .B1(\i56/n44 ),
    .B2(\i56/n514 ),
    .Y(\i56/n273 ));
 OAI211xp5_ASAP7_75t_SL \i56/i216  (.A1(\i56/n74 ),
    .A2(\i56/n189 ),
    .B(\i56/n93 ),
    .C(\i56/n147 ),
    .Y(\i56/n272 ));
 NAND4xp25_ASAP7_75t_SL \i56/i217  (.A(\i56/n9 ),
    .B(\i56/n161 ),
    .C(\i56/n173 ),
    .D(\i56/n526 ),
    .Y(\i56/n271 ));
 OAI22xp5_ASAP7_75t_SL \i56/i218  (.A1(\i56/n549 ),
    .A2(\i56/n164 ),
    .B1(\i56/n4 ),
    .B2(\i56/n124 ),
    .Y(\i56/n270 ));
 OAI22xp5_ASAP7_75t_SL \i56/i219  (.A1(\i56/n83 ),
    .A2(\i56/n116 ),
    .B1(\i56/n79 ),
    .B2(\i56/n39 ),
    .Y(\i56/n269 ));
 NOR2xp33_ASAP7_75t_SL \i56/i22  (.A(\i56/n442 ),
    .B(\i56/n439 ),
    .Y(\i56/n469 ));
 AOI211x1_ASAP7_75t_SL \i56/i220  (.A1(\i56/n174 ),
    .A2(\i56/n89 ),
    .B(\i56/n546 ),
    .C(\i56/n191 ),
    .Y(\i56/n268 ));
 NAND4xp25_ASAP7_75t_SL \i56/i221  (.A(\i56/n181 ),
    .B(\i56/n530 ),
    .C(\i56/n117 ),
    .D(\i56/n135 ),
    .Y(\i56/n267 ));
 OAI22xp5_ASAP7_75t_SL \i56/i222  (.A1(\i56/n68 ),
    .A2(\i56/n101 ),
    .B1(\i56/n86 ),
    .B2(\i56/n4 ),
    .Y(\i56/n266 ));
 OAI221xp5_ASAP7_75t_R \i56/i223  (.A1(\i56/n119 ),
    .A2(\i56/n501 ),
    .B1(\i56/n76 ),
    .B2(\i56/n88 ),
    .C(\i56/n165 ),
    .Y(\i56/n265 ));
 OAI221xp5_ASAP7_75t_SL \i56/i224  (.A1(\i56/n68 ),
    .A2(\i56/n549 ),
    .B1(\i56/n501 ),
    .B2(\i56/n45 ),
    .C(\i56/n154 ),
    .Y(\i56/n264 ));
 AOI222xp33_ASAP7_75t_SL \i56/i225  (.A1(\i56/n60 ),
    .A2(\i56/n87 ),
    .B1(\i56/n65 ),
    .B2(\i56/n77 ),
    .C1(\i56/n46 ),
    .C2(\i56/n53 ),
    .Y(\i56/n263 ));
 OAI221xp5_ASAP7_75t_SL \i56/i226  (.A1(\i56/n39 ),
    .A2(\i56/n8 ),
    .B1(\i56/n83 ),
    .B2(\i56/n58 ),
    .C(\i56/n112 ),
    .Y(\i56/n262 ));
 OAI211xp5_ASAP7_75t_SL \i56/i227  (.A1(\i56/n58 ),
    .A2(\i56/n146 ),
    .B(\i56/n142 ),
    .C(\i56/n97 ),
    .Y(\i56/n261 ));
 AOI22xp33_ASAP7_75t_SL \i56/i228  (.A1(\i56/n51 ),
    .A2(\i56/n200 ),
    .B1(\i56/n77 ),
    .B2(\i56/n60 ),
    .Y(\i56/n260 ));
 OAI221xp5_ASAP7_75t_SL \i56/i229  (.A1(\i56/n68 ),
    .A2(\i56/n76 ),
    .B1(\i56/n72 ),
    .B2(\i56/n536 ),
    .C(\i56/n528 ),
    .Y(\i56/n299 ));
 NAND2xp5_ASAP7_75t_SL \i56/i23  (.A(\i56/n444 ),
    .B(\i56/n433 ),
    .Y(\i56/n468 ));
 OAI221xp5_ASAP7_75t_SL \i56/i230  (.A1(\i56/n50 ),
    .A2(\i56/n43 ),
    .B1(\i56/n549 ),
    .B2(\i56/n61 ),
    .C(\i56/n106 ),
    .Y(\i56/n297 ));
 AOI221x1_ASAP7_75t_SL \i56/i231  (.A1(\i56/n1 ),
    .A2(\i56/n49 ),
    .B1(\i56/n6 ),
    .B2(\i56/n60 ),
    .C(\i56/n507 ),
    .Y(\i56/n295 ));
 OAI21xp5_ASAP7_75t_L \i56/i232  (.A1(\i56/n192 ),
    .A2(\i56/n61 ),
    .B(\i56/n113 ),
    .Y(\i56/n293 ));
 AOI221x1_ASAP7_75t_SL \i56/i233  (.A1(\i56/n1 ),
    .A2(\i56/n60 ),
    .B1(\i56/n78 ),
    .B2(\i56/n170 ),
    .C(\i56/n162 ),
    .Y(\i56/n291 ));
 OAI221xp5_ASAP7_75t_SL \i56/i234  (.A1(\i56/n163 ),
    .A2(\i56/n519 ),
    .B1(\i56/n86 ),
    .B2(\i56/n45 ),
    .C(\i56/n185 ),
    .Y(\i56/n289 ));
 AOI22xp5_ASAP7_75t_SL \i56/i235  (.A1(\i56/n78 ),
    .A2(\i56/n175 ),
    .B1(\i56/n53 ),
    .B2(\i56/n80 ),
    .Y(\i56/n288 ));
 INVxp67_ASAP7_75t_SL \i56/i236  (.A(\i56/n256 ),
    .Y(\i56/n257 ));
 INVxp67_ASAP7_75t_SL \i56/i237  (.A(\i56/n523 ),
    .Y(\i56/n254 ));
 INVxp67_ASAP7_75t_SL \i56/i238  (.A(\i56/n252 ),
    .Y(\i56/n253 ));
 INVx1_ASAP7_75t_SL \i56/i239  (.A(\i56/n248 ),
    .Y(\i56/n249 ));
 NOR2xp33_ASAP7_75t_SL \i56/i24  (.A(\i56/n422 ),
    .B(\i56/n447 ),
    .Y(\i56/n467 ));
 INVxp67_ASAP7_75t_SL \i56/i240  (.A(\i56/n246 ),
    .Y(\i56/n247 ));
 INVxp67_ASAP7_75t_SL \i56/i241  (.A(\i56/n496 ),
    .Y(\i56/n242 ));
 NOR2xp33_ASAP7_75t_SL \i56/i242  (.A(\i56/n506 ),
    .B(\i56/n179 ),
    .Y(\i56/n241 ));
 OAI21xp5_ASAP7_75t_SL \i56/i243  (.A1(\i56/n47 ),
    .A2(\i56/n44 ),
    .B(\i56/n85 ),
    .Y(\i56/n240 ));
 OAI21xp5_ASAP7_75t_SL \i56/i244  (.A1(\i56/n519 ),
    .A2(\i56/n43 ),
    .B(\i56/n147 ),
    .Y(\i56/n239 ));
 AOI21xp33_ASAP7_75t_SL \i56/i245  (.A1(\i56/n70 ),
    .A2(\i56/n61 ),
    .B(\i56/n176 ),
    .Y(\i56/n238 ));
 OAI21xp5_ASAP7_75t_SL \i56/i246  (.A1(\i56/n83 ),
    .A2(\i56/n66 ),
    .B(\i56/n186 ),
    .Y(\i56/n259 ));
 NAND2xp5_ASAP7_75t_L \i56/i247  (.A(\i56/n490 ),
    .B(\i56/n156 ),
    .Y(\i56/n237 ));
 OAI21xp33_ASAP7_75t_SL \i56/i248  (.A1(\i56/n63 ),
    .A2(\i56/n66 ),
    .B(\i56/n493 ),
    .Y(\i56/n236 ));
 AOI21xp5_ASAP7_75t_SL \i56/i249  (.A1(\i56/n41 ),
    .A2(\i56/n79 ),
    .B(\i56/n549 ),
    .Y(\i56/n258 ));
 NOR2xp33_ASAP7_75t_SL \i56/i25  (.A(\i56/n455 ),
    .B(\i56/n449 ),
    .Y(\i56/n466 ));
 AOI21xp33_ASAP7_75t_SL \i56/i250  (.A1(\i56/n79 ),
    .A2(\i56/n48 ),
    .B(\i56/n176 ),
    .Y(\i56/n235 ));
 OAI21xp5_ASAP7_75t_SL \i56/i251  (.A1(\i56/n62 ),
    .A2(\i56/n66 ),
    .B(\i56/n140 ),
    .Y(\i56/n234 ));
 NOR2xp33_ASAP7_75t_SL \i56/i252  (.A(\i56/n152 ),
    .B(\i56/n182 ),
    .Y(\i56/n233 ));
 OAI22xp5_ASAP7_75t_SL \i56/i253  (.A1(\i56/n536 ),
    .A2(\i56/n61 ),
    .B1(\i56/n81 ),
    .B2(\i56/n41 ),
    .Y(\i56/n232 ));
 OAI21xp5_ASAP7_75t_SL \i56/i254  (.A1(\i56/n55 ),
    .A2(\i56/n52 ),
    .B(\i56/n196 ),
    .Y(\i56/n231 ));
 OAI21xp33_ASAP7_75t_SL \i56/i255  (.A1(\i56/n55 ),
    .A2(\i56/n62 ),
    .B(\i56/n7 ),
    .Y(\i56/n256 ));
 OAI21xp5_ASAP7_75t_SL \i56/i256  (.A1(\i56/n86 ),
    .A2(\i56/n68 ),
    .B(\i56/n199 ),
    .Y(\i56/n255 ));
 OAI22xp5_ASAP7_75t_SL \i56/i257  (.A1(\i56/n70 ),
    .A2(\i56/n63 ),
    .B1(\i56/n501 ),
    .B2(\i56/n68 ),
    .Y(\i56/n252 ));
 AO22x2_ASAP7_75t_SL \i56/i258  (.A1(\i56/n514 ),
    .A2(\i56/n60 ),
    .B1(\i56/n51 ),
    .B2(\i56/n65 ),
    .Y(\i56/n251 ));
 AOI22xp5_ASAP7_75t_SL \i56/i259  (.A1(\i56/n78 ),
    .A2(\i56/n64 ),
    .B1(\i56/n77 ),
    .B2(\i56/n80 ),
    .Y(\i56/n250 ));
 AND2x2_ASAP7_75t_SL \i56/i26  (.A(\i56/n413 ),
    .B(\i56/n446 ),
    .Y(\i56/n471 ));
 OAI22xp5_ASAP7_75t_SL \i56/i260  (.A1(\i56/n57 ),
    .A2(\i56/n61 ),
    .B1(\i56/n74 ),
    .B2(\i56/n4 ),
    .Y(\i56/n230 ));
 OAI21xp5_ASAP7_75t_SL \i56/i261  (.A1(\i56/n55 ),
    .A2(\i56/n39 ),
    .B(\i56/n10 ),
    .Y(\i56/n248 ));
 NAND2xp5_ASAP7_75t_SL \i56/i262  (.A(\i56/n44 ),
    .B(\i56/n6 ),
    .Y(\i56/n246 ));
 OAI21xp5_ASAP7_75t_SL \i56/i263  (.A1(\i56/n78 ),
    .A2(\i56/n69 ),
    .B(\i56/n1 ),
    .Y(\i56/n245 ));
 NAND2xp5_ASAP7_75t_SL \i56/i264  (.A(\i56/n89 ),
    .B(\i56/n175 ),
    .Y(\i56/n244 ));
 AOI22xp5_ASAP7_75t_SL \i56/i265  (.A1(\i56/n54 ),
    .A2(\i56/n84 ),
    .B1(\i56/n56 ),
    .B2(\i56/n71 ),
    .Y(\i56/n243 ));
 INVxp67_ASAP7_75t_SL \i56/i266  (.A(\i56/n228 ),
    .Y(\i56/n229 ));
 INVxp67_ASAP7_75t_SL \i56/i267  (.A(\i56/n508 ),
    .Y(\i56/n222 ));
 INVxp67_ASAP7_75t_SL \i56/i268  (.A(\i56/n542 ),
    .Y(\i56/n221 ));
 INVx1_ASAP7_75t_SL \i56/i269  (.A(\i56/n543 ),
    .Y(\i56/n217 ));
 NOR2xp33_ASAP7_75t_SL \i56/i27  (.A(\i56/n454 ),
    .B(\i56/n436 ),
    .Y(\i56/n464 ));
 AOI22xp33_ASAP7_75t_SL \i56/i270  (.A1(\i56/n40 ),
    .A2(\i56/n60 ),
    .B1(\i56/n54 ),
    .B2(\i56/n56 ),
    .Y(\i56/n214 ));
 OAI21xp5_ASAP7_75t_SL \i56/i271  (.A1(\i56/n44 ),
    .A2(\i56/n42 ),
    .B(\i56/n53 ),
    .Y(\i56/n213 ));
 AOI21xp33_ASAP7_75t_SL \i56/i272  (.A1(\i56/n66 ),
    .A2(\i56/n79 ),
    .B(\i56/n39 ),
    .Y(\i56/n212 ));
 AOI22xp5_ASAP7_75t_SL \i56/i273  (.A1(\i56/n89 ),
    .A2(\i56/n84 ),
    .B1(\i56/n51 ),
    .B2(\i56/n73 ),
    .Y(\i56/n211 ));
 AOI22xp5_ASAP7_75t_SL \i56/i274  (.A1(\i56/n59 ),
    .A2(\i56/n64 ),
    .B1(\i56/n80 ),
    .B2(\i56/n514 ),
    .Y(\i56/n210 ));
 AOI22xp5_ASAP7_75t_SL \i56/i275  (.A1(\i56/n89 ),
    .A2(\i56/n64 ),
    .B1(\i56/n87 ),
    .B2(\i56/n44 ),
    .Y(\i56/n228 ));
 OAI22xp5_ASAP7_75t_SL \i56/i276  (.A1(\i56/n39 ),
    .A2(\i56/n66 ),
    .B1(\i56/n483 ),
    .B2(\i56/n63 ),
    .Y(\i56/n209 ));
 OAI22xp5_ASAP7_75t_R \i56/i277  (.A1(\i56/n501 ),
    .A2(\i56/n58 ),
    .B1(\i56/n55 ),
    .B2(\i56/n549 ),
    .Y(\i56/n208 ));
 OAI21xp5_ASAP7_75t_SL \i56/i278  (.A1(\i56/n536 ),
    .A2(\i56/n41 ),
    .B(\i56/n126 ),
    .Y(\i56/n207 ));
 AOI22xp5_ASAP7_75t_SL \i56/i279  (.A1(\i56/n514 ),
    .A2(\i56/n71 ),
    .B1(\i56/n40 ),
    .B2(\i56/n47 ),
    .Y(\i56/n206 ));
 NOR2xp33_ASAP7_75t_SL \i56/i28  (.A(\i56/n435 ),
    .B(\i56/n430 ),
    .Y(\i56/n463 ));
 OAI22xp5_ASAP7_75t_SL \i56/i280  (.A1(\i56/n88 ),
    .A2(\i56/n536 ),
    .B1(\i56/n43 ),
    .B2(\i56/n63 ),
    .Y(\i56/n227 ));
 OAI22xp5_ASAP7_75t_SL \i56/i281  (.A1(\i56/n76 ),
    .A2(\i56/n66 ),
    .B1(\i56/n39 ),
    .B2(\i56/n70 ),
    .Y(\i56/n226 ));
 NAND2xp5_ASAP7_75t_SL \i56/i282  (.A(\i56/n545 ),
    .B(\i56/n495 ),
    .Y(\i56/n205 ));
 AOI22xp5_ASAP7_75t_SL \i56/i283  (.A1(\i56/n51 ),
    .A2(\i56/n67 ),
    .B1(\i56/n47 ),
    .B2(\i56/n1 ),
    .Y(\i56/n225 ));
 NAND2xp5_ASAP7_75t_SL \i56/i284  (.A(\i56/n201 ),
    .B(\i56/n151 ),
    .Y(\i56/n204 ));
 OAI22xp5_ASAP7_75t_SL \i56/i285  (.A1(\i56/n55 ),
    .A2(\i56/n536 ),
    .B1(\i56/n74 ),
    .B2(\i56/n72 ),
    .Y(\i56/n224 ));
 OAI22xp33_ASAP7_75t_SL \i56/i286  (.A1(\i56/n549 ),
    .A2(\i56/n48 ),
    .B1(\i56/n483 ),
    .B2(\i56/n74 ),
    .Y(\i56/n203 ));
 OAI22xp5_ASAP7_75t_SL \i56/i287  (.A1(\i56/n66 ),
    .A2(\i56/n74 ),
    .B1(\i56/n43 ),
    .B2(\i56/n39 ),
    .Y(\i56/n223 ));
 OAI22xp5_ASAP7_75t_SL \i56/i288  (.A1(\i56/n501 ),
    .A2(\i56/n41 ),
    .B1(\i56/n72 ),
    .B2(\i56/n57 ),
    .Y(\i56/n220 ));
 OAI22xp5_ASAP7_75t_SL \i56/i289  (.A1(\i56/n48 ),
    .A2(\i56/n50 ),
    .B1(\i56/n4 ),
    .B2(\i56/n39 ),
    .Y(\i56/n219 ));
 NOR2xp33_ASAP7_75t_SL \i56/i29  (.A(\i56/n429 ),
    .B(\i56/n448 ),
    .Y(\i56/n462 ));
 AOI22xp5_ASAP7_75t_SL \i56/i290  (.A1(\i56/n64 ),
    .A2(\i56/n60 ),
    .B1(\i56/n40 ),
    .B2(\i56/n69 ),
    .Y(\i56/n218 ));
 AOI22xp5_ASAP7_75t_SL \i56/i291  (.A1(\i56/n49 ),
    .A2(\i56/n40 ),
    .B1(\i56/n56 ),
    .B2(\i56/n47 ),
    .Y(\i56/n202 ));
 AOI22xp5_ASAP7_75t_SL \i56/i292  (.A1(\i56/n42 ),
    .A2(\i56/n64 ),
    .B1(\i56/n82 ),
    .B2(\i56/n80 ),
    .Y(\i56/n216 ));
 AOI22xp5_ASAP7_75t_SL \i56/i293  (.A1(\i56/n71 ),
    .A2(\i56/n85 ),
    .B1(\i56/n75 ),
    .B2(\i56/n59 ),
    .Y(\i56/n215 ));
 INVxp67_ASAP7_75t_SL \i56/i294  (.A(\i56/n197 ),
    .Y(\i56/n198 ));
 INVxp67_ASAP7_75t_SL \i56/i295  (.A(\i56/n530 ),
    .Y(\i56/n195 ));
 INVxp67_ASAP7_75t_SL \i56/i296  (.A(\i56/n506 ),
    .Y(\i56/n194 ));
 INVxp67_ASAP7_75t_SL \i56/i297  (.A(\i56/n546 ),
    .Y(\i56/n193 ));
 INVxp67_ASAP7_75t_SL \i56/i298  (.A(\i56/n547 ),
    .Y(\i56/n187 ));
 INVx1_ASAP7_75t_SL \i56/i299  (.A(\i56/n183 ),
    .Y(\i56/n184 ));
 AND2x4_ASAP7_75t_SL \i56/i3  (.A(\i56/n480 ),
    .B(\i56/n472 ),
    .Y(n8[3]));
 AND4x1_ASAP7_75t_SL \i56/i30  (.A(\i56/n418 ),
    .B(\i56/n414 ),
    .C(\i56/n374 ),
    .D(\i56/n367 ),
    .Y(\i56/n461 ));
 INVxp67_ASAP7_75t_SL \i56/i300  (.A(\i56/n181 ),
    .Y(\i56/n182 ));
 INVxp67_ASAP7_75t_SL \i56/i301  (.A(\i56/n179 ),
    .Y(\i56/n180 ));
 INVx1_ASAP7_75t_SL \i56/i302  (.A(\i56/n177 ),
    .Y(\i56/n178 ));
 NAND2xp5_ASAP7_75t_L \i56/i303  (.A(\i56/n86 ),
    .B(\i56/n76 ),
    .Y(\i56/n174 ));
 NAND2xp5_ASAP7_75t_SL \i56/i304  (.A(\i56/n84 ),
    .B(\i56/n42 ),
    .Y(\i56/n173 ));
 NAND2xp33_ASAP7_75t_L \i56/i305  (.A(\i56/n536 ),
    .B(\i56/n81 ),
    .Y(\i56/n172 ));
 NOR2xp33_ASAP7_75t_L \i56/i306  (.A(\i56/n47 ),
    .B(\i56/n65 ),
    .Y(\i56/n171 ));
 NAND2xp5_ASAP7_75t_SL \i56/i307  (.A(\i56/n52 ),
    .B(\i56/n83 ),
    .Y(\i56/n170 ));
 NAND2xp5_ASAP7_75t_SL \i56/i308  (.A(\i56/n63 ),
    .B(\i56/n83 ),
    .Y(\i56/n169 ));
 NAND2xp5_ASAP7_75t_SL \i56/i309  (.A(\i56/n73 ),
    .B(\i56/n84 ),
    .Y(\i56/n168 ));
 NOR3xp33_ASAP7_75t_SL \i56/i31  (.A(\i56/n399 ),
    .B(\i56/n343 ),
    .C(\i56/n411 ),
    .Y(\i56/n460 ));
 NOR2xp33_ASAP7_75t_SL \i56/i310  (.A(\i56/n82 ),
    .B(\i56/n85 ),
    .Y(\i56/n167 ));
 NAND2xp5_ASAP7_75t_SL \i56/i311  (.A(\i56/n59 ),
    .B(\i56/n514 ),
    .Y(\i56/n166 ));
 NAND2xp5_ASAP7_75t_SL \i56/i312  (.A(\i56/n65 ),
    .B(\i56/n53 ),
    .Y(\i56/n165 ));
 NOR2xp33_ASAP7_75t_SL \i56/i313  (.A(\i56/n54 ),
    .B(\i56/n42 ),
    .Y(\i56/n164 ));
 NOR2xp33_ASAP7_75t_SL \i56/i314  (.A(\i56/n67 ),
    .B(\i56/n47 ),
    .Y(\i56/n163 ));
 NOR2xp67_ASAP7_75t_SL \i56/i315  (.A(\i56/n501 ),
    .B(\i56/n72 ),
    .Y(\i56/n162 ));
 NAND2xp5_ASAP7_75t_SL \i56/i316  (.A(\i56/n85 ),
    .B(\i56/n46 ),
    .Y(\i56/n161 ));
 NOR2xp33_ASAP7_75t_SL \i56/i317  (.A(\i56/n67 ),
    .B(\i56/n73 ),
    .Y(\i56/n160 ));
 NOR2xp33_ASAP7_75t_SL \i56/i318  (.A(\i56/n44 ),
    .B(\i56/n67 ),
    .Y(\i56/n159 ));
 NAND2xp5_ASAP7_75t_SL \i56/i319  (.A(\i56/n49 ),
    .B(\i56/n75 ),
    .Y(\i56/n158 ));
 NAND2xp33_ASAP7_75t_SL \i56/i32  (.A(\i56/n15 ),
    .B(\i56/n431 ),
    .Y(\i56/n459 ));
 NOR2xp33_ASAP7_75t_SL \i56/i320  (.A(\i56/n78 ),
    .B(\i56/n73 ),
    .Y(\i56/n157 ));
 NAND2xp5_ASAP7_75t_SL \i56/i321  (.A(\i56/n75 ),
    .B(\i56/n47 ),
    .Y(\i56/n201 ));
 NAND2xp5_ASAP7_75t_SL \i56/i322  (.A(\i56/n80 ),
    .B(\i56/n64 ),
    .Y(\i56/n156 ));
 NAND2xp5_ASAP7_75t_SL \i56/i323  (.A(\i56/n75 ),
    .B(\i56/n69 ),
    .Y(\i56/n155 ));
 NAND2xp5_ASAP7_75t_SL \i56/i324  (.A(\i56/n54 ),
    .B(\i56/n75 ),
    .Y(\i56/n154 ));
 NAND2xp5_ASAP7_75t_SL \i56/i325  (.A(\i56/n65 ),
    .B(\i56/n84 ),
    .Y(\i56/n12 ));
 NAND2xp5_ASAP7_75t_SL \i56/i326  (.A(\i56/n1 ),
    .B(\i56/n71 ),
    .Y(\i56/n11 ));
 NAND2xp33_ASAP7_75t_SL \i56/i327  (.A(\i56/n43 ),
    .B(\i56/n79 ),
    .Y(\i56/n200 ));
 NAND2xp5_ASAP7_75t_SL \i56/i328  (.A(\i56/n56 ),
    .B(\i56/n67 ),
    .Y(\i56/n10 ));
 NAND2xp5_ASAP7_75t_SL \i56/i329  (.A(\i56/n80 ),
    .B(\i56/n1 ),
    .Y(\i56/n9 ));
 AND3x1_ASAP7_75t_SL \i56/i33  (.A(\i56/n417 ),
    .B(\i56/n2 ),
    .C(\i56/n410 ),
    .Y(\i56/n465 ));
 NOR2xp33_ASAP7_75t_SL \i56/i330  (.A(\i56/n79 ),
    .B(\i56/n76 ),
    .Y(\i56/n153 ));
 NAND2xp5_ASAP7_75t_SL \i56/i331  (.A(\i56/n89 ),
    .B(\i56/n56 ),
    .Y(\i56/n199 ));
 NAND2xp5_ASAP7_75t_L \i56/i332  (.A(\i56/n85 ),
    .B(\i56/n89 ),
    .Y(\i56/n197 ));
 NAND2xp5_ASAP7_75t_SL \i56/i333  (.A(\i56/n82 ),
    .B(\i56/n78 ),
    .Y(\i56/n196 ));
 NOR2x1_ASAP7_75t_SL \i56/i334  (.A(\i56/n75 ),
    .B(\i56/n53 ),
    .Y(\i56/n192 ));
 AND2x2_ASAP7_75t_SL \i56/i335  (.A(\i56/n514 ),
    .B(\i56/n73 ),
    .Y(\i56/n191 ));
 NAND2xp5_ASAP7_75t_SL \i56/i336  (.A(\i56/n75 ),
    .B(\i56/n46 ),
    .Y(\i56/n190 ));
 NOR2xp33_ASAP7_75t_L \i56/i337  (.A(\i56/n44 ),
    .B(\i56/n65 ),
    .Y(\i56/n189 ));
 NAND2xp5_ASAP7_75t_SL \i56/i338  (.A(\i56/n80 ),
    .B(\i56/n84 ),
    .Y(\i56/n188 ));
 NAND2xp5_ASAP7_75t_SL \i56/i339  (.A(\i56/n65 ),
    .B(\i56/n40 ),
    .Y(\i56/n186 ));
 INVxp67_ASAP7_75t_SL \i56/i34  (.A(\i56/n457 ),
    .Y(\i56/n458 ));
 NAND2xp5_ASAP7_75t_SL \i56/i340  (.A(\i56/n65 ),
    .B(\i56/n85 ),
    .Y(\i56/n185 ));
 NOR2xp33_ASAP7_75t_SL \i56/i341  (.A(\i56/n50 ),
    .B(\i56/n483 ),
    .Y(\i56/n152 ));
 NOR2xp33_ASAP7_75t_L \i56/i342  (.A(\i56/n40 ),
    .B(\i56/n75 ),
    .Y(\i56/n183 ));
 NAND2xp5_ASAP7_75t_SL \i56/i343  (.A(\i56/n89 ),
    .B(\i56/n1 ),
    .Y(\i56/n181 ));
 NAND2xp5_ASAP7_75t_L \i56/i344  (.A(\i56/n83 ),
    .B(\i56/n81 ),
    .Y(\i56/n179 ));
 NOR2xp33_ASAP7_75t_L \i56/i345  (.A(\i56/n87 ),
    .B(\i56/n82 ),
    .Y(\i56/n177 ));
 NOR2xp33_ASAP7_75t_L \i56/i346  (.A(\i56/n87 ),
    .B(\i56/n75 ),
    .Y(\i56/n176 ));
 NAND2xp5_ASAP7_75t_SL \i56/i347  (.A(\i56/n50 ),
    .B(\i56/n519 ),
    .Y(\i56/n175 ));
 INVxp67_ASAP7_75t_SL \i56/i348  (.A(\i56/n490 ),
    .Y(\i56/n148 ));
 INVxp67_ASAP7_75t_SL \i56/i349  (.A(\i56/n142 ),
    .Y(\i56/n143 ));
 INVxp67_ASAP7_75t_SL \i56/i35  (.A(\i56/n455 ),
    .Y(\i56/n456 ));
 INVxp67_ASAP7_75t_SL \i56/i350  (.A(\i56/n136 ),
    .Y(\i56/n137 ));
 INVxp67_ASAP7_75t_SL \i56/i351  (.A(\i56/n133 ),
    .Y(\i56/n134 ));
 INVxp67_ASAP7_75t_SL \i56/i352  (.A(\i56/n5 ),
    .Y(\i56/n130 ));
 NOR2xp33_ASAP7_75t_SL \i56/i353  (.A(\i56/n44 ),
    .B(\i56/n59 ),
    .Y(\i56/n129 ));
 NOR2xp33_ASAP7_75t_SL \i56/i354  (.A(\i56/n86 ),
    .B(\i56/n548 ),
    .Y(\i56/n128 ));
 NAND2xp33_ASAP7_75t_SL \i56/i355  (.A(\i56/n57 ),
    .B(\i56/n81 ),
    .Y(\i56/n127 ));
 NAND2xp5_ASAP7_75t_SL \i56/i356  (.A(\i56/n44 ),
    .B(\i56/n85 ),
    .Y(\i56/n126 ));
 NAND2xp5_ASAP7_75t_SL \i56/i357  (.A(\i56/n87 ),
    .B(\i56/n42 ),
    .Y(\i56/n125 ));
 NOR2xp33_ASAP7_75t_SL \i56/i358  (.A(\i56/n87 ),
    .B(\i56/n53 ),
    .Y(\i56/n124 ));
 NAND2xp5_ASAP7_75t_SL \i56/i359  (.A(\i56/n49 ),
    .B(\i56/n40 ),
    .Y(\i56/n123 ));
 NAND3xp33_ASAP7_75t_SL \i56/i36  (.A(\i56/n407 ),
    .B(\i56/n358 ),
    .C(\i56/n366 ),
    .Y(\i56/n453 ));
 NAND2xp33_ASAP7_75t_L \i56/i360  (.A(\i56/n61 ),
    .B(\i56/n58 ),
    .Y(\i56/n122 ));
 NAND2xp5_ASAP7_75t_SL \i56/i361  (.A(\i56/n77 ),
    .B(\i56/n78 ),
    .Y(\i56/n121 ));
 NAND2xp33_ASAP7_75t_SL \i56/i362  (.A(\i56/n62 ),
    .B(\i56/n57 ),
    .Y(\i56/n120 ));
 NOR2xp33_ASAP7_75t_SL \i56/i363  (.A(\i56/n49 ),
    .B(\i56/n46 ),
    .Y(\i56/n119 ));
 NOR2xp33_ASAP7_75t_SL \i56/i364  (.A(\i56/n1 ),
    .B(\i56/n40 ),
    .Y(\i56/n118 ));
 NAND2xp5_ASAP7_75t_SL \i56/i365  (.A(\i56/n77 ),
    .B(\i56/n49 ),
    .Y(\i56/n117 ));
 NOR2xp33_ASAP7_75t_L \i56/i366  (.A(\i56/n49 ),
    .B(\i56/n69 ),
    .Y(\i56/n116 ));
 NAND2xp5_ASAP7_75t_SL \i56/i367  (.A(\i56/n49 ),
    .B(\i56/n53 ),
    .Y(\i56/n115 ));
 NAND2xp5_ASAP7_75t_SL \i56/i368  (.A(\i56/n78 ),
    .B(\i56/n56 ),
    .Y(\i56/n114 ));
 NAND2xp5_ASAP7_75t_SL \i56/i369  (.A(\i56/n1 ),
    .B(\i56/n59 ),
    .Y(\i56/n113 ));
 NAND3xp33_ASAP7_75t_SL \i56/i37  (.A(\i56/n359 ),
    .B(\i56/n345 ),
    .C(\i56/n322 ),
    .Y(\i56/n452 ));
 NAND2xp5_ASAP7_75t_SL \i56/i370  (.A(\i56/n49 ),
    .B(\i56/n82 ),
    .Y(\i56/n112 ));
 NAND2xp33_ASAP7_75t_SL \i56/i371  (.A(\i56/n43 ),
    .B(\i56/n70 ),
    .Y(\i56/n111 ));
 NAND2xp33_ASAP7_75t_SL \i56/i372  (.A(\i56/n76 ),
    .B(\i56/n72 ),
    .Y(\i56/n110 ));
 NOR2xp33_ASAP7_75t_SL \i56/i373  (.A(\i56/n46 ),
    .B(\i56/n71 ),
    .Y(\i56/n109 ));
 NAND2xp33_ASAP7_75t_L \i56/i374  (.A(\i56/n45 ),
    .B(\i56/n55 ),
    .Y(\i56/n108 ));
 NAND2xp5_ASAP7_75t_SL \i56/i375  (.A(\i56/n46 ),
    .B(\i56/n64 ),
    .Y(\i56/n151 ));
 NAND2xp33_ASAP7_75t_SL \i56/i376  (.A(\i56/n548 ),
    .B(\i56/n45 ),
    .Y(\i56/n107 ));
 NAND2xp5_ASAP7_75t_SL \i56/i377  (.A(\i56/n53 ),
    .B(\i56/n73 ),
    .Y(\i56/n106 ));
 NAND2xp5_ASAP7_75t_SL \i56/i378  (.A(\i56/n46 ),
    .B(\i56/n51 ),
    .Y(\i56/n150 ));
 NOR2xp33_ASAP7_75t_SL \i56/i379  (.A(\i56/n50 ),
    .B(\i56/n70 ),
    .Y(\i56/n105 ));
 NAND2xp5_ASAP7_75t_L \i56/i38  (.A(\i56/n553 ),
    .B(\i56/n386 ),
    .Y(\i56/n451 ));
 NOR2xp33_ASAP7_75t_SL \i56/i380  (.A(\i56/n59 ),
    .B(\i56/n42 ),
    .Y(\i56/n104 ));
 NAND2xp5_ASAP7_75t_R \i56/i381  (.A(\i56/n548 ),
    .B(\i56/n68 ),
    .Y(\i56/n103 ));
 NAND2xp5_ASAP7_75t_SL \i56/i382  (.A(\i56/n56 ),
    .B(\i56/n47 ),
    .Y(\i56/n102 ));
 NOR2xp33_ASAP7_75t_SL \i56/i383  (.A(\i56/n56 ),
    .B(\i56/n40 ),
    .Y(\i56/n101 ));
 NAND2xp5_ASAP7_75t_L \i56/i384  (.A(\i56/n57 ),
    .B(\i56/n76 ),
    .Y(\i56/n100 ));
 NAND2xp5_ASAP7_75t_SL \i56/i385  (.A(\i56/n82 ),
    .B(\i56/n69 ),
    .Y(\i56/n99 ));
 NOR2xp33_ASAP7_75t_SL \i56/i386  (.A(\i56/n78 ),
    .B(\i56/n71 ),
    .Y(\i56/n8 ));
 NAND2xp5_ASAP7_75t_SL \i56/i387  (.A(\i56/n53 ),
    .B(\i56/n71 ),
    .Y(\i56/n149 ));
 NOR2xp33_ASAP7_75t_SL \i56/i388  (.A(\i56/n57 ),
    .B(\i56/n70 ),
    .Y(\i56/n98 ));
 NAND2xp5_ASAP7_75t_SL \i56/i389  (.A(\i56/n51 ),
    .B(\i56/n60 ),
    .Y(\i56/n97 ));
 NOR2xp33_ASAP7_75t_SL \i56/i39  (.A(\i56/n415 ),
    .B(\i56/n341 ),
    .Y(\i56/n450 ));
 NOR2xp33_ASAP7_75t_SL \i56/i390  (.A(\i56/n81 ),
    .B(\i56/n41 ),
    .Y(\i56/n96 ));
 NOR2xp33_ASAP7_75t_SL \i56/i391  (.A(\i56/n501 ),
    .B(\i56/n68 ),
    .Y(\i56/n95 ));
 NAND2xp5_ASAP7_75t_SL \i56/i392  (.A(\i56/n54 ),
    .B(\i56/n82 ),
    .Y(\i56/n147 ));
 NAND2xp5_ASAP7_75t_SL \i56/i393  (.A(\i56/n64 ),
    .B(\i56/n73 ),
    .Y(\i56/n7 ));
 NAND2x1p5_ASAP7_75t_SL \i56/i394  (.A(\i56/n81 ),
    .B(\i56/n76 ),
    .Y(\i56/n6 ));
 NOR2xp33_ASAP7_75t_L \i56/i395  (.A(\i56/n1 ),
    .B(\i56/n77 ),
    .Y(\i56/n146 ));
 NAND2xp5_ASAP7_75t_SL \i56/i396  (.A(\i56/n77 ),
    .B(\i56/n42 ),
    .Y(\i56/n145 ));
 NAND2xp5_ASAP7_75t_SL \i56/i397  (.A(\i56/n56 ),
    .B(\i56/n42 ),
    .Y(\i56/n144 ));
 NOR2xp33_ASAP7_75t_SL \i56/i398  (.A(\i56/n55 ),
    .B(\i56/n63 ),
    .Y(\i56/n94 ));
 NAND2xp5_ASAP7_75t_SL \i56/i399  (.A(\i56/n54 ),
    .B(\i56/n87 ),
    .Y(\i56/n93 ));
 AND3x4_ASAP7_75t_SL \i56/i4  (.A(\i56/n465 ),
    .B(\i56/n474 ),
    .C(\i56/n471 ),
    .Y(n8[4]));
 NAND2xp33_ASAP7_75t_L \i56/i40  (.A(\i56/n391 ),
    .B(\i56/n409 ),
    .Y(\i56/n449 ));
 NAND2xp5_ASAP7_75t_SL \i56/i400  (.A(\i56/n40 ),
    .B(\i56/n60 ),
    .Y(\i56/n92 ));
 NAND2xp5_ASAP7_75t_SL \i56/i401  (.A(\i56/n51 ),
    .B(\i56/n47 ),
    .Y(\i56/n142 ));
 NAND2xp5_ASAP7_75t_SL \i56/i402  (.A(\i56/n51 ),
    .B(\i56/n69 ),
    .Y(\i56/n141 ));
 NAND2xp5_ASAP7_75t_SL \i56/i403  (.A(\i56/n64 ),
    .B(\i56/n47 ),
    .Y(\i56/n140 ));
 NOR2xp33_ASAP7_75t_SL \i56/i404  (.A(\i56/n548 ),
    .B(\i56/n52 ),
    .Y(\i56/n91 ));
 NAND2xp5_ASAP7_75t_SL \i56/i405  (.A(\i56/n40 ),
    .B(\i56/n59 ),
    .Y(\i56/n139 ));
 NAND2xp5_ASAP7_75t_SL \i56/i406  (.A(\i56/n53 ),
    .B(\i56/n59 ),
    .Y(\i56/n138 ));
 AND2x2_ASAP7_75t_SL \i56/i407  (.A(\i56/n56 ),
    .B(\i56/n44 ),
    .Y(\i56/n136 ));
 NAND4xp25_ASAP7_75t_SL \i56/i408  (.A(\i56/n33 ),
    .B(\i56/n37 ),
    .C(\i56/n533 ),
    .D(\i56/n25 ),
    .Y(\i56/n135 ));
 NAND2xp5_ASAP7_75t_SL \i56/i409  (.A(\i56/n46 ),
    .B(\i56/n40 ),
    .Y(\i56/n133 ));
 NAND3xp33_ASAP7_75t_SL \i56/i41  (.A(\i56/n420 ),
    .B(\i56/n540 ),
    .C(\i56/n288 ),
    .Y(\i56/n448 ));
 NAND2xp5_ASAP7_75t_SL \i56/i410  (.A(\i56/n49 ),
    .B(\i56/n64 ),
    .Y(\i56/n90 ));
 AND2x2_ASAP7_75t_SL \i56/i411  (.A(\i56/n53 ),
    .B(\i56/n44 ),
    .Y(\i56/n132 ));
 AND2x2_ASAP7_75t_SL \i56/i412  (.A(\i56/n51 ),
    .B(\i56/n59 ),
    .Y(\i56/n131 ));
 NAND2xp5_ASAP7_75t_SL \i56/i413  (.A(\i56/n85 ),
    .B(\i56/n59 ),
    .Y(\i56/n5 ));
 INVx2_ASAP7_75t_SL \i56/i414  (.A(\i56/n89 ),
    .Y(\i56/n88 ));
 INVx4_ASAP7_75t_SL \i56/i415  (.A(\i56/n87 ),
    .Y(\i56/n86 ));
 INVx3_ASAP7_75t_SL \i56/i416  (.A(\i56/n82 ),
    .Y(\i56/n81 ));
 INVx2_ASAP7_75t_SL \i56/i417  (.A(\i56/n80 ),
    .Y(\i56/n79 ));
 INVx3_ASAP7_75t_SL \i56/i418  (.A(\i56/n77 ),
    .Y(\i56/n76 ));
 INVx2_ASAP7_75t_SL \i56/i419  (.A(\i56/n75 ),
    .Y(\i56/n74 ));
 NAND2xp33_ASAP7_75t_SL \i56/i42  (.A(\i56/n402 ),
    .B(\i56/n406 ),
    .Y(\i56/n447 ));
 INVx2_ASAP7_75t_SL \i56/i420  (.A(\i56/n73 ),
    .Y(\i56/n72 ));
 INVx2_ASAP7_75t_SL \i56/i421  (.A(\i56/n71 ),
    .Y(\i56/n70 ));
 INVx3_ASAP7_75t_SL \i56/i422  (.A(\i56/n69 ),
    .Y(\i56/n68 ));
 INVx3_ASAP7_75t_SL \i56/i423  (.A(\i56/n67 ),
    .Y(\i56/n66 ));
 AND2x4_ASAP7_75t_SL \i56/i424  (.A(\i56/n29 ),
    .B(\i56/n31 ),
    .Y(\i56/n89 ));
 AND2x4_ASAP7_75t_SL \i56/i425  (.A(\i56/n488 ),
    .B(\i56/n38 ),
    .Y(\i56/n87 ));
 AND2x4_ASAP7_75t_SL \i56/i426  (.A(\i56/n517 ),
    .B(\i56/n25 ),
    .Y(\i56/n85 ));
 AND2x4_ASAP7_75t_SL \i56/i427  (.A(\i56/n516 ),
    .B(\i56/n533 ),
    .Y(\i56/n84 ));
 AND2x4_ASAP7_75t_SL \i56/i428  (.A(\i56/n34 ),
    .B(\i56/n25 ),
    .Y(\i56/n82 ));
 AND2x4_ASAP7_75t_SL \i56/i429  (.A(\i56/n36 ),
    .B(\i56/n35 ),
    .Y(\i56/n80 ));
 NOR2xp33_ASAP7_75t_SL \i56/i43  (.A(\i56/n404 ),
    .B(\i56/n403 ),
    .Y(\i56/n446 ));
 AND2x2_ASAP7_75t_SL \i56/i430  (.A(\i56/n36 ),
    .B(\i56/n27 ),
    .Y(\i56/n78 ));
 NAND2x1_ASAP7_75t_SL \i56/i431  (.A(\i56/n36 ),
    .B(\i56/n27 ),
    .Y(\i56/n4 ));
 AND2x4_ASAP7_75t_SL \i56/i432  (.A(\i56/n488 ),
    .B(\i56/n516 ),
    .Y(\i56/n77 ));
 AND2x4_ASAP7_75t_SL \i56/i433  (.A(\i56/n488 ),
    .B(\i56/n25 ),
    .Y(\i56/n75 ));
 AND2x4_ASAP7_75t_SL \i56/i434  (.A(\i56/n36 ),
    .B(\i56/n26 ),
    .Y(\i56/n73 ));
 AND2x4_ASAP7_75t_SL \i56/i435  (.A(\i56/n33 ),
    .B(\i56/n27 ),
    .Y(\i56/n71 ));
 AND2x4_ASAP7_75t_SL \i56/i436  (.A(\i56/n36 ),
    .B(\i56/n37 ),
    .Y(\i56/n69 ));
 AND2x4_ASAP7_75t_SL \i56/i437  (.A(\i56/n33 ),
    .B(\i56/n37 ),
    .Y(\i56/n67 ));
 INVx2_ASAP7_75t_SL \i56/i438  (.A(\i56/n64 ),
    .Y(\i56/n63 ));
 INVx2_ASAP7_75t_SL \i56/i439  (.A(\i56/n59 ),
    .Y(\i56/n58 ));
 NAND4xp25_ASAP7_75t_SL \i56/i44  (.A(\i56/n381 ),
    .B(\i56/n317 ),
    .C(\i56/n242 ),
    .D(\i56/n281 ),
    .Y(\i56/n445 ));
 INVx3_ASAP7_75t_SL \i56/i440  (.A(\i56/n55 ),
    .Y(\i56/n54 ));
 INVx2_ASAP7_75t_SL \i56/i441  (.A(\i56/n53 ),
    .Y(\i56/n52 ));
 INVx3_ASAP7_75t_SL \i56/i442  (.A(\i56/n51 ),
    .Y(\i56/n50 ));
 INVx3_ASAP7_75t_SL \i56/i443  (.A(\i56/n49 ),
    .Y(\i56/n48 ));
 INVx3_ASAP7_75t_SL \i56/i444  (.A(\i56/n46 ),
    .Y(\i56/n45 ));
 INVx2_ASAP7_75t_SL \i56/i445  (.A(\i56/n44 ),
    .Y(\i56/n43 ));
 INVx3_ASAP7_75t_SL \i56/i446  (.A(\i56/n42 ),
    .Y(\i56/n41 ));
 INVx3_ASAP7_75t_SL \i56/i447  (.A(\i56/n40 ),
    .Y(\i56/n39 ));
 AND2x4_ASAP7_75t_SL \i56/i448  (.A(\i56/n23 ),
    .B(\i56/n35 ),
    .Y(\i56/n65 ));
 AND2x4_ASAP7_75t_SL \i56/i449  (.A(\i56/n25 ),
    .B(\i56/n533 ),
    .Y(\i56/n64 ));
 NOR2xp33_ASAP7_75t_SL \i56/i45  (.A(\i56/n419 ),
    .B(\i56/n396 ),
    .Y(\i56/n444 ));
 NAND2x1p5_ASAP7_75t_SL \i56/i450  (.A(\i56/n34 ),
    .B(\i56/n516 ),
    .Y(\i56/n62 ));
 AND2x4_ASAP7_75t_SL \i56/i451  (.A(\i56/n33 ),
    .B(\i56/n26 ),
    .Y(\i56/n60 ));
 AND2x4_ASAP7_75t_SL \i56/i452  (.A(\i56/n28 ),
    .B(\i56/n27 ),
    .Y(\i56/n59 ));
 NAND2xp5_ASAP7_75t_SL \i56/i453  (.A(\i56/n517 ),
    .B(\i56/n532 ),
    .Y(\i56/n57 ));
 AND4x1_ASAP7_75t_SL \i56/i454  (.A(n9[6]),
    .B(\i56/n0 ),
    .C(\i56/n3 ),
    .D(n9[4]),
    .Y(\i56/n56 ));
 OR2x6_ASAP7_75t_SL \i56/i455  (.A(\i56/n30 ),
    .B(\i56/n24 ),
    .Y(\i56/n55 ));
 AND2x4_ASAP7_75t_SL \i56/i456  (.A(\i56/n38 ),
    .B(\i56/n517 ),
    .Y(\i56/n53 ));
 AND2x4_ASAP7_75t_SL \i56/i457  (.A(\i56/n532 ),
    .B(\i56/n34 ),
    .Y(\i56/n51 ));
 AND2x4_ASAP7_75t_SL \i56/i458  (.A(\i56/n32 ),
    .B(\i56/n29 ),
    .Y(\i56/n49 ));
 AND2x4_ASAP7_75t_SL \i56/i459  (.A(\i56/n22 ),
    .B(\i56/n26 ),
    .Y(\i56/n47 ));
 NAND3xp33_ASAP7_75t_SL \i56/i46  (.A(\i56/n362 ),
    .B(\i56/n352 ),
    .C(\i56/n288 ),
    .Y(\i56/n443 ));
 AND2x4_ASAP7_75t_SL \i56/i460  (.A(\i56/n35 ),
    .B(\i56/n28 ),
    .Y(\i56/n46 ));
 AND2x4_ASAP7_75t_SL \i56/i461  (.A(\i56/n35 ),
    .B(\i56/n33 ),
    .Y(\i56/n44 ));
 AND2x4_ASAP7_75t_SL \i56/i462  (.A(\i56/n37 ),
    .B(\i56/n28 ),
    .Y(\i56/n42 ));
 AND2x4_ASAP7_75t_SL \i56/i463  (.A(\i56/n38 ),
    .B(\i56/n34 ),
    .Y(\i56/n40 ));
 AND2x2_ASAP7_75t_SL \i56/i464  (.A(n9[1]),
    .B(n9[0]),
    .Y(\i56/n32 ));
 AND2x2_ASAP7_75t_SL \i56/i465  (.A(n9[5]),
    .B(\i56/n18 ),
    .Y(\i56/n38 ));
 AND2x2_ASAP7_75t_SL \i56/i466  (.A(\i56/n21 ),
    .B(\i56/n17 ),
    .Y(\i56/n37 ));
 AND2x2_ASAP7_75t_SL \i56/i467  (.A(n9[2]),
    .B(n9[0]),
    .Y(\i56/n36 ));
 AND2x2_ASAP7_75t_SL \i56/i468  (.A(n9[3]),
    .B(n9[1]),
    .Y(\i56/n35 ));
 AND2x4_ASAP7_75t_SL \i56/i469  (.A(n9[7]),
    .B(\i56/n19 ),
    .Y(\i56/n34 ));
 NAND3xp33_ASAP7_75t_SL \i56/i47  (.A(\i56/n381 ),
    .B(\i56/n363 ),
    .C(\i56/n349 ),
    .Y(\i56/n442 ));
 AND2x4_ASAP7_75t_L \i56/i470  (.A(\i56/n20 ),
    .B(\i56/n16 ),
    .Y(\i56/n33 ));
 INVx1_ASAP7_75t_SL \i56/i471  (.A(\i56/n30 ),
    .Y(\i56/n31 ));
 NAND2xp5_ASAP7_75t_SL \i56/i472  (.A(n9[3]),
    .B(\i56/n20 ),
    .Y(\i56/n24 ));
 NOR2xp33_ASAP7_75t_SL \i56/i473  (.A(\i56/n16 ),
    .B(n9[2]),
    .Y(\i56/n23 ));
 NOR2xp33_ASAP7_75t_SL \i56/i474  (.A(\i56/n20 ),
    .B(n9[0]),
    .Y(\i56/n22 ));
 OR2x2_ASAP7_75t_SL \i56/i475  (.A(\i56/n16 ),
    .B(n9[1]),
    .Y(\i56/n30 ));
 AND2x2_ASAP7_75t_SL \i56/i476  (.A(\i56/n21 ),
    .B(\i56/n20 ),
    .Y(\i56/n29 ));
 AND2x2_ASAP7_75t_SL \i56/i477  (.A(n9[2]),
    .B(\i56/n16 ),
    .Y(\i56/n28 ));
 AND2x2_ASAP7_75t_SL \i56/i478  (.A(n9[1]),
    .B(\i56/n21 ),
    .Y(\i56/n27 ));
 AND2x2_ASAP7_75t_SL \i56/i479  (.A(n9[3]),
    .B(\i56/n17 ),
    .Y(\i56/n26 ));
 NOR3xp33_ASAP7_75t_SL \i56/i48  (.A(\i56/n330 ),
    .B(\i56/n496 ),
    .C(\i56/n369 ),
    .Y(\i56/n457 ));
 AND2x2_ASAP7_75t_SL \i56/i480  (.A(n9[5]),
    .B(n9[4]),
    .Y(\i56/n25 ));
 INVx3_ASAP7_75t_SL \i56/i481  (.A(n9[7]),
    .Y(\i56/n3 ));
 INVx2_ASAP7_75t_SL \i56/i482  (.A(n9[3]),
    .Y(\i56/n21 ));
 INVx4_ASAP7_75t_SL \i56/i483  (.A(n9[2]),
    .Y(\i56/n20 ));
 INVx1_ASAP7_75t_SL \i56/i484  (.A(n9[6]),
    .Y(\i56/n19 ));
 INVx2_ASAP7_75t_SL \i56/i485  (.A(n9[4]),
    .Y(\i56/n18 ));
 INVx2_ASAP7_75t_SL \i56/i486  (.A(n9[1]),
    .Y(\i56/n17 ));
 INVx3_ASAP7_75t_SL \i56/i487  (.A(n9[0]),
    .Y(\i56/n16 ));
 AND2x2_ASAP7_75t_SL \i56/i488  (.A(\i56/n531 ),
    .B(\i56/n15 ),
    .Y(\i56/n2 ));
 INVx2_ASAP7_75t_SL \i56/i489  (.A(\i56/n65 ),
    .Y(\i56/n483 ));
 NAND2xp5_ASAP7_75t_SL \i56/i49  (.A(\i56/n347 ),
    .B(\i56/n420 ),
    .Y(\i56/n455 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i56/i490  (.A1(\i56/n78 ),
    .A2(\i56/n484 ),
    .B(\i56/n1 ),
    .C(\i56/n73 ),
    .Y(\i56/n485 ));
 NAND2x1_ASAP7_75t_SL \i56/i491  (.A(\i56/n41 ),
    .B(\i56/n483 ),
    .Y(\i56/n484 ));
 NAND2xp5_ASAP7_75t_SL \i56/i492  (.A(\i56/n87 ),
    .B(\i56/n484 ),
    .Y(\i56/n486 ));
 OAI31xp33_ASAP7_75t_SL \i56/i493  (.A1(\i56/n484 ),
    .A2(\i56/n73 ),
    .A3(\i56/n60 ),
    .B(\i56/n489 ),
    .Y(\i56/n487 ));
 AND2x2_ASAP7_75t_SL \i56/i494  (.A(n9[7]),
    .B(n9[6]),
    .Y(\i56/n488 ));
 NAND2xp5_ASAP7_75t_SL \i56/i495  (.A(\i56/n489 ),
    .B(\i56/n44 ),
    .Y(\i56/n490 ));
 AND2x4_ASAP7_75t_SL \i56/i496  (.A(\i56/n488 ),
    .B(\i56/n532 ),
    .Y(\i56/n489 ));
 NAND2xp5_ASAP7_75t_SL \i56/i497  (.A(\i56/n49 ),
    .B(\i56/n489 ),
    .Y(\i56/n491 ));
 NOR2xp33_ASAP7_75t_SL \i56/i498  (.A(\i56/n489 ),
    .B(\i56/n1 ),
    .Y(\i56/n492 ));
 NAND2xp5_ASAP7_75t_SL \i56/i499  (.A(\i56/n78 ),
    .B(\i56/n489 ),
    .Y(\i56/n493 ));
 AND5x2_ASAP7_75t_SL \i56/i5  (.A(\i56/n461 ),
    .B(\i56/n460 ),
    .C(\i56/n428 ),
    .D(\i56/n462 ),
    .E(\i56/n438 ),
    .Y(n8[1]));
 NAND2xp5_ASAP7_75t_SL \i56/i50  (.A(\i56/n362 ),
    .B(\i56/n394 ),
    .Y(\i56/n454 ));
 NAND2xp5_ASAP7_75t_SL \i56/i500  (.A(\i56/n89 ),
    .B(\i56/n489 ),
    .Y(\i56/n494 ));
 NAND2xp5_ASAP7_75t_SL \i56/i501  (.A(\i56/n489 ),
    .B(\i56/n67 ),
    .Y(\i56/n495 ));
 AO22x1_ASAP7_75t_SL \i56/i502  (.A1(\i56/n64 ),
    .A2(\i56/n69 ),
    .B1(\i56/n489 ),
    .B2(\i56/n47 ),
    .Y(\i56/n496 ));
 AOI22xp5_ASAP7_75t_SL \i56/i503  (.A1(\i56/n54 ),
    .A2(\i56/n87 ),
    .B1(\i56/n489 ),
    .B2(\i56/n80 ),
    .Y(\i56/n497 ));
 AOI22xp5_ASAP7_75t_SL \i56/i504  (.A1(\i56/n84 ),
    .A2(\i56/n69 ),
    .B1(\i56/n489 ),
    .B2(\i56/n47 ),
    .Y(\i56/n498 ));
 AOI222xp33_ASAP7_75t_R \i56/i505  (.A1(\i56/n71 ),
    .A2(\i56/n77 ),
    .B1(\i56/n60 ),
    .B2(\i56/n489 ),
    .C1(\i56/n47 ),
    .C2(\i56/n82 ),
    .Y(\i56/n499 ));
 AOI222xp33_ASAP7_75t_SL \i56/i506  (.A1(\i56/n59 ),
    .A2(\i56/n100 ),
    .B1(\i56/n71 ),
    .B2(\i56/n489 ),
    .C1(\i56/n73 ),
    .C2(\i56/n40 ),
    .Y(\i56/n500 ));
 INVx3_ASAP7_75t_SL \i56/i507  (.A(\i56/n489 ),
    .Y(\i56/n501 ));
 OAI211xp5_ASAP7_75t_SL \i56/i508  (.A1(\i56/n505 ),
    .A2(\i56/n159 ),
    .B(\i56/n11 ),
    .C(\i56/n185 ),
    .Y(\i56/n502 ));
 OR2x2_ASAP7_75t_SL \i56/i509  (.A(n9[7]),
    .B(n9[6]),
    .Y(\i56/n503 ));
 INVx1_ASAP7_75t_SL \i56/i51  (.A(\i56/n440 ),
    .Y(\i56/n441 ));
 NAND2xp33_ASAP7_75t_SL \i56/i510  (.A(\i56/n50 ),
    .B(\i56/n505 ),
    .Y(\i56/n506 ));
 OR2x6_ASAP7_75t_SL \i56/i511  (.A(\i56/n503 ),
    .B(\i56/n504 ),
    .Y(\i56/n505 ));
 INVx2_ASAP7_75t_SL \i56/i512  (.A(\i56/n38 ),
    .Y(\i56/n504 ));
 NOR2xp67_ASAP7_75t_SL \i56/i513  (.A(\i56/n505 ),
    .B(\i56/n4 ),
    .Y(\i56/n507 ));
 OAI22xp5_ASAP7_75t_SL \i56/i514  (.A1(\i56/n55 ),
    .A2(\i56/n505 ),
    .B1(\i56/n88 ),
    .B2(\i56/n74 ),
    .Y(\i56/n508 ));
 OAI22xp5_ASAP7_75t_SL \i56/i515  (.A1(\i56/n50 ),
    .A2(\i56/n41 ),
    .B1(\i56/n48 ),
    .B2(\i56/n505 ),
    .Y(\i56/n509 ));
 OAI22xp5_ASAP7_75t_SL \i56/i516  (.A1(\i56/n505 ),
    .A2(\i56/n66 ),
    .B1(\i56/n74 ),
    .B2(\i56/n41 ),
    .Y(\i56/n510 ));
 OAI22xp5_ASAP7_75t_SL \i56/i517  (.A1(\i56/n505 ),
    .A2(\i56/n171 ),
    .B1(\i56/n86 ),
    .B2(\i56/n66 ),
    .Y(\i56/n511 ));
 OAI222xp33_ASAP7_75t_SL \i56/i518  (.A1(\i56/n74 ),
    .A2(\i56/n79 ),
    .B1(\i56/n41 ),
    .B2(\i56/n505 ),
    .C1(\i56/n39 ),
    .C2(\i56/n88 ),
    .Y(\i56/n512 ));
 OAI211xp5_ASAP7_75t_SL \i56/i519  (.A1(\i56/n68 ),
    .A2(\i56/n505 ),
    .B(\i56/n190 ),
    .C(\i56/n494 ),
    .Y(\i56/n513 ));
 INVxp67_ASAP7_75t_SL \i56/i52  (.A(\i56/n438 ),
    .Y(\i56/n439 ));
 INVx3_ASAP7_75t_SL \i56/i520  (.A(\i56/n505 ),
    .Y(\i56/n514 ));
 OAI22x1_ASAP7_75t_SL \i56/i521  (.A1(\i56/n45 ),
    .A2(\i56/n505 ),
    .B1(\i56/n86 ),
    .B2(\i56/n48 ),
    .Y(\i56/n515 ));
 AND2x2_ASAP7_75t_SL \i56/i522  (.A(\i56/n0 ),
    .B(\i56/n18 ),
    .Y(\i56/n516 ));
 AND2x2_ASAP7_75t_SL \i56/i523  (.A(\i56/n3 ),
    .B(n9[6]),
    .Y(\i56/n517 ));
 INVx2_ASAP7_75t_SL \i56/i524  (.A(\i56/n518 ),
    .Y(\i56/n519 ));
 AND2x4_ASAP7_75t_SL \i56/i525  (.A(\i56/n516 ),
    .B(\i56/n517 ),
    .Y(\i56/n518 ));
 AOI221xp5_ASAP7_75t_SL \i56/i526  (.A1(\i56/n175 ),
    .A2(\i56/n80 ),
    .B1(\i56/n518 ),
    .B2(\i56/n67 ),
    .C(\i56/n95 ),
    .Y(\i56/n520 ));
 O2A1O1Ixp5_ASAP7_75t_SL \i56/i527  (.A1(\i56/n73 ),
    .A2(\i56/n69 ),
    .B(\i56/n518 ),
    .C(\i56/n508 ),
    .Y(\i56/n521 ));
 AOI22xp5_ASAP7_75t_SL \i56/i528  (.A1(\i56/n49 ),
    .A2(\i56/n518 ),
    .B1(\i56/n54 ),
    .B2(\i56/n64 ),
    .Y(\i56/n522 ));
 AOI22xp5_ASAP7_75t_SL \i56/i529  (.A1(\i56/n518 ),
    .A2(\i56/n60 ),
    .B1(\i56/n47 ),
    .B2(\i56/n53 ),
    .Y(\i56/n523 ));
 NAND3xp33_ASAP7_75t_L \i56/i53  (.A(\i56/n376 ),
    .B(\i56/n338 ),
    .C(\i56/n387 ),
    .Y(\i56/n437 ));
 AOI22xp5_ASAP7_75t_SL \i56/i530  (.A1(\i56/n1 ),
    .A2(\i56/n44 ),
    .B1(\i56/n518 ),
    .B2(\i56/n69 ),
    .Y(\i56/n524 ));
 NAND2xp5_ASAP7_75t_SL \i56/i531  (.A(\i56/n65 ),
    .B(\i56/n518 ),
    .Y(\i56/n525 ));
 NAND2xp5_ASAP7_75t_SL \i56/i532  (.A(\i56/n73 ),
    .B(\i56/n518 ),
    .Y(\i56/n526 ));
 NOR2xp33_ASAP7_75t_SL \i56/i533  (.A(\i56/n85 ),
    .B(\i56/n518 ),
    .Y(\i56/n527 ));
 NAND2xp5_ASAP7_75t_SL \i56/i534  (.A(\i56/n80 ),
    .B(\i56/n518 ),
    .Y(\i56/n528 ));
 NAND2xp5_ASAP7_75t_SL \i56/i535  (.A(\i56/n518 ),
    .B(\i56/n42 ),
    .Y(\i56/n529 ));
 NAND2xp5_ASAP7_75t_SL \i56/i536  (.A(\i56/n71 ),
    .B(\i56/n518 ),
    .Y(\i56/n530 ));
 NAND2xp5_ASAP7_75t_SL \i56/i537  (.A(\i56/n46 ),
    .B(\i56/n518 ),
    .Y(\i56/n531 ));
 AND2x2_ASAP7_75t_SL \i56/i538  (.A(n9[4]),
    .B(\i56/n0 ),
    .Y(\i56/n532 ));
 INVx3_ASAP7_75t_SL \i56/i539  (.A(\i56/n503 ),
    .Y(\i56/n533 ));
 NAND3xp33_ASAP7_75t_L \i56/i54  (.A(\i56/n384 ),
    .B(\i56/n531 ),
    .C(\i56/n15 ),
    .Y(\i56/n436 ));
 AOI22xp33_ASAP7_75t_SL \i56/i540  (.A1(\i56/n534 ),
    .A2(\i56/n73 ),
    .B1(\i56/n80 ),
    .B2(\i56/n518 ),
    .Y(\i56/n535 ));
 AND2x4_ASAP7_75t_SL \i56/i541  (.A(\i56/n532 ),
    .B(\i56/n533 ),
    .Y(\i56/n534 ));
 INVx2_ASAP7_75t_SL \i56/i542  (.A(\i56/n534 ),
    .Y(\i56/n536 ));
 AOI222xp33_ASAP7_75t_SL \i56/i543  (.A1(\i56/n534 ),
    .A2(\i56/n71 ),
    .B1(\i56/n42 ),
    .B2(\i56/n53 ),
    .C1(\i56/n64 ),
    .C2(\i56/n49 ),
    .Y(\i56/n537 ));
 AOI222xp33_ASAP7_75t_SL \i56/i544  (.A1(\i56/n65 ),
    .A2(\i56/n534 ),
    .B1(\i56/n85 ),
    .B2(\i56/n49 ),
    .C1(\i56/n75 ),
    .C2(\i56/n65 ),
    .Y(\i56/n538 ));
 AOI222xp33_ASAP7_75t_SL \i56/i545  (.A1(\i56/n120 ),
    .A2(\i56/n46 ),
    .B1(\i56/n67 ),
    .B2(\i56/n85 ),
    .C1(\i56/n69 ),
    .C2(\i56/n534 ),
    .Y(\i56/n539 ));
 AOI221xp5_ASAP7_75t_SL \i56/i546  (.A1(\i56/n200 ),
    .A2(\i56/n64 ),
    .B1(\i56/n534 ),
    .B2(\i56/n71 ),
    .C(\i56/n134 ),
    .Y(\i56/n540 ));
 AOI22xp5_ASAP7_75t_SL \i56/i547  (.A1(\i56/n60 ),
    .A2(\i56/n51 ),
    .B1(\i56/n534 ),
    .B2(\i56/n59 ),
    .Y(\i56/n541 ));
 AOI22xp5_ASAP7_75t_SL \i56/i548  (.A1(\i56/n67 ),
    .A2(\i56/n534 ),
    .B1(\i56/n89 ),
    .B2(\i56/n82 ),
    .Y(\i56/n542 ));
 AO22x1_ASAP7_75t_SL \i56/i549  (.A1(\i56/n53 ),
    .A2(\i56/n67 ),
    .B1(\i56/n80 ),
    .B2(\i56/n534 ),
    .Y(\i56/n543 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i56/i55  (.A1(\i56/n62 ),
    .A2(\i56/n52 ),
    .B(\i56/n485 ),
    .C(\i56/n395 ),
    .Y(\i56/n435 ));
 AND2x2_ASAP7_75t_SL \i56/i550  (.A(\i56/n44 ),
    .B(\i56/n534 ),
    .Y(\i56/n544 ));
 NAND2xp5_ASAP7_75t_SL \i56/i551  (.A(\i56/n46 ),
    .B(\i56/n534 ),
    .Y(\i56/n545 ));
 AND2x2_ASAP7_75t_SL \i56/i552  (.A(\i56/n534 ),
    .B(\i56/n78 ),
    .Y(\i56/n546 ));
 NAND2xp5_ASAP7_75t_SL \i56/i553  (.A(\i56/n49 ),
    .B(\i56/n534 ),
    .Y(\i56/n547 ));
 INVx5_ASAP7_75t_SL \i56/i554  (.A(\i56/n84 ),
    .Y(\i56/n83 ));
 INVx5_ASAP7_75t_SL \i56/i555  (.A(\i56/n60 ),
    .Y(\i56/n61 ));
 INVx3_ASAP7_75t_SL \i56/i556  (.A(\i56/n47 ),
    .Y(\i56/n548 ));
 INVx3_ASAP7_75t_SL \i56/i557  (.A(\i56/n85 ),
    .Y(\i56/n549 ));
 NOR2xp67_ASAP7_75t_SL \i56/i558  (.A(\i56/n515 ),
    .B(\i56/n550 ),
    .Y(\i56/n551 ));
 OAI22x1_ASAP7_75t_SL \i56/i559  (.A1(\i56/n83 ),
    .A2(\i56/n61 ),
    .B1(\i56/n548 ),
    .B2(\i56/n549 ),
    .Y(\i56/n550 ));
 NAND2xp33_ASAP7_75t_SL \i56/i56  (.A(\i56/n401 ),
    .B(\i56/n552 ),
    .Y(\i56/n434 ));
 NOR4xp25_ASAP7_75t_SL \i56/i560  (.A(\i56/n372 ),
    .B(\i56/n330 ),
    .C(\i56/n221 ),
    .D(\i56/n550 ),
    .Y(\i56/n552 ));
 NOR4xp25_ASAP7_75t_SL \i56/i561  (.A(\i56/n375 ),
    .B(\i56/n299 ),
    .C(\i56/n131 ),
    .D(\i56/n226 ),
    .Y(\i56/n553 ));
 AND3x1_ASAP7_75t_SL \i56/i562  (.A(\i56/n11 ),
    .B(\i56/n150 ),
    .C(\i56/n529 ),
    .Y(\i56/n554 ));
 AND4x1_ASAP7_75t_SL \i56/i563  (.A(\i56/n197 ),
    .B(\i56/n196 ),
    .C(\i56/n149 ),
    .D(\i56/n12 ),
    .Y(\i56/n555 ));
 NOR2xp33_ASAP7_75t_SL \i56/i564  (.A(\i56/n556 ),
    .B(\i56/n231 ),
    .Y(\i56/n557 ));
 OAI21xp5_ASAP7_75t_SL \i56/i565  (.A1(\i56/n74 ),
    .A2(\i56/n4 ),
    .B(\i56/n495 ),
    .Y(\i56/n556 ));
 NOR2xp33_ASAP7_75t_SL \i56/i57  (.A(\i56/n379 ),
    .B(\i56/n397 ),
    .Y(\i56/n433 ));
 NAND5xp2_ASAP7_75t_SL \i56/i58  (.A(\i56/n333 ),
    .B(\i56/n294 ),
    .C(\i56/n284 ),
    .D(\i56/n305 ),
    .E(\i56/n313 ),
    .Y(\i56/n432 ));
 NOR3xp33_ASAP7_75t_SL \i56/i59  (.A(\i56/n348 ),
    .B(\i56/n261 ),
    .C(\i56/n319 ),
    .Y(\i56/n431 ));
 NOR2xp33_ASAP7_75t_SL \i56/i6  (.A(\i56/n451 ),
    .B(\i56/n481 ),
    .Y(\i56/n482 ));
 NAND2xp33_ASAP7_75t_SL \i56/i60  (.A(\i56/n378 ),
    .B(\i56/n401 ),
    .Y(\i56/n430 ));
 NAND4xp25_ASAP7_75t_SL \i56/i61  (.A(\i56/n388 ),
    .B(\i56/n363 ),
    .C(\i56/n290 ),
    .D(\i56/n557 ),
    .Y(\i56/n429 ));
 NOR3xp33_ASAP7_75t_SL \i56/i62  (.A(\i56/n400 ),
    .B(\i56/n360 ),
    .C(\i56/n383 ),
    .Y(\i56/n428 ));
 NAND5xp2_ASAP7_75t_SL \i56/i63  (.A(\i56/n368 ),
    .B(\i56/n334 ),
    .C(\i56/n329 ),
    .D(\i56/n215 ),
    .E(\i56/n298 ),
    .Y(\i56/n427 ));
 NAND5xp2_ASAP7_75t_SL \i56/i64  (.A(\i56/n356 ),
    .B(\i56/n326 ),
    .C(\i56/n302 ),
    .D(\i56/n300 ),
    .E(\i56/n551 ),
    .Y(\i56/n426 ));
 NOR4xp25_ASAP7_75t_SL \i56/i65  (.A(\i56/n353 ),
    .B(\i56/n354 ),
    .C(\i56/n543 ),
    .D(\i56/n191 ),
    .Y(\i56/n425 ));
 NAND2xp33_ASAP7_75t_SL \i56/i66  (.A(\i56/n405 ),
    .B(\i56/n382 ),
    .Y(\i56/n424 ));
 NAND4xp25_ASAP7_75t_SL \i56/i67  (.A(\i56/n387 ),
    .B(\i56/n359 ),
    .C(\i56/n390 ),
    .D(\i56/n312 ),
    .Y(\i56/n440 ));
 NOR3x1_ASAP7_75t_SL \i56/i68  (.A(\i56/n364 ),
    .B(\i56/n332 ),
    .C(\i56/n373 ),
    .Y(\i56/n438 ));
 INVxp67_ASAP7_75t_SL \i56/i69  (.A(\i56/n422 ),
    .Y(\i56/n423 ));
 AND4x2_ASAP7_75t_SL \i56/i7  (.A(\i56/n471 ),
    .B(\i56/n479 ),
    .C(\i56/n478 ),
    .D(\i56/n425 ),
    .Y(n8[5]));
 INVx1_ASAP7_75t_SL \i56/i70  (.A(\i56/n418 ),
    .Y(\i56/n419 ));
 INVxp67_ASAP7_75t_SL \i56/i71  (.A(\i56/n416 ),
    .Y(\i56/n417 ));
 INVxp67_ASAP7_75t_SL \i56/i72  (.A(\i56/n414 ),
    .Y(\i56/n415 ));
 NOR3xp33_ASAP7_75t_SL \i56/i73  (.A(\i56/n377 ),
    .B(\i56/n14 ),
    .C(\i56/n229 ),
    .Y(\i56/n413 ));
 NAND3xp33_ASAP7_75t_SL \i56/i74  (.A(\i56/n260 ),
    .B(\i56/n487 ),
    .C(\i56/n278 ),
    .Y(\i56/n412 ));
 NAND2xp5_ASAP7_75t_SL \i56/i75  (.A(\i56/n365 ),
    .B(\i56/n380 ),
    .Y(\i56/n411 ));
 NOR2xp33_ASAP7_75t_SL \i56/i76  (.A(\i56/n389 ),
    .B(\i56/n355 ),
    .Y(\i56/n410 ));
 NOR2xp33_ASAP7_75t_SL \i56/i77  (.A(\i56/n346 ),
    .B(\i56/n289 ),
    .Y(\i56/n409 ));
 NOR5xp2_ASAP7_75t_SL \i56/i78  (.A(\i56/n280 ),
    .B(\i56/n496 ),
    .C(\i56/n543 ),
    .D(\i56/n256 ),
    .E(\i56/n254 ),
    .Y(\i56/n408 ));
 NOR2xp33_ASAP7_75t_SL \i56/i79  (.A(\i56/n331 ),
    .B(\i56/n357 ),
    .Y(\i56/n407 ));
 AND3x4_ASAP7_75t_SL \i56/i8  (.A(\i56/n473 ),
    .B(\i56/n477 ),
    .C(\i56/n441 ),
    .Y(n8[0]));
 AOI211xp5_ASAP7_75t_SL \i56/i80  (.A1(\i56/n318 ),
    .A2(\i56/n110 ),
    .B(\i56/n272 ),
    .C(\i56/n230 ),
    .Y(\i56/n406 ));
 NAND2xp5_ASAP7_75t_SL \i56/i81  (.A(\i56/n283 ),
    .B(\i56/n381 ),
    .Y(\i56/n422 ));
 NAND3xp33_ASAP7_75t_SL \i56/i82  (.A(\i56/n339 ),
    .B(\i56/n361 ),
    .C(\i56/n311 ),
    .Y(\i56/n421 ));
 NOR2x1_ASAP7_75t_SL \i56/i83  (.A(\i56/n370 ),
    .B(\i56/n293 ),
    .Y(\i56/n420 ));
 AND3x1_ASAP7_75t_SL \i56/i84  (.A(\i56/n486 ),
    .B(\i56/n295 ),
    .C(\i56/n273 ),
    .Y(\i56/n418 ));
 NAND3xp33_ASAP7_75t_SL \i56/i85  (.A(\i56/n290 ),
    .B(\i56/n288 ),
    .C(\i56/n555 ),
    .Y(\i56/n416 ));
 NOR3x1_ASAP7_75t_SL \i56/i86  (.A(\i56/n292 ),
    .B(\i56/n315 ),
    .C(\i56/n224 ),
    .Y(\i56/n414 ));
 INVxp33_ASAP7_75t_SL \i56/i87  (.A(\i56/n402 ),
    .Y(\i56/n403 ));
 OAI211xp5_ASAP7_75t_SL \i56/i88  (.A1(\i56/n548 ),
    .A2(\i56/n183 ),
    .B(\i56/n308 ),
    .C(\i56/n246 ),
    .Y(\i56/n399 ));
 AOI211xp5_ASAP7_75t_SL \i56/i89  (.A1(\i56/n184 ),
    .A2(\i56/n49 ),
    .B(\i56/n270 ),
    .C(\i56/n513 ),
    .Y(\i56/n398 ));
 AND4x2_ASAP7_75t_SL \i56/i9  (.A(\i56/n466 ),
    .B(\i56/n467 ),
    .C(\i56/n463 ),
    .D(\i56/n464 ),
    .Y(n8[7]));
 NAND4xp25_ASAP7_75t_SL \i56/i90  (.A(\i56/n521 ),
    .B(\i56/n316 ),
    .C(\i56/n282 ),
    .D(\i56/n244 ),
    .Y(\i56/n397 ));
 NAND4xp25_ASAP7_75t_SL \i56/i91  (.A(\i56/n339 ),
    .B(\i56/n243 ),
    .C(\i56/n304 ),
    .D(\i56/n202 ),
    .Y(\i56/n396 ));
 NOR3xp33_ASAP7_75t_SL \i56/i92  (.A(\i56/n307 ),
    .B(\i56/n262 ),
    .C(\i56/n265 ),
    .Y(\i56/n395 ));
 NOR3xp33_ASAP7_75t_SL \i56/i93  (.A(\i56/n511 ),
    .B(\i56/n248 ),
    .C(\i56/n271 ),
    .Y(\i56/n405 ));
 NOR2xp67_ASAP7_75t_SL \i56/i94  (.A(\i56/n383 ),
    .B(\i56/n344 ),
    .Y(\i56/n394 ));
 NOR2xp33_ASAP7_75t_SL \i56/i95  (.A(\i56/n371 ),
    .B(\i56/n351 ),
    .Y(\i56/n393 ));
 NAND5xp2_ASAP7_75t_SL \i56/i96  (.A(\i56/n286 ),
    .B(\i56/n537 ),
    .C(\i56/n214 ),
    .D(\i56/n542 ),
    .E(\i56/n215 ),
    .Y(\i56/n404 ));
 NAND2xp5_ASAP7_75t_SL \i56/i97  (.A(\i56/n359 ),
    .B(\i56/n390 ),
    .Y(\i56/n392 ));
 NOR3xp33_ASAP7_75t_SL \i56/i98  (.A(\i56/n340 ),
    .B(\i56/n220 ),
    .C(\i56/n105 ),
    .Y(\i56/n402 ));
 NOR2xp33_ASAP7_75t_L \i56/i99  (.A(\i56/n342 ),
    .B(\i56/n325 ),
    .Y(\i56/n401 ));
 AOI22xp5_ASAP7_75t_SL i560 (.A1(n765),
    .A2(n506),
    .B1(n764),
    .B2(n507),
    .Y(n912));
 OAI22xp5_ASAP7_75t_SL i561 (.A1(n759),
    .A2(n803),
    .B1(n758),
    .B2(n802),
    .Y(n911));
 OAI22xp5_ASAP7_75t_SL i562 (.A1(n794),
    .A2(n756),
    .B1(n793),
    .B2(n757),
    .Y(n910));
 AOI22xp33_ASAP7_75t_SL i563 (.A1(n758),
    .A2(n1232),
    .B1(n777),
    .B2(n759),
    .Y(n909));
 AOI22xp5_ASAP7_75t_SL i564 (.A1(n757),
    .A2(n802),
    .B1(n756),
    .B2(n803),
    .Y(n908));
 OAI22xp5_ASAP7_75t_SL i565 (.A1(n478),
    .A2(n507),
    .B1(n477),
    .B2(n506),
    .Y(n907));
 AOI22xp5_ASAP7_75t_SL i566 (.A1(n497),
    .A2(n763),
    .B1(n498),
    .B2(n762),
    .Y(n906));
 OAI22xp5_ASAP7_75t_SL i567 (.A1(n493),
    .A2(n762),
    .B1(n492),
    .B2(n763),
    .Y(n905));
 AOI22xp5_ASAP7_75t_SL i568 (.A1(n763),
    .A2(n505),
    .B1(n762),
    .B2(n504),
    .Y(n904));
 OAI22xp5_ASAP7_75t_SL i569 (.A1(n1175),
    .A2(n572),
    .B1(n571),
    .B2(n792),
    .Y(n903));
 INVx1_ASAP7_75t_SL \i57/i0  (.A(n7[5]),
    .Y(\i57/n0 ));
 INVx2_ASAP7_75t_SL \i57/i1  (.A(n7[1]),
    .Y(\i57/n1 ));
 AND3x4_ASAP7_75t_SL \i57/i10  (.A(\i57/n474 ),
    .B(\i57/n478 ),
    .C(\i57/n444 ),
    .Y(n6[0]));
 INVxp33_ASAP7_75t_SL \i57/i100  (.A(\i57/n393 ),
    .Y(\i57/n394 ));
 INVxp67_ASAP7_75t_SL \i57/i101  (.A(\i57/n389 ),
    .Y(\i57/n390 ));
 NOR3xp33_ASAP7_75t_SL \i57/i102  (.A(\i57/n256 ),
    .B(\i57/n215 ),
    .C(\i57/n94 ),
    .Y(\i57/n385 ));
 OAI211xp5_ASAP7_75t_SL \i57/i103  (.A1(\i57/n66 ),
    .A2(\i57/n174 ),
    .B(\i57/n545 ),
    .C(\i57/n300 ),
    .Y(\i57/n384 ));
 NOR2xp33_ASAP7_75t_SL \i57/i104  (.A(\i57/n340 ),
    .B(\i57/n17 ),
    .Y(\i57/n383 ));
 OAI21xp5_ASAP7_75t_SL \i57/i105  (.A1(\i57/n57 ),
    .A2(\i57/n78 ),
    .B(\i57/n343 ),
    .Y(\i57/n382 ));
 NOR4xp25_ASAP7_75t_SL \i57/i106  (.A(\i57/n241 ),
    .B(\i57/n242 ),
    .C(\i57/n207 ),
    .D(\i57/n535 ),
    .Y(\i57/n381 ));
 NAND2xp33_ASAP7_75t_SL \i57/i107  (.A(\i57/n557 ),
    .B(\i57/n345 ),
    .Y(\i57/n380 ));
 NOR3xp33_ASAP7_75t_SL \i57/i108  (.A(\i57/n308 ),
    .B(\i57/n128 ),
    .C(\i57/n184 ),
    .Y(\i57/n379 ));
 NAND2xp5_ASAP7_75t_SL \i57/i109  (.A(\i57/n228 ),
    .B(\i57/n274 ),
    .Y(\i57/n378 ));
 AND4x2_ASAP7_75t_SL \i57/i11  (.A(\i57/n467 ),
    .B(\i57/n468 ),
    .C(\i57/n465 ),
    .D(\i57/n466 ),
    .Y(n6[7]));
 NOR2xp33_ASAP7_75t_L \i57/i110  (.A(\i57/n285 ),
    .B(\i57/n307 ),
    .Y(\i57/n395 ));
 OAI211xp5_ASAP7_75t_SL \i57/i111  (.A1(\i57/n48 ),
    .A2(\i57/n57 ),
    .B(\i57/n514 ),
    .C(\i57/n219 ),
    .Y(\i57/n377 ));
 NAND3xp33_ASAP7_75t_L \i57/i112  (.A(\i57/n258 ),
    .B(\i57/n493 ),
    .C(\i57/n310 ),
    .Y(\i57/n376 ));
 NAND2xp5_ASAP7_75t_SL \i57/i113  (.A(\i57/n509 ),
    .B(\i57/n514 ),
    .Y(\i57/n375 ));
 NAND2xp5_ASAP7_75t_L \i57/i114  (.A(\i57/n250 ),
    .B(\i57/n270 ),
    .Y(\i57/n374 ));
 NOR3xp33_ASAP7_75t_SL \i57/i115  (.A(\i57/n304 ),
    .B(\i57/n208 ),
    .C(\i57/n224 ),
    .Y(\i57/n373 ));
 NOR3xp33_ASAP7_75t_SL \i57/i116  (.A(\i57/n16 ),
    .B(\i57/n195 ),
    .C(\i57/n179 ),
    .Y(\i57/n372 ));
 NOR4xp25_ASAP7_75t_SL \i57/i117  (.A(\i57/n16 ),
    .B(\i57/n209 ),
    .C(\i57/n199 ),
    .D(\i57/n97 ),
    .Y(\i57/n371 ));
 AOI211x1_ASAP7_75t_SL \i57/i118  (.A1(\i57/n113 ),
    .A2(\i57/n74 ),
    .B(\i57/n237 ),
    .C(\i57/n229 ),
    .Y(\i57/n393 ));
 NOR3xp33_ASAP7_75t_SL \i57/i119  (.A(\i57/n263 ),
    .B(\i57/n128 ),
    .C(\i57/n245 ),
    .Y(\i57/n392 ));
 NAND4xp25_ASAP7_75t_SL \i57/i12  (.A(\i57/n459 ),
    .B(\i57/n397 ),
    .C(\i57/n387 ),
    .D(\i57/n489 ),
    .Y(\i57/n482 ));
 NOR2xp33_ASAP7_75t_L \i57/i120  (.A(\i57/n224 ),
    .B(\i57/n349 ),
    .Y(\i57/n370 ));
 NOR2x1_ASAP7_75t_SL \i57/i121  (.A(\i57/n272 ),
    .B(\i57/n337 ),
    .Y(\i57/n391 ));
 NOR2x1_ASAP7_75t_SL \i57/i122  (.A(\i57/n278 ),
    .B(\i57/n344 ),
    .Y(\i57/n389 ));
 NAND2xp5_ASAP7_75t_SL \i57/i123  (.A(\i57/n219 ),
    .B(\i57/n284 ),
    .Y(\i57/n388 ));
 NOR2xp67_ASAP7_75t_SL \i57/i124  (.A(\i57/n323 ),
    .B(\i57/n346 ),
    .Y(\i57/n387 ));
 NOR3x1_ASAP7_75t_SL \i57/i125  (.A(\i57/n271 ),
    .B(\i57/n256 ),
    .C(\i57/n230 ),
    .Y(\i57/n386 ));
 INVx1_ASAP7_75t_SL \i57/i126  (.A(\i57/n366 ),
    .Y(\i57/n367 ));
 NOR2xp33_ASAP7_75t_SL \i57/i127  (.A(\i57/n528 ),
    .B(\i57/n318 ),
    .Y(\i57/n365 ));
 NAND5xp2_ASAP7_75t_SL \i57/i128  (.A(\i57/n95 ),
    .B(\i57/n200 ),
    .C(\i57/n163 ),
    .D(\i57/n554 ),
    .E(\i57/n191 ),
    .Y(\i57/n364 ));
 NOR2xp33_ASAP7_75t_SL \i57/i129  (.A(\i57/n319 ),
    .B(\i57/n332 ),
    .Y(\i57/n363 ));
 NOR3xp33_ASAP7_75t_SL \i57/i13  (.A(\i57/n540 ),
    .B(\i57/n471 ),
    .C(\i57/n455 ),
    .Y(\i57/n481 ));
 OAI211xp5_ASAP7_75t_SL \i57/i130  (.A1(\i57/n48 ),
    .A2(\i57/n177 ),
    .B(\i57/n487 ),
    .C(\i57/n262 ),
    .Y(\i57/n362 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i57/i131  (.A1(\i57/n75 ),
    .A2(\i57/n193 ),
    .B(\i57/n8 ),
    .C(\i57/n254 ),
    .Y(\i57/n361 ));
 NAND3xp33_ASAP7_75t_SL \i57/i132  (.A(\i57/n265 ),
    .B(\i57/n510 ),
    .C(\i57/n238 ),
    .Y(\i57/n360 ));
 NOR3xp33_ASAP7_75t_SL \i57/i133  (.A(\i57/n275 ),
    .B(\i57/n223 ),
    .C(\i57/n231 ),
    .Y(\i57/n359 ));
 NAND3xp33_ASAP7_75t_L \i57/i134  (.A(\i57/n222 ),
    .B(\i57/n219 ),
    .C(\i57/n312 ),
    .Y(\i57/n358 ));
 NOR3xp33_ASAP7_75t_SL \i57/i135  (.A(\i57/n287 ),
    .B(\i57/n260 ),
    .C(\i57/n223 ),
    .Y(\i57/n357 ));
 AOI211xp5_ASAP7_75t_SL \i57/i136  (.A1(\i57/n526 ),
    .A2(\i57/n81 ),
    .B(\i57/n330 ),
    .C(\i57/n129 ),
    .Y(\i57/n356 ));
 OAI221xp5_ASAP7_75t_SL \i57/i137  (.A1(\i57/n174 ),
    .A2(\i57/n48 ),
    .B1(\i57/n116 ),
    .B2(\i57/n2 ),
    .C(\i57/n183 ),
    .Y(\i57/n355 ));
 NAND2xp33_ASAP7_75t_SL \i57/i138  (.A(\i57/n286 ),
    .B(\i57/n282 ),
    .Y(\i57/n354 ));
 NOR2xp33_ASAP7_75t_SL \i57/i139  (.A(\i57/n329 ),
    .B(\i57/n294 ),
    .Y(\i57/n353 ));
 AND2x2_ASAP7_75t_SL \i57/i14  (.A(\i57/n476 ),
    .B(\i57/n477 ),
    .Y(n6[2]));
 OAI221xp5_ASAP7_75t_SL \i57/i140  (.A1(\i57/n247 ),
    .A2(\i57/n92 ),
    .B1(\i57/n12 ),
    .B2(\i57/n84 ),
    .C(\i57/n206 ),
    .Y(\i57/n352 ));
 NAND4xp25_ASAP7_75t_SL \i57/i141  (.A(\i57/n210 ),
    .B(\i57/n548 ),
    .C(\i57/n550 ),
    .D(\i57/n201 ),
    .Y(\i57/n351 ));
 NOR2xp67_ASAP7_75t_SL \i57/i142  (.A(\i57/n296 ),
    .B(\i57/n305 ),
    .Y(\i57/n369 ));
 NAND2xp33_ASAP7_75t_L \i57/i143  (.A(\i57/n336 ),
    .B(\i57/n233 ),
    .Y(\i57/n350 ));
 NOR2x1_ASAP7_75t_SL \i57/i144  (.A(\i57/n314 ),
    .B(\i57/n333 ),
    .Y(\i57/n368 ));
 NAND2xp5_ASAP7_75t_SL \i57/i145  (.A(\i57/n277 ),
    .B(\i57/n221 ),
    .Y(\i57/n366 ));
 NOR2xp67_ASAP7_75t_SL \i57/i146  (.A(\i57/n276 ),
    .B(\i57/n283 ),
    .Y(\i57/n18 ));
 INVxp67_ASAP7_75t_SL \i57/i147  (.A(\i57/n346 ),
    .Y(\i57/n347 ));
 INVxp33_ASAP7_75t_SL \i57/i148  (.A(\i57/n344 ),
    .Y(\i57/n345 ));
 INVx1_ASAP7_75t_SL \i57/i149  (.A(\i57/n341 ),
    .Y(\i57/n342 ));
 NOR3xp33_ASAP7_75t_SL \i57/i15  (.A(\i57/n456 ),
    .B(\i57/n405 ),
    .C(\i57/n460 ),
    .Y(\i57/n480 ));
 INVxp67_ASAP7_75t_SL \i57/i150  (.A(\i57/n337 ),
    .Y(\i57/n338 ));
 INVxp67_ASAP7_75t_SL \i57/i151  (.A(\i57/n17 ),
    .Y(\i57/n336 ));
 INVxp67_ASAP7_75t_SL \i57/i152  (.A(\i57/n334 ),
    .Y(\i57/n335 ));
 NAND2xp5_ASAP7_75t_SL \i57/i153  (.A(\i57/n493 ),
    .B(\i57/n511 ),
    .Y(\i57/n333 ));
 NAND2xp33_ASAP7_75t_SL \i57/i154  (.A(\i57/n534 ),
    .B(\i57/n547 ),
    .Y(\i57/n332 ));
 AOI21xp5_ASAP7_75t_SL \i57/i155  (.A1(\i57/n181 ),
    .A2(\i57/n93 ),
    .B(\i57/n260 ),
    .Y(\i57/n331 ));
 OAI22xp5_ASAP7_75t_SL \i57/i156  (.A1(\i57/n111 ),
    .A2(\i57/n141 ),
    .B1(\i57/n86 ),
    .B2(\i57/n126 ),
    .Y(\i57/n330 ));
 NAND4xp25_ASAP7_75t_SL \i57/i157  (.A(\i57/n187 ),
    .B(\i57/n137 ),
    .C(\i57/n520 ),
    .D(\i57/n501 ),
    .Y(\i57/n329 ));
 NAND3xp33_ASAP7_75t_SL \i57/i158  (.A(\i57/n134 ),
    .B(\i57/n145 ),
    .C(\i57/n9 ),
    .Y(\i57/n328 ));
 NAND3xp33_ASAP7_75t_SL \i57/i159  (.A(\i57/n173 ),
    .B(\i57/n186 ),
    .C(\i57/n508 ),
    .Y(\i57/n327 ));
 NOR3xp33_ASAP7_75t_SL \i57/i16  (.A(\i57/n436 ),
    .B(\i57/n441 ),
    .C(\i57/n420 ),
    .Y(\i57/n479 ));
 OAI211xp5_ASAP7_75t_SL \i57/i160  (.A1(\i57/n68 ),
    .A2(\i57/n89 ),
    .B(\i57/n187 ),
    .C(\i57/n201 ),
    .Y(\i57/n326 ));
 NOR2xp33_ASAP7_75t_SL \i57/i161  (.A(\i57/n230 ),
    .B(\i57/n239 ),
    .Y(\i57/n325 ));
 OAI21xp5_ASAP7_75t_SL \i57/i162  (.A1(\i57/n86 ),
    .A2(\i57/n154 ),
    .B(\i57/n102 ),
    .Y(\i57/n324 ));
 NAND4xp25_ASAP7_75t_SL \i57/i163  (.A(\i57/n517 ),
    .B(\i57/n147 ),
    .C(\i57/n135 ),
    .D(\i57/n170 ),
    .Y(\i57/n323 ));
 AOI211xp5_ASAP7_75t_SL \i57/i164  (.A1(\i57/n45 ),
    .A2(\i57/n7 ),
    .B(\i57/n144 ),
    .C(\i57/n138 ),
    .Y(\i57/n322 ));
 NOR2xp33_ASAP7_75t_L \i57/i165  (.A(\i57/n213 ),
    .B(\i57/n252 ),
    .Y(\i57/n321 ));
 NOR2xp33_ASAP7_75t_L \i57/i166  (.A(\i57/n212 ),
    .B(\i57/n232 ),
    .Y(\i57/n320 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i57/i167  (.A1(\i57/n66 ),
    .A2(\i57/n44 ),
    .B(\i57/n50 ),
    .C(\i57/n255 ),
    .Y(\i57/n319 ));
 NAND3xp33_ASAP7_75t_SL \i57/i168  (.A(\i57/n250 ),
    .B(\i57/n550 ),
    .C(\i57/n503 ),
    .Y(\i57/n318 ));
 NOR3xp33_ASAP7_75t_SL \i57/i169  (.A(\i57/n236 ),
    .B(\i57/n150 ),
    .C(\i57/n202 ),
    .Y(\i57/n317 ));
 NOR3xp33_ASAP7_75t_SL \i57/i17  (.A(\i57/n446 ),
    .B(\i57/n448 ),
    .C(\i57/n431 ),
    .Y(\i57/n478 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i57/i170  (.A1(\i57/n63 ),
    .A2(\i57/n69 ),
    .B(\i57/n56 ),
    .C(\i57/n127 ),
    .Y(\i57/n316 ));
 NAND4xp25_ASAP7_75t_SL \i57/i171  (.A(\i57/n495 ),
    .B(\i57/n121 ),
    .C(\i57/n15 ),
    .D(\i57/n549 ),
    .Y(\i57/n315 ));
 OAI211xp5_ASAP7_75t_SL \i57/i172  (.A1(\i57/n58 ),
    .A2(\i57/n64 ),
    .B(\i57/n518 ),
    .C(\i57/n497 ),
    .Y(\i57/n314 ));
 AOI221xp5_ASAP7_75t_SL \i57/i173  (.A1(\i57/n166 ),
    .A2(\i57/n59 ),
    .B1(\i57/n53 ),
    .B2(\i57/n93 ),
    .C(\i57/n149 ),
    .Y(\i57/n313 ));
 NOR2xp33_ASAP7_75t_SL \i57/i174  (.A(\i57/n133 ),
    .B(\i57/n211 ),
    .Y(\i57/n312 ));
 OAI221xp5_ASAP7_75t_SL \i57/i175  (.A1(\i57/n44 ),
    .A2(\i57/n42 ),
    .B1(\i57/n52 ),
    .B2(\i57/n68 ),
    .C(\i57/n494 ),
    .Y(\i57/n349 ));
 AOI222xp33_ASAP7_75t_SL \i57/i176  (.A1(\i57/n6 ),
    .A2(\i57/n56 ),
    .B1(\i57/n77 ),
    .B2(\i57/n74 ),
    .C1(\i57/n63 ),
    .C2(\i57/n81 ),
    .Y(\i57/n348 ));
 NAND2xp5_ASAP7_75t_SL \i57/i177  (.A(\i57/n249 ),
    .B(\i57/n513 ),
    .Y(\i57/n346 ));
 OAI221xp5_ASAP7_75t_SL \i57/i178  (.A1(\i57/n64 ),
    .A2(\i57/n55 ),
    .B1(\i57/n530 ),
    .B2(\i57/n57 ),
    .C(\i57/n9 ),
    .Y(\i57/n344 ));
 OAI21xp5_ASAP7_75t_SL \i57/i179  (.A1(\i57/n59 ),
    .A2(\i57/n125 ),
    .B(\i57/n175 ),
    .Y(\i57/n343 ));
 NOR4xp25_ASAP7_75t_SL \i57/i18  (.A(\i57/n417 ),
    .B(\i57/n429 ),
    .C(\i57/n421 ),
    .D(\i57/n525 ),
    .Y(\i57/n477 ));
 NOR2xp33_ASAP7_75t_SL \i57/i180  (.A(\i57/n128 ),
    .B(\i57/n263 ),
    .Y(\i57/n311 ));
 NAND2xp5_ASAP7_75t_SL \i57/i181  (.A(\i57/n214 ),
    .B(\i57/n547 ),
    .Y(\i57/n341 ));
 NOR2xp33_ASAP7_75t_SL \i57/i182  (.A(\i57/n536 ),
    .B(\i57/n535 ),
    .Y(\i57/n310 ));
 NAND2xp5_ASAP7_75t_SL \i57/i183  (.A(\i57/n216 ),
    .B(\i57/n218 ),
    .Y(\i57/n340 ));
 NAND2xp5_ASAP7_75t_SL \i57/i184  (.A(\i57/n240 ),
    .B(\i57/n255 ),
    .Y(\i57/n339 ));
 OAI221xp5_ASAP7_75t_SL \i57/i185  (.A1(\i57/n508 ),
    .A2(\i57/n90 ),
    .B1(\i57/n70 ),
    .B2(\i57/n86 ),
    .C(\i57/n140 ),
    .Y(\i57/n337 ));
 NAND2xp5_ASAP7_75t_SL \i57/i186  (.A(\i57/n246 ),
    .B(\i57/n222 ),
    .Y(\i57/n17 ));
 NAND3xp33_ASAP7_75t_SL \i57/i187  (.A(\i57/n139 ),
    .B(\i57/n136 ),
    .C(\i57/n132 ),
    .Y(\i57/n16 ));
 NOR2xp33_ASAP7_75t_SL \i57/i188  (.A(\i57/n264 ),
    .B(\i57/n257 ),
    .Y(\i57/n309 ));
 OAI211xp5_ASAP7_75t_SL \i57/i189  (.A1(\i57/n80 ),
    .A2(\i57/n71 ),
    .B(\i57/n205 ),
    .C(\i57/n13 ),
    .Y(\i57/n334 ));
 NOR5xp2_ASAP7_75t_SL \i57/i19  (.A(\i57/n539 ),
    .B(\i57/n426 ),
    .C(\i57/n456 ),
    .D(\i57/n409 ),
    .E(\i57/n390 ),
    .Y(\i57/n476 ));
 INVxp67_ASAP7_75t_SL \i57/i190  (.A(\i57/n305 ),
    .Y(\i57/n306 ));
 INVxp67_ASAP7_75t_SL \i57/i191  (.A(\i57/n492 ),
    .Y(\i57/n304 ));
 INVxp67_ASAP7_75t_SL \i57/i192  (.A(\i57/n302 ),
    .Y(\i57/n303 ));
 INVx2_ASAP7_75t_SL \i57/i193  (.A(\i57/n300 ),
    .Y(\i57/n301 ));
 INVx1_ASAP7_75t_SL \i57/i194  (.A(\i57/n298 ),
    .Y(\i57/n299 ));
 OAI22xp5_ASAP7_75t_SL \i57/i195  (.A1(\i57/n530 ),
    .A2(\i57/n123 ),
    .B1(\i57/n75 ),
    .B2(\i57/n71 ),
    .Y(\i57/n296 ));
 AOI21xp5_ASAP7_75t_SL \i57/i196  (.A1(\i57/n109 ),
    .A2(\i57/n76 ),
    .B(\i57/n129 ),
    .Y(\i57/n295 ));
 OAI22xp5_ASAP7_75t_SL \i57/i197  (.A1(\i57/n57 ),
    .A2(\i57/n106 ),
    .B1(\i57/n55 ),
    .B2(\i57/n189 ),
    .Y(\i57/n294 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i57/i198  (.A1(\i57/n526 ),
    .A2(\i57/n67 ),
    .B(\i57/n74 ),
    .C(\i57/n99 ),
    .Y(\i57/n293 ));
 AOI21xp5_ASAP7_75t_SL \i57/i199  (.A1(\i57/n176 ),
    .A2(\i57/n526 ),
    .B(\i57/n243 ),
    .Y(\i57/n292 ));
 INVx3_ASAP7_75t_SL \i57/i2  (.A(\i57/n6 ),
    .Y(\i57/n2 ));
 NOR3xp33_ASAP7_75t_SL \i57/i20  (.A(\i57/n541 ),
    .B(\i57/n457 ),
    .C(\i57/n469 ),
    .Y(\i57/n475 ));
 AOI22xp5_ASAP7_75t_SL \i57/i200  (.A1(\i57/n51 ),
    .A2(\i57/n110 ),
    .B1(\i57/n79 ),
    .B2(\i57/n169 ),
    .Y(\i57/n291 ));
 AOI211xp5_ASAP7_75t_SL \i57/i201  (.A1(\i57/n51 ),
    .A2(\i57/n54 ),
    .B(\i57/n129 ),
    .C(\i57/n101 ),
    .Y(\i57/n290 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i57/i202  (.A1(\i57/n72 ),
    .A2(\i57/n69 ),
    .B(\i57/n65 ),
    .C(\i57/n227 ),
    .Y(\i57/n289 ));
 OAI22xp5_ASAP7_75t_SL \i57/i203  (.A1(\i57/n66 ),
    .A2(\i57/n165 ),
    .B1(\i57/n8 ),
    .B2(\i57/n164 ),
    .Y(\i57/n288 ));
 OAI22xp5_ASAP7_75t_SL \i57/i204  (.A1(\i57/n60 ),
    .A2(\i57/n157 ),
    .B1(\i57/n55 ),
    .B2(\i57/n75 ),
    .Y(\i57/n287 ));
 AND4x1_ASAP7_75t_SL \i57/i205  (.A(\i57/n135 ),
    .B(\i57/n11 ),
    .C(\i57/n14 ),
    .D(\i57/n140 ),
    .Y(\i57/n286 ));
 NAND4xp25_ASAP7_75t_SL \i57/i206  (.A(\i57/n130 ),
    .B(\i57/n152 ),
    .C(\i57/n118 ),
    .D(\i57/n496 ),
    .Y(\i57/n285 ));
 AOI222xp33_ASAP7_75t_SL \i57/i207  (.A1(\i57/n117 ),
    .A2(\i57/n49 ),
    .B1(\i57/n67 ),
    .B2(\i57/n85 ),
    .C1(\i57/n69 ),
    .C2(\i57/n91 ),
    .Y(\i57/n284 ));
 NAND4xp25_ASAP7_75t_SL \i57/i208  (.A(\i57/n139 ),
    .B(\i57/n137 ),
    .C(\i57/n197 ),
    .D(\i57/n136 ),
    .Y(\i57/n283 ));
 AOI22xp5_ASAP7_75t_SL \i57/i209  (.A1(\i57/n88 ),
    .A2(\i57/n105 ),
    .B1(\i57/n81 ),
    .B2(\i57/n119 ),
    .Y(\i57/n282 ));
 NOR3xp33_ASAP7_75t_SL \i57/i21  (.A(\i57/n438 ),
    .B(\i57/n426 ),
    .C(\i57/n461 ),
    .Y(\i57/n474 ));
 OAI211xp5_ASAP7_75t_SL \i57/i210  (.A1(\i57/n73 ),
    .A2(\i57/n186 ),
    .B(\i57/n96 ),
    .C(\i57/n142 ),
    .Y(\i57/n281 ));
 NAND4xp25_ASAP7_75t_SL \i57/i211  (.A(\i57/n14 ),
    .B(\i57/n158 ),
    .C(\i57/n551 ),
    .D(\i57/n168 ),
    .Y(\i57/n280 ));
 OAI22xp5_ASAP7_75t_SL \i57/i212  (.A1(\i57/n84 ),
    .A2(\i57/n160 ),
    .B1(\i57/n8 ),
    .B2(\i57/n120 ),
    .Y(\i57/n279 ));
 OAI22xp5_ASAP7_75t_SL \i57/i213  (.A1(\i57/n3 ),
    .A2(\i57/n500 ),
    .B1(\i57/n78 ),
    .B2(\i57/n42 ),
    .Y(\i57/n278 ));
 AOI211x1_ASAP7_75t_SL \i57/i214  (.A1(\i57/n171 ),
    .A2(\i57/n93 ),
    .B(\i57/n190 ),
    .C(\i57/n188 ),
    .Y(\i57/n277 ));
 NAND4xp25_ASAP7_75t_SL \i57/i215  (.A(\i57/n178 ),
    .B(\i57/n194 ),
    .C(\i57/n499 ),
    .D(\i57/n132 ),
    .Y(\i57/n276 ));
 OAI22xp5_ASAP7_75t_SL \i57/i216  (.A1(\i57/n68 ),
    .A2(\i57/n104 ),
    .B1(\i57/n86 ),
    .B2(\i57/n8 ),
    .Y(\i57/n275 ));
 AOI222xp33_ASAP7_75t_SL \i57/i217  (.A1(\i57/n59 ),
    .A2(\i57/n103 ),
    .B1(\i57/n526 ),
    .B2(\i57/n83 ),
    .C1(\i57/n72 ),
    .C2(\i57/n43 ),
    .Y(\i57/n274 ));
 OAI221xp5_ASAP7_75t_R \i57/i218  (.A1(\i57/n498 ),
    .A2(\i57/n82 ),
    .B1(\i57/n75 ),
    .B2(\i57/n92 ),
    .C(\i57/n161 ),
    .Y(\i57/n273 ));
 OAI221xp5_ASAP7_75t_SL \i57/i219  (.A1(\i57/n68 ),
    .A2(\i57/n84 ),
    .B1(\i57/n82 ),
    .B2(\i57/n48 ),
    .C(\i57/n151 ),
    .Y(\i57/n272 ));
 AND4x1_ASAP7_75t_SL \i57/i22  (.A(\i57/n453 ),
    .B(\i57/n458 ),
    .C(\i57/n442 ),
    .D(\i57/n428 ),
    .Y(\i57/n473 ));
 OAI222xp33_ASAP7_75t_SL \i57/i220  (.A1(\i57/n73 ),
    .A2(\i57/n78 ),
    .B1(\i57/n44 ),
    .B2(\i57/n89 ),
    .C1(\i57/n42 ),
    .C2(\i57/n92 ),
    .Y(\i57/n271 ));
 AOI222xp33_ASAP7_75t_SL \i57/i221  (.A1(\i57/n6 ),
    .A2(\i57/n87 ),
    .B1(\i57/n63 ),
    .B2(\i57/n76 ),
    .C1(\i57/n49 ),
    .C2(\i57/n53 ),
    .Y(\i57/n270 ));
 OAI221xp5_ASAP7_75t_SL \i57/i222  (.A1(\i57/n12 ),
    .A2(\i57/n42 ),
    .B1(\i57/n3 ),
    .B2(\i57/n58 ),
    .C(\i57/n502 ),
    .Y(\i57/n269 ));
 OAI211xp5_ASAP7_75t_SL \i57/i223  (.A1(\i57/n58 ),
    .A2(\i57/n141 ),
    .B(\i57/n519 ),
    .C(\i57/n100 ),
    .Y(\i57/n268 ));
 AOI221xp5_ASAP7_75t_SL \i57/i224  (.A1(\i57/n203 ),
    .A2(\i57/n62 ),
    .B1(\i57/n91 ),
    .B2(\i57/n526 ),
    .C(\i57/n131 ),
    .Y(\i57/n267 ));
 AOI22xp33_ASAP7_75t_SL \i57/i225  (.A1(\i57/n51 ),
    .A2(\i57/n203 ),
    .B1(\i57/n76 ),
    .B2(\i57/n6 ),
    .Y(\i57/n266 ));
 AOI221xp5_ASAP7_75t_SL \i57/i226  (.A1(\i57/n172 ),
    .A2(\i57/n79 ),
    .B1(\i57/n65 ),
    .B2(\i57/n67 ),
    .C(\i57/n98 ),
    .Y(\i57/n265 ));
 OAI22xp5_ASAP7_75t_SL \i57/i227  (.A1(\i57/n89 ),
    .A2(\i57/n515 ),
    .B1(\i57/n86 ),
    .B2(\i57/n66 ),
    .Y(\i57/n308 ));
 OAI221xp5_ASAP7_75t_SL \i57/i228  (.A1(\i57/n68 ),
    .A2(\i57/n75 ),
    .B1(\i57/n71 ),
    .B2(\i57/n90 ),
    .C(\i57/n155 ),
    .Y(\i57/n307 ));
 OAI221xp5_ASAP7_75t_SL \i57/i229  (.A1(\i57/n50 ),
    .A2(\i57/n46 ),
    .B1(\i57/n84 ),
    .B2(\i57/n2 ),
    .C(\i57/n108 ),
    .Y(\i57/n305 ));
 NAND3xp33_ASAP7_75t_SL \i57/i23  (.A(\i57/n413 ),
    .B(\i57/n387 ),
    .C(\i57/n410 ),
    .Y(\i57/n471 ));
 OAI21xp5_ASAP7_75t_L \i57/i230  (.A1(\i57/n189 ),
    .A2(\i57/n2 ),
    .B(\i57/n114 ),
    .Y(\i57/n302 ));
 AOI221x1_ASAP7_75t_SL \i57/i231  (.A1(\i57/n7 ),
    .A2(\i57/n6 ),
    .B1(\i57/n77 ),
    .B2(\i57/n167 ),
    .C(\i57/n159 ),
    .Y(\i57/n300 ));
 OAI221xp5_ASAP7_75t_SL \i57/i232  (.A1(\i57/n516 ),
    .A2(\i57/n64 ),
    .B1(\i57/n86 ),
    .B2(\i57/n48 ),
    .C(\i57/n182 ),
    .Y(\i57/n298 ));
 AOI22xp5_ASAP7_75t_SL \i57/i233  (.A1(\i57/n77 ),
    .A2(\i57/n172 ),
    .B1(\i57/n53 ),
    .B2(\i57/n79 ),
    .Y(\i57/n297 ));
 INVxp67_ASAP7_75t_SL \i57/i234  (.A(\i57/n261 ),
    .Y(\i57/n262 ));
 INVxp67_ASAP7_75t_SL \i57/i235  (.A(\i57/n511 ),
    .Y(\i57/n259 ));
 INVxp67_ASAP7_75t_SL \i57/i236  (.A(\i57/n257 ),
    .Y(\i57/n258 ));
 INVx1_ASAP7_75t_SL \i57/i237  (.A(\i57/n253 ),
    .Y(\i57/n254 ));
 INVxp67_ASAP7_75t_SL \i57/i238  (.A(\i57/n251 ),
    .Y(\i57/n252 ));
 INVxp67_ASAP7_75t_SL \i57/i239  (.A(\i57/n512 ),
    .Y(\i57/n248 ));
 NOR2xp33_ASAP7_75t_SL \i57/i24  (.A(\i57/n445 ),
    .B(\i57/n443 ),
    .Y(\i57/n470 ));
 NOR2xp33_ASAP7_75t_SL \i57/i240  (.A(\i57/n192 ),
    .B(\i57/n176 ),
    .Y(\i57/n247 ));
 AOI22xp5_ASAP7_75t_SL \i57/i241  (.A1(\i57/n51 ),
    .A2(\i57/n6 ),
    .B1(\i57/n91 ),
    .B2(\i57/n59 ),
    .Y(\i57/n246 ));
 OAI21xp5_ASAP7_75t_SL \i57/i242  (.A1(\i57/n64 ),
    .A2(\i57/n46 ),
    .B(\i57/n142 ),
    .Y(\i57/n245 ));
 AOI21xp33_ASAP7_75t_SL \i57/i243  (.A1(\i57/n70 ),
    .A2(\i57/n2 ),
    .B(\i57/n173 ),
    .Y(\i57/n244 ));
 OAI21xp5_ASAP7_75t_SL \i57/i244  (.A1(\i57/n3 ),
    .A2(\i57/n66 ),
    .B(\i57/n183 ),
    .Y(\i57/n264 ));
 NAND2xp5_ASAP7_75t_L \i57/i245  (.A(\i57/n143 ),
    .B(\i57/n153 ),
    .Y(\i57/n243 ));
 OAI21xp33_ASAP7_75t_SL \i57/i246  (.A1(\i57/n61 ),
    .A2(\i57/n66 ),
    .B(\i57/n197 ),
    .Y(\i57/n242 ));
 AOI21xp5_ASAP7_75t_SL \i57/i247  (.A1(\i57/n44 ),
    .A2(\i57/n78 ),
    .B(\i57/n84 ),
    .Y(\i57/n263 ));
 AOI21xp33_ASAP7_75t_SL \i57/i248  (.A1(\i57/n78 ),
    .A2(\i57/n488 ),
    .B(\i57/n173 ),
    .Y(\i57/n241 ));
 AOI22xp5_ASAP7_75t_SL \i57/i249  (.A1(\i57/n54 ),
    .A2(\i57/n87 ),
    .B1(\i57/n83 ),
    .B2(\i57/n79 ),
    .Y(\i57/n240 ));
 NAND2xp33_ASAP7_75t_SL \i57/i25  (.A(\i57/n447 ),
    .B(\i57/n437 ),
    .Y(\i57/n469 ));
 OAI21xp33_ASAP7_75t_SL \i57/i250  (.A1(\i57/n60 ),
    .A2(\i57/n66 ),
    .B(\i57/n520 ),
    .Y(\i57/n239 ));
 NOR2xp33_ASAP7_75t_SL \i57/i251  (.A(\i57/n148 ),
    .B(\i57/n179 ),
    .Y(\i57/n238 ));
 OAI22xp5_ASAP7_75t_SL \i57/i252  (.A1(\i57/n90 ),
    .A2(\i57/n2 ),
    .B1(\i57/n80 ),
    .B2(\i57/n44 ),
    .Y(\i57/n237 ));
 OAI21xp5_ASAP7_75t_SL \i57/i253  (.A1(\i57/n55 ),
    .A2(\i57/n52 ),
    .B(\i57/n196 ),
    .Y(\i57/n236 ));
 OAI21xp5_ASAP7_75t_SL \i57/i254  (.A1(\i57/n55 ),
    .A2(\i57/n60 ),
    .B(\i57/n11 ),
    .Y(\i57/n261 ));
 OAI21xp5_ASAP7_75t_SL \i57/i255  (.A1(\i57/n86 ),
    .A2(\i57/n68 ),
    .B(\i57/n200 ),
    .Y(\i57/n260 ));
 OAI22xp5_ASAP7_75t_SL \i57/i256  (.A1(\i57/n70 ),
    .A2(\i57/n61 ),
    .B1(\i57/n82 ),
    .B2(\i57/n68 ),
    .Y(\i57/n257 ));
 AO22x1_ASAP7_75t_SL \i57/i257  (.A1(\i57/n88 ),
    .A2(\i57/n6 ),
    .B1(\i57/n51 ),
    .B2(\i57/n63 ),
    .Y(\i57/n256 ));
 AOI22xp5_ASAP7_75t_SL \i57/i258  (.A1(\i57/n77 ),
    .A2(\i57/n62 ),
    .B1(\i57/n76 ),
    .B2(\i57/n79 ),
    .Y(\i57/n255 ));
 OAI22xp5_ASAP7_75t_SL \i57/i259  (.A1(\i57/n57 ),
    .A2(\i57/n2 ),
    .B1(\i57/n73 ),
    .B2(\i57/n8 ),
    .Y(\i57/n235 ));
 NOR2xp33_ASAP7_75t_SL \i57/i26  (.A(\i57/n427 ),
    .B(\i57/n450 ),
    .Y(\i57/n468 ));
 OAI21xp5_ASAP7_75t_SL \i57/i260  (.A1(\i57/n55 ),
    .A2(\i57/n42 ),
    .B(\i57/n15 ),
    .Y(\i57/n253 ));
 NAND2xp5_ASAP7_75t_SL \i57/i261  (.A(\i57/n47 ),
    .B(\i57/n10 ),
    .Y(\i57/n251 ));
 OAI21xp5_ASAP7_75t_SL \i57/i262  (.A1(\i57/n77 ),
    .A2(\i57/n69 ),
    .B(\i57/n7 ),
    .Y(\i57/n250 ));
 NAND2xp5_ASAP7_75t_SL \i57/i263  (.A(\i57/n93 ),
    .B(\i57/n172 ),
    .Y(\i57/n249 ));
 INVxp67_ASAP7_75t_SL \i57/i264  (.A(\i57/n233 ),
    .Y(\i57/n234 ));
 INVxp67_ASAP7_75t_SL \i57/i265  (.A(\i57/n227 ),
    .Y(\i57/n228 ));
 INVxp67_ASAP7_75t_SL \i57/i266  (.A(\i57/n225 ),
    .Y(\i57/n226 ));
 INVx1_ASAP7_75t_SL \i57/i267  (.A(\i57/n220 ),
    .Y(\i57/n221 ));
 AOI22xp33_ASAP7_75t_SL \i57/i268  (.A1(\i57/n43 ),
    .A2(\i57/n6 ),
    .B1(\i57/n54 ),
    .B2(\i57/n56 ),
    .Y(\i57/n217 ));
 OAI21xp5_ASAP7_75t_SL \i57/i269  (.A1(\i57/n47 ),
    .A2(\i57/n45 ),
    .B(\i57/n53 ),
    .Y(\i57/n216 ));
 NOR2xp33_ASAP7_75t_SL \i57/i27  (.A(\i57/n457 ),
    .B(\i57/n452 ),
    .Y(\i57/n467 ));
 AOI21xp33_ASAP7_75t_SL \i57/i270  (.A1(\i57/n66 ),
    .A2(\i57/n78 ),
    .B(\i57/n42 ),
    .Y(\i57/n215 ));
 AOI22xp5_ASAP7_75t_SL \i57/i271  (.A1(\i57/n59 ),
    .A2(\i57/n62 ),
    .B1(\i57/n79 ),
    .B2(\i57/n88 ),
    .Y(\i57/n214 ));
 AOI22xp5_ASAP7_75t_SL \i57/i272  (.A1(\i57/n93 ),
    .A2(\i57/n62 ),
    .B1(\i57/n87 ),
    .B2(\i57/n47 ),
    .Y(\i57/n233 ));
 OAI22xp5_ASAP7_75t_SL \i57/i273  (.A1(\i57/n82 ),
    .A2(\i57/n58 ),
    .B1(\i57/n55 ),
    .B2(\i57/n84 ),
    .Y(\i57/n213 ));
 OAI21xp5_ASAP7_75t_SL \i57/i274  (.A1(\i57/n90 ),
    .A2(\i57/n44 ),
    .B(\i57/n122 ),
    .Y(\i57/n212 ));
 OAI22xp5_ASAP7_75t_SL \i57/i275  (.A1(\i57/n89 ),
    .A2(\i57/n66 ),
    .B1(\i57/n73 ),
    .B2(\i57/n44 ),
    .Y(\i57/n211 ));
 AOI22xp5_ASAP7_75t_SL \i57/i276  (.A1(\i57/n7 ),
    .A2(\i57/n47 ),
    .B1(\i57/n65 ),
    .B2(\i57/n69 ),
    .Y(\i57/n210 ));
 OAI22xp5_ASAP7_75t_SL \i57/i277  (.A1(\i57/n75 ),
    .A2(\i57/n66 ),
    .B1(\i57/n42 ),
    .B2(\i57/n70 ),
    .Y(\i57/n232 ));
 NAND2xp5_ASAP7_75t_SL \i57/i278  (.A(\i57/n205 ),
    .B(\i57/n13 ),
    .Y(\i57/n209 ));
 NAND2xp5_ASAP7_75t_SL \i57/i279  (.A(\i57/n517 ),
    .B(\i57/n147 ),
    .Y(\i57/n208 ));
 AND2x2_ASAP7_75t_SL \i57/i28  (.A(\i57/n418 ),
    .B(\i57/n449 ),
    .Y(\i57/n472 ));
 OAI22xp5_ASAP7_75t_SL \i57/i280  (.A1(\i57/n55 ),
    .A2(\i57/n90 ),
    .B1(\i57/n73 ),
    .B2(\i57/n71 ),
    .Y(\i57/n231 ));
 OAI22xp5_ASAP7_75t_SL \i57/i281  (.A1(\i57/n50 ),
    .A2(\i57/n44 ),
    .B1(\i57/n488 ),
    .B2(\i57/n89 ),
    .Y(\i57/n230 ));
 OAI22xp33_ASAP7_75t_SL \i57/i282  (.A1(\i57/n84 ),
    .A2(\i57/n488 ),
    .B1(\i57/n530 ),
    .B2(\i57/n73 ),
    .Y(\i57/n207 ));
 OAI22xp5_ASAP7_75t_SL \i57/i283  (.A1(\i57/n66 ),
    .A2(\i57/n73 ),
    .B1(\i57/n46 ),
    .B2(\i57/n42 ),
    .Y(\i57/n229 ));
 OAI22xp5_ASAP7_75t_SL \i57/i284  (.A1(\i57/n55 ),
    .A2(\i57/n89 ),
    .B1(\i57/n92 ),
    .B2(\i57/n73 ),
    .Y(\i57/n227 ));
 AOI22xp5_ASAP7_75t_SL \i57/i285  (.A1(\i57/n67 ),
    .A2(\i57/n91 ),
    .B1(\i57/n93 ),
    .B2(\i57/n81 ),
    .Y(\i57/n225 ));
 OAI22xp5_ASAP7_75t_SL \i57/i286  (.A1(\i57/n82 ),
    .A2(\i57/n44 ),
    .B1(\i57/n71 ),
    .B2(\i57/n57 ),
    .Y(\i57/n224 ));
 OAI22xp5_ASAP7_75t_SL \i57/i287  (.A1(\i57/n488 ),
    .A2(\i57/n50 ),
    .B1(\i57/n8 ),
    .B2(\i57/n42 ),
    .Y(\i57/n223 ));
 AOI22xp5_ASAP7_75t_SL \i57/i288  (.A1(\i57/n62 ),
    .A2(\i57/n6 ),
    .B1(\i57/n43 ),
    .B2(\i57/n69 ),
    .Y(\i57/n222 ));
 AOI22xp33_ASAP7_75t_SL \i57/i289  (.A1(\i57/n91 ),
    .A2(\i57/n72 ),
    .B1(\i57/n79 ),
    .B2(\i57/n65 ),
    .Y(\i57/n206 ));
 NOR2xp33_ASAP7_75t_SL \i57/i29  (.A(\i57/n456 ),
    .B(\i57/n440 ),
    .Y(\i57/n466 ));
 AO22x1_ASAP7_75t_SL \i57/i290  (.A1(\i57/n53 ),
    .A2(\i57/n67 ),
    .B1(\i57/n79 ),
    .B2(\i57/n91 ),
    .Y(\i57/n220 ));
 AOI22xp5_ASAP7_75t_SL \i57/i291  (.A1(\i57/n45 ),
    .A2(\i57/n62 ),
    .B1(\i57/n81 ),
    .B2(\i57/n79 ),
    .Y(\i57/n219 ));
 AOI22xp5_ASAP7_75t_SL \i57/i292  (.A1(\i57/n526 ),
    .A2(\i57/n85 ),
    .B1(\i57/n74 ),
    .B2(\i57/n59 ),
    .Y(\i57/n218 ));
 INVxp67_ASAP7_75t_SL \i57/i293  (.A(\i57/n13 ),
    .Y(\i57/n202 ));
 INVxp67_ASAP7_75t_SL \i57/i294  (.A(\i57/n198 ),
    .Y(\i57/n199 ));
 INVxp67_ASAP7_75t_SL \i57/i295  (.A(\i57/n194 ),
    .Y(\i57/n195 ));
 INVxp67_ASAP7_75t_SL \i57/i296  (.A(\i57/n192 ),
    .Y(\i57/n193 ));
 INVxp67_ASAP7_75t_SL \i57/i297  (.A(\i57/n190 ),
    .Y(\i57/n191 ));
 INVxp67_ASAP7_75t_SL \i57/i298  (.A(\i57/n495 ),
    .Y(\i57/n184 ));
 INVx1_ASAP7_75t_SL \i57/i299  (.A(\i57/n180 ),
    .Y(\i57/n181 ));
 INVx3_ASAP7_75t_SL \i57/i3  (.A(\i57/n544 ),
    .Y(\i57/n3 ));
 NOR2xp33_ASAP7_75t_SL \i57/i30  (.A(\i57/n439 ),
    .B(\i57/n434 ),
    .Y(\i57/n465 ));
 INVxp67_ASAP7_75t_SL \i57/i300  (.A(\i57/n178 ),
    .Y(\i57/n179 ));
 INVxp67_ASAP7_75t_SL \i57/i301  (.A(\i57/n176 ),
    .Y(\i57/n177 ));
 INVx1_ASAP7_75t_SL \i57/i302  (.A(\i57/n174 ),
    .Y(\i57/n175 ));
 NAND2xp5_ASAP7_75t_L \i57/i303  (.A(\i57/n86 ),
    .B(\i57/n75 ),
    .Y(\i57/n171 ));
 NAND2xp5_ASAP7_75t_SL \i57/i304  (.A(\i57/n63 ),
    .B(\i57/n65 ),
    .Y(\i57/n170 ));
 NAND2xp33_ASAP7_75t_L \i57/i305  (.A(\i57/n90 ),
    .B(\i57/n80 ),
    .Y(\i57/n169 ));
 NAND2xp5_ASAP7_75t_SL \i57/i306  (.A(\i57/n72 ),
    .B(\i57/n65 ),
    .Y(\i57/n168 ));
 NAND2xp5_ASAP7_75t_SL \i57/i307  (.A(\i57/n52 ),
    .B(\i57/n3 ),
    .Y(\i57/n167 ));
 NAND2xp5_ASAP7_75t_SL \i57/i308  (.A(\i57/n61 ),
    .B(\i57/n3 ),
    .Y(\i57/n166 ));
 NOR2xp33_ASAP7_75t_SL \i57/i309  (.A(\i57/n81 ),
    .B(\i57/n85 ),
    .Y(\i57/n165 ));
 NOR2xp33_ASAP7_75t_SL \i57/i31  (.A(\i57/n433 ),
    .B(\i57/n451 ),
    .Y(\i57/n464 ));
 NOR2xp33_ASAP7_75t_SL \i57/i310  (.A(\i57/n85 ),
    .B(\i57/n65 ),
    .Y(\i57/n164 ));
 NAND2xp5_ASAP7_75t_SL \i57/i311  (.A(\i57/n49 ),
    .B(\i57/n91 ),
    .Y(\i57/n205 ));
 NAND2xp5_ASAP7_75t_SL \i57/i312  (.A(\i57/n59 ),
    .B(\i57/n88 ),
    .Y(\i57/n163 ));
 NOR2xp67_ASAP7_75t_L \i57/i313  (.A(\i57/n89 ),
    .B(\i57/n8 ),
    .Y(\i57/n162 ));
 NAND2xp5_ASAP7_75t_SL \i57/i314  (.A(\i57/n63 ),
    .B(\i57/n53 ),
    .Y(\i57/n161 ));
 NOR2xp33_ASAP7_75t_SL \i57/i315  (.A(\i57/n54 ),
    .B(\i57/n45 ),
    .Y(\i57/n160 ));
 NOR2xp67_ASAP7_75t_SL \i57/i316  (.A(\i57/n82 ),
    .B(\i57/n71 ),
    .Y(\i57/n159 ));
 NAND2xp5_ASAP7_75t_SL \i57/i317  (.A(\i57/n85 ),
    .B(\i57/n49 ),
    .Y(\i57/n158 ));
 NOR2xp33_ASAP7_75t_SL \i57/i318  (.A(\i57/n67 ),
    .B(\i57/n72 ),
    .Y(\i57/n157 ));
 NOR2xp33_ASAP7_75t_SL \i57/i319  (.A(\i57/n47 ),
    .B(\i57/n67 ),
    .Y(\i57/n156 ));
 AND4x1_ASAP7_75t_SL \i57/i32  (.A(\i57/n423 ),
    .B(\i57/n419 ),
    .C(\i57/n379 ),
    .D(\i57/n372 ),
    .Y(\i57/n463 ));
 NAND2xp5_ASAP7_75t_SL \i57/i320  (.A(\i57/n79 ),
    .B(\i57/n65 ),
    .Y(\i57/n155 ));
 NOR2xp33_ASAP7_75t_SL \i57/i321  (.A(\i57/n77 ),
    .B(\i57/n72 ),
    .Y(\i57/n154 ));
 NAND2xp5_ASAP7_75t_SL \i57/i322  (.A(\i57/n65 ),
    .B(\i57/n45 ),
    .Y(\i57/n204 ));
 NAND2xp5_ASAP7_75t_SL \i57/i323  (.A(\i57/n79 ),
    .B(\i57/n62 ),
    .Y(\i57/n153 ));
 NAND2xp5_ASAP7_75t_SL \i57/i324  (.A(\i57/n74 ),
    .B(\i57/n69 ),
    .Y(\i57/n152 ));
 NAND2xp5_ASAP7_75t_SL \i57/i325  (.A(\i57/n54 ),
    .B(\i57/n74 ),
    .Y(\i57/n151 ));
 NOR2xp33_ASAP7_75t_SL \i57/i326  (.A(\i57/n73 ),
    .B(\i57/n8 ),
    .Y(\i57/n150 ));
 NAND2xp33_ASAP7_75t_SL \i57/i327  (.A(\i57/n46 ),
    .B(\i57/n78 ),
    .Y(\i57/n203 ));
 NAND2xp5_ASAP7_75t_SL \i57/i328  (.A(\i57/n56 ),
    .B(\i57/n67 ),
    .Y(\i57/n15 ));
 NAND2xp5_ASAP7_75t_SL \i57/i329  (.A(\i57/n79 ),
    .B(\i57/n7 ),
    .Y(\i57/n14 ));
 NOR3xp33_ASAP7_75t_SL \i57/i33  (.A(\i57/n416 ),
    .B(\i57/n352 ),
    .C(\i57/n404 ),
    .Y(\i57/n462 ));
 NOR2xp33_ASAP7_75t_SL \i57/i330  (.A(\i57/n78 ),
    .B(\i57/n75 ),
    .Y(\i57/n149 ));
 NAND2xp5_ASAP7_75t_SL \i57/i331  (.A(\i57/n83 ),
    .B(\i57/n67 ),
    .Y(\i57/n13 ));
 NAND2xp5_ASAP7_75t_SL \i57/i332  (.A(\i57/n93 ),
    .B(\i57/n83 ),
    .Y(\i57/n201 ));
 NAND2xp5_ASAP7_75t_SL \i57/i333  (.A(\i57/n93 ),
    .B(\i57/n56 ),
    .Y(\i57/n200 ));
 NAND2xp5_ASAP7_75t_L \i57/i334  (.A(\i57/n85 ),
    .B(\i57/n93 ),
    .Y(\i57/n198 ));
 NAND2xp5_ASAP7_75t_SL \i57/i335  (.A(\i57/n77 ),
    .B(\i57/n83 ),
    .Y(\i57/n197 ));
 NAND2xp5_ASAP7_75t_SL \i57/i336  (.A(\i57/n81 ),
    .B(\i57/n77 ),
    .Y(\i57/n196 ));
 NAND2xp5_ASAP7_75t_SL \i57/i337  (.A(\i57/n526 ),
    .B(\i57/n65 ),
    .Y(\i57/n194 ));
 NAND2xp33_ASAP7_75t_SL \i57/i338  (.A(\i57/n50 ),
    .B(\i57/n89 ),
    .Y(\i57/n192 ));
 AND2x2_ASAP7_75t_SL \i57/i339  (.A(\i57/n91 ),
    .B(\i57/n77 ),
    .Y(\i57/n190 ));
 NAND2xp33_ASAP7_75t_SL \i57/i34  (.A(\i57/n18 ),
    .B(\i57/n435 ),
    .Y(\i57/n461 ));
 NOR2xp33_ASAP7_75t_SL \i57/i340  (.A(\i57/n74 ),
    .B(\i57/n53 ),
    .Y(\i57/n189 ));
 AND2x2_ASAP7_75t_SL \i57/i341  (.A(\i57/n88 ),
    .B(\i57/n72 ),
    .Y(\i57/n188 ));
 NAND2xp5_ASAP7_75t_SL \i57/i342  (.A(\i57/n74 ),
    .B(\i57/n49 ),
    .Y(\i57/n187 ));
 NOR2xp33_ASAP7_75t_L \i57/i343  (.A(\i57/n47 ),
    .B(\i57/n63 ),
    .Y(\i57/n186 ));
 NAND2xp5_ASAP7_75t_SL \i57/i344  (.A(\i57/n49 ),
    .B(\i57/n65 ),
    .Y(\i57/n185 ));
 NAND2xp5_ASAP7_75t_SL \i57/i345  (.A(\i57/n63 ),
    .B(\i57/n43 ),
    .Y(\i57/n183 ));
 NAND2xp5_ASAP7_75t_SL \i57/i346  (.A(\i57/n63 ),
    .B(\i57/n85 ),
    .Y(\i57/n182 ));
 NOR2xp33_ASAP7_75t_SL \i57/i347  (.A(\i57/n50 ),
    .B(\i57/n530 ),
    .Y(\i57/n148 ));
 NOR2xp33_ASAP7_75t_L \i57/i348  (.A(\i57/n43 ),
    .B(\i57/n74 ),
    .Y(\i57/n180 ));
 NAND2xp5_ASAP7_75t_SL \i57/i349  (.A(\i57/n93 ),
    .B(\i57/n7 ),
    .Y(\i57/n178 ));
 INVxp67_ASAP7_75t_SL \i57/i35  (.A(\i57/n459 ),
    .Y(\i57/n460 ));
 NAND2xp5_ASAP7_75t_L \i57/i350  (.A(\i57/n3 ),
    .B(\i57/n80 ),
    .Y(\i57/n176 ));
 NOR2xp33_ASAP7_75t_L \i57/i351  (.A(\i57/n87 ),
    .B(\i57/n81 ),
    .Y(\i57/n174 ));
 NOR2xp33_ASAP7_75t_L \i57/i352  (.A(\i57/n87 ),
    .B(\i57/n74 ),
    .Y(\i57/n173 ));
 NAND2xp5_ASAP7_75t_SL \i57/i353  (.A(\i57/n50 ),
    .B(\i57/n64 ),
    .Y(\i57/n172 ));
 INVxp67_ASAP7_75t_SL \i57/i354  (.A(\i57/n143 ),
    .Y(\i57/n144 ));
 INVxp67_ASAP7_75t_SL \i57/i355  (.A(\i57/n519 ),
    .Y(\i57/n138 ));
 INVxp67_ASAP7_75t_SL \i57/i356  (.A(\i57/n133 ),
    .Y(\i57/n134 ));
 INVxp67_ASAP7_75t_SL \i57/i357  (.A(\i57/n130 ),
    .Y(\i57/n131 ));
 INVxp67_ASAP7_75t_SL \i57/i358  (.A(\i57/n9 ),
    .Y(\i57/n127 ));
 NOR2xp33_ASAP7_75t_SL \i57/i359  (.A(\i57/n47 ),
    .B(\i57/n59 ),
    .Y(\i57/n126 ));
 INVxp67_ASAP7_75t_SL \i57/i36  (.A(\i57/n457 ),
    .Y(\i57/n458 ));
 NOR2xp33_ASAP7_75t_SL \i57/i360  (.A(\i57/n86 ),
    .B(\i57/n508 ),
    .Y(\i57/n125 ));
 NAND2xp33_ASAP7_75t_SL \i57/i361  (.A(\i57/n57 ),
    .B(\i57/n80 ),
    .Y(\i57/n124 ));
 NOR2xp33_ASAP7_75t_SL \i57/i362  (.A(\i57/n83 ),
    .B(\i57/n7 ),
    .Y(\i57/n123 ));
 NAND2xp5_ASAP7_75t_SL \i57/i363  (.A(\i57/n47 ),
    .B(\i57/n85 ),
    .Y(\i57/n122 ));
 NAND2xp5_ASAP7_75t_SL \i57/i364  (.A(\i57/n87 ),
    .B(\i57/n45 ),
    .Y(\i57/n121 ));
 NOR2xp33_ASAP7_75t_SL \i57/i365  (.A(\i57/n87 ),
    .B(\i57/n53 ),
    .Y(\i57/n120 ));
 NAND2xp33_ASAP7_75t_L \i57/i366  (.A(\i57/n2 ),
    .B(\i57/n58 ),
    .Y(\i57/n119 ));
 NAND2xp5_ASAP7_75t_SL \i57/i367  (.A(\i57/n76 ),
    .B(\i57/n77 ),
    .Y(\i57/n118 ));
 NAND2xp33_ASAP7_75t_SL \i57/i368  (.A(\i57/n60 ),
    .B(\i57/n57 ),
    .Y(\i57/n117 ));
 NOR2xp33_ASAP7_75t_SL \i57/i369  (.A(\i57/n7 ),
    .B(\i57/n43 ),
    .Y(\i57/n116 ));
 NAND3xp33_ASAP7_75t_SL \i57/i37  (.A(\i57/n412 ),
    .B(\i57/n365 ),
    .C(\i57/n371 ),
    .Y(\i57/n455 ));
 NAND2xp5_ASAP7_75t_SL \i57/i370  (.A(\i57/n77 ),
    .B(\i57/n56 ),
    .Y(\i57/n115 ));
 NAND2xp5_ASAP7_75t_SL \i57/i371  (.A(\i57/n7 ),
    .B(\i57/n59 ),
    .Y(\i57/n114 ));
 NAND2xp33_ASAP7_75t_SL \i57/i372  (.A(\i57/n46 ),
    .B(\i57/n70 ),
    .Y(\i57/n113 ));
 NAND2xp33_ASAP7_75t_SL \i57/i373  (.A(\i57/n75 ),
    .B(\i57/n71 ),
    .Y(\i57/n112 ));
 NOR2xp33_ASAP7_75t_SL \i57/i374  (.A(\i57/n49 ),
    .B(\i57/n526 ),
    .Y(\i57/n111 ));
 NAND2xp33_ASAP7_75t_L \i57/i375  (.A(\i57/n48 ),
    .B(\i57/n55 ),
    .Y(\i57/n110 ));
 NAND2xp5_ASAP7_75t_SL \i57/i376  (.A(\i57/n49 ),
    .B(\i57/n62 ),
    .Y(\i57/n147 ));
 NAND2xp33_ASAP7_75t_SL \i57/i377  (.A(\i57/n508 ),
    .B(\i57/n48 ),
    .Y(\i57/n109 ));
 NAND2xp5_ASAP7_75t_SL \i57/i378  (.A(\i57/n53 ),
    .B(\i57/n72 ),
    .Y(\i57/n108 ));
 NAND2xp5_ASAP7_75t_SL \i57/i379  (.A(\i57/n49 ),
    .B(\i57/n51 ),
    .Y(\i57/n146 ));
 NAND2xp5_ASAP7_75t_L \i57/i38  (.A(\i57/n402 ),
    .B(\i57/n391 ),
    .Y(\i57/n454 ));
 NOR2xp33_ASAP7_75t_SL \i57/i380  (.A(\i57/n50 ),
    .B(\i57/n70 ),
    .Y(\i57/n107 ));
 NOR2xp33_ASAP7_75t_SL \i57/i381  (.A(\i57/n59 ),
    .B(\i57/n45 ),
    .Y(\i57/n106 ));
 NAND2xp33_ASAP7_75t_SL \i57/i382  (.A(\i57/n508 ),
    .B(\i57/n68 ),
    .Y(\i57/n105 ));
 NOR2xp33_ASAP7_75t_SL \i57/i383  (.A(\i57/n56 ),
    .B(\i57/n43 ),
    .Y(\i57/n104 ));
 NAND2xp5_ASAP7_75t_L \i57/i384  (.A(\i57/n57 ),
    .B(\i57/n75 ),
    .Y(\i57/n103 ));
 NAND2xp5_ASAP7_75t_SL \i57/i385  (.A(\i57/n81 ),
    .B(\i57/n69 ),
    .Y(\i57/n102 ));
 NOR2xp33_ASAP7_75t_SL \i57/i386  (.A(\i57/n77 ),
    .B(\i57/n526 ),
    .Y(\i57/n12 ));
 NAND2xp5_ASAP7_75t_SL \i57/i387  (.A(\i57/n53 ),
    .B(\i57/n526 ),
    .Y(\i57/n145 ));
 NOR2xp33_ASAP7_75t_SL \i57/i388  (.A(\i57/n57 ),
    .B(\i57/n70 ),
    .Y(\i57/n101 ));
 NAND2xp5_ASAP7_75t_SL \i57/i389  (.A(\i57/n51 ),
    .B(\i57/n6 ),
    .Y(\i57/n100 ));
 NOR2xp33_ASAP7_75t_SL \i57/i39  (.A(\i57/n420 ),
    .B(\i57/n350 ),
    .Y(\i57/n453 ));
 NOR2xp33_ASAP7_75t_SL \i57/i390  (.A(\i57/n80 ),
    .B(\i57/n44 ),
    .Y(\i57/n99 ));
 NAND2xp5_ASAP7_75t_SL \i57/i391  (.A(\i57/n83 ),
    .B(\i57/n47 ),
    .Y(\i57/n143 ));
 NOR2xp33_ASAP7_75t_SL \i57/i392  (.A(\i57/n82 ),
    .B(\i57/n68 ),
    .Y(\i57/n98 ));
 NAND2xp5_ASAP7_75t_SL \i57/i393  (.A(\i57/n54 ),
    .B(\i57/n81 ),
    .Y(\i57/n142 ));
 NAND2xp5_ASAP7_75t_SL \i57/i394  (.A(\i57/n62 ),
    .B(\i57/n72 ),
    .Y(\i57/n11 ));
 NAND2x1p5_ASAP7_75t_SL \i57/i395  (.A(\i57/n80 ),
    .B(\i57/n75 ),
    .Y(\i57/n10 ));
 NOR2xp33_ASAP7_75t_L \i57/i396  (.A(\i57/n7 ),
    .B(\i57/n76 ),
    .Y(\i57/n141 ));
 NAND2xp5_ASAP7_75t_SL \i57/i397  (.A(\i57/n76 ),
    .B(\i57/n45 ),
    .Y(\i57/n140 ));
 NAND2xp5_ASAP7_75t_SL \i57/i398  (.A(\i57/n56 ),
    .B(\i57/n45 ),
    .Y(\i57/n139 ));
 NOR2xp33_ASAP7_75t_SL \i57/i399  (.A(\i57/n55 ),
    .B(\i57/n61 ),
    .Y(\i57/n97 ));
 AND3x2_ASAP7_75t_SL \i57/i4  (.A(\i57/n470 ),
    .B(\i57/n483 ),
    .C(\i57/n556 ),
    .Y(n6[6]));
 NAND2xp33_ASAP7_75t_SL \i57/i40  (.A(\i57/n396 ),
    .B(\i57/n414 ),
    .Y(\i57/n452 ));
 NAND2xp5_ASAP7_75t_SL \i57/i400  (.A(\i57/n54 ),
    .B(\i57/n87 ),
    .Y(\i57/n96 ));
 NAND2xp5_ASAP7_75t_SL \i57/i401  (.A(\i57/n43 ),
    .B(\i57/n6 ),
    .Y(\i57/n95 ));
 NAND2xp5_ASAP7_75t_SL \i57/i402  (.A(\i57/n51 ),
    .B(\i57/n69 ),
    .Y(\i57/n137 ));
 NOR2xp33_ASAP7_75t_SL \i57/i403  (.A(\i57/n508 ),
    .B(\i57/n52 ),
    .Y(\i57/n94 ));
 NAND2xp5_ASAP7_75t_SL \i57/i404  (.A(\i57/n43 ),
    .B(\i57/n59 ),
    .Y(\i57/n136 ));
 NAND2xp5_ASAP7_75t_SL \i57/i405  (.A(\i57/n53 ),
    .B(\i57/n59 ),
    .Y(\i57/n135 ));
 AND2x2_ASAP7_75t_SL \i57/i406  (.A(\i57/n56 ),
    .B(\i57/n47 ),
    .Y(\i57/n133 ));
 NAND4xp25_ASAP7_75t_SL \i57/i407  (.A(\i57/n32 ),
    .B(\i57/n37 ),
    .C(\i57/n543 ),
    .D(\i57/n27 ),
    .Y(\i57/n132 ));
 NAND2xp5_ASAP7_75t_SL \i57/i408  (.A(\i57/n49 ),
    .B(\i57/n43 ),
    .Y(\i57/n130 ));
 AND2x2_ASAP7_75t_SL \i57/i409  (.A(\i57/n53 ),
    .B(\i57/n47 ),
    .Y(\i57/n129 ));
 NAND3xp33_ASAP7_75t_SL \i57/i41  (.A(\i57/n425 ),
    .B(\i57/n267 ),
    .C(\i57/n297 ),
    .Y(\i57/n451 ));
 AND2x2_ASAP7_75t_SL \i57/i410  (.A(\i57/n51 ),
    .B(\i57/n59 ),
    .Y(\i57/n128 ));
 NAND2xp5_ASAP7_75t_SL \i57/i411  (.A(\i57/n85 ),
    .B(\i57/n59 ),
    .Y(\i57/n9 ));
 INVx2_ASAP7_75t_SL \i57/i412  (.A(\i57/n93 ),
    .Y(\i57/n92 ));
 INVx2_ASAP7_75t_SL \i57/i413  (.A(\i57/n91 ),
    .Y(\i57/n90 ));
 INVx3_ASAP7_75t_SL \i57/i414  (.A(\i57/n89 ),
    .Y(\i57/n88 ));
 INVx4_ASAP7_75t_SL \i57/i415  (.A(\i57/n87 ),
    .Y(\i57/n86 ));
 INVx3_ASAP7_75t_SL \i57/i416  (.A(\i57/n85 ),
    .Y(\i57/n84 ));
 INVx3_ASAP7_75t_SL \i57/i417  (.A(\i57/n83 ),
    .Y(\i57/n82 ));
 INVx3_ASAP7_75t_SL \i57/i418  (.A(\i57/n81 ),
    .Y(\i57/n80 ));
 INVx2_ASAP7_75t_SL \i57/i419  (.A(\i57/n79 ),
    .Y(\i57/n78 ));
 NAND2xp33_ASAP7_75t_SL \i57/i42  (.A(\i57/n407 ),
    .B(\i57/n411 ),
    .Y(\i57/n450 ));
 INVx3_ASAP7_75t_SL \i57/i420  (.A(\i57/n76 ),
    .Y(\i57/n75 ));
 INVx2_ASAP7_75t_SL \i57/i421  (.A(\i57/n74 ),
    .Y(\i57/n73 ));
 INVx2_ASAP7_75t_SL \i57/i422  (.A(\i57/n72 ),
    .Y(\i57/n71 ));
 INVx2_ASAP7_75t_SL \i57/i423  (.A(\i57/n526 ),
    .Y(\i57/n70 ));
 INVx3_ASAP7_75t_SL \i57/i424  (.A(\i57/n69 ),
    .Y(\i57/n68 ));
 INVx3_ASAP7_75t_SL \i57/i425  (.A(\i57/n67 ),
    .Y(\i57/n66 ));
 AND2x4_ASAP7_75t_SL \i57/i426  (.A(\i57/n484 ),
    .B(\i57/n31 ),
    .Y(\i57/n93 ));
 AND2x4_ASAP7_75t_SL \i57/i427  (.A(\i57/n38 ),
    .B(\i57/n543 ),
    .Y(\i57/n91 ));
 OR2x6_ASAP7_75t_SL \i57/i428  (.A(\i57/n26 ),
    .B(\i57/n39 ),
    .Y(\i57/n89 ));
 AND2x4_ASAP7_75t_SL \i57/i429  (.A(\i57/n40 ),
    .B(\i57/n33 ),
    .Y(\i57/n87 ));
 NOR2xp33_ASAP7_75t_SL \i57/i43  (.A(\i57/n409 ),
    .B(\i57/n408 ),
    .Y(\i57/n449 ));
 AND2x4_ASAP7_75t_SL \i57/i430  (.A(\i57/n41 ),
    .B(\i57/n27 ),
    .Y(\i57/n85 ));
 AND2x4_ASAP7_75t_SL \i57/i431  (.A(\i57/n33 ),
    .B(\i57/n38 ),
    .Y(\i57/n83 ));
 AND2x4_ASAP7_75t_SL \i57/i432  (.A(\i57/n34 ),
    .B(\i57/n27 ),
    .Y(\i57/n81 ));
 AND2x4_ASAP7_75t_SL \i57/i433  (.A(\i57/n36 ),
    .B(\i57/n35 ),
    .Y(\i57/n79 ));
 AND2x2_ASAP7_75t_SL \i57/i434  (.A(\i57/n36 ),
    .B(\i57/n28 ),
    .Y(\i57/n77 ));
 NAND2x1_ASAP7_75t_SL \i57/i435  (.A(\i57/n36 ),
    .B(\i57/n28 ),
    .Y(\i57/n8 ));
 AND2x4_ASAP7_75t_SL \i57/i436  (.A(\i57/n33 ),
    .B(\i57/n542 ),
    .Y(\i57/n76 ));
 AND2x4_ASAP7_75t_SL \i57/i437  (.A(\i57/n33 ),
    .B(\i57/n27 ),
    .Y(\i57/n74 ));
 AND2x4_ASAP7_75t_SL \i57/i438  (.A(\i57/n36 ),
    .B(\i57/n504 ),
    .Y(\i57/n72 ));
 AND2x4_ASAP7_75t_SL \i57/i439  (.A(\i57/n36 ),
    .B(\i57/n37 ),
    .Y(\i57/n69 ));
 NAND4xp25_ASAP7_75t_SL \i57/i44  (.A(\i57/n386 ),
    .B(\i57/n546 ),
    .C(\i57/n248 ),
    .D(\i57/n290 ),
    .Y(\i57/n448 ));
 AND2x4_ASAP7_75t_SL \i57/i440  (.A(\i57/n32 ),
    .B(\i57/n37 ),
    .Y(\i57/n67 ));
 INVx3_ASAP7_75t_SL \i57/i441  (.A(\i57/n65 ),
    .Y(\i57/n64 ));
 INVx2_ASAP7_75t_SL \i57/i442  (.A(\i57/n62 ),
    .Y(\i57/n61 ));
 INVx2_ASAP7_75t_SL \i57/i443  (.A(\i57/n59 ),
    .Y(\i57/n58 ));
 INVx2_ASAP7_75t_SL \i57/i444  (.A(\i57/n55 ),
    .Y(\i57/n54 ));
 INVx2_ASAP7_75t_SL \i57/i445  (.A(\i57/n53 ),
    .Y(\i57/n52 ));
 INVx3_ASAP7_75t_SL \i57/i446  (.A(\i57/n51 ),
    .Y(\i57/n50 ));
 INVx4_ASAP7_75t_SL \i57/i447  (.A(\i57/n49 ),
    .Y(\i57/n48 ));
 INVx2_ASAP7_75t_SL \i57/i448  (.A(\i57/n47 ),
    .Y(\i57/n46 ));
 INVx4_ASAP7_75t_SL \i57/i449  (.A(\i57/n45 ),
    .Y(\i57/n44 ));
 NOR2xp33_ASAP7_75t_SL \i57/i45  (.A(\i57/n424 ),
    .B(\i57/n401 ),
    .Y(\i57/n447 ));
 INVx3_ASAP7_75t_SL \i57/i450  (.A(\i57/n43 ),
    .Y(\i57/n42 ));
 AND2x4_ASAP7_75t_SL \i57/i451  (.A(\i57/n542 ),
    .B(\i57/n41 ),
    .Y(\i57/n65 ));
 AND2x4_ASAP7_75t_SL \i57/i452  (.A(\i57/n24 ),
    .B(\i57/n35 ),
    .Y(\i57/n63 ));
 AND2x4_ASAP7_75t_SL \i57/i453  (.A(\i57/n27 ),
    .B(\i57/n543 ),
    .Y(\i57/n62 ));
 NAND2x1p5_ASAP7_75t_SL \i57/i454  (.A(\i57/n34 ),
    .B(\i57/n542 ),
    .Y(\i57/n60 ));
 AND2x4_ASAP7_75t_SL \i57/i455  (.A(\i57/n32 ),
    .B(\i57/n504 ),
    .Y(\i57/n6 ));
 AND2x4_ASAP7_75t_SL \i57/i456  (.A(\i57/n29 ),
    .B(\i57/n28 ),
    .Y(\i57/n59 ));
 NAND2xp5_ASAP7_75t_SL \i57/i457  (.A(\i57/n41 ),
    .B(\i57/n38 ),
    .Y(\i57/n57 ));
 AND4x1_ASAP7_75t_SL \i57/i458  (.A(n7[6]),
    .B(\i57/n0 ),
    .C(\i57/n5 ),
    .D(n7[4]),
    .Y(\i57/n56 ));
 OR2x6_ASAP7_75t_SL \i57/i459  (.A(\i57/n30 ),
    .B(\i57/n25 ),
    .Y(\i57/n55 ));
 NAND3xp33_ASAP7_75t_SL \i57/i46  (.A(\i57/n368 ),
    .B(\i57/n359 ),
    .C(\i57/n297 ),
    .Y(\i57/n446 ));
 AND2x4_ASAP7_75t_SL \i57/i460  (.A(\i57/n40 ),
    .B(\i57/n41 ),
    .Y(\i57/n53 ));
 AND2x4_ASAP7_75t_SL \i57/i461  (.A(\i57/n38 ),
    .B(\i57/n34 ),
    .Y(\i57/n51 ));
 AND2x4_ASAP7_75t_SL \i57/i462  (.A(\i57/n35 ),
    .B(\i57/n29 ),
    .Y(\i57/n49 ));
 AND2x4_ASAP7_75t_SL \i57/i463  (.A(\i57/n35 ),
    .B(\i57/n32 ),
    .Y(\i57/n47 ));
 AND2x4_ASAP7_75t_SL \i57/i464  (.A(\i57/n37 ),
    .B(\i57/n29 ),
    .Y(\i57/n45 ));
 AND2x4_ASAP7_75t_SL \i57/i465  (.A(\i57/n40 ),
    .B(\i57/n34 ),
    .Y(\i57/n43 ));
 INVx2_ASAP7_75t_SL \i57/i466  (.A(\i57/n40 ),
    .Y(\i57/n39 ));
 AND2x2_ASAP7_75t_SL \i57/i467  (.A(n7[6]),
    .B(\i57/n5 ),
    .Y(\i57/n41 ));
 AND2x2_ASAP7_75t_SL \i57/i468  (.A(n7[5]),
    .B(\i57/n20 ),
    .Y(\i57/n40 ));
 AND2x2_ASAP7_75t_SL \i57/i469  (.A(n7[4]),
    .B(\i57/n0 ),
    .Y(\i57/n38 ));
 NAND3xp33_ASAP7_75t_SL \i57/i47  (.A(\i57/n386 ),
    .B(\i57/n369 ),
    .C(\i57/n356 ),
    .Y(\i57/n445 ));
 AND2x2_ASAP7_75t_SL \i57/i470  (.A(\i57/n23 ),
    .B(\i57/n1 ),
    .Y(\i57/n37 ));
 AND2x2_ASAP7_75t_SL \i57/i471  (.A(n7[2]),
    .B(n7[0]),
    .Y(\i57/n36 ));
 AND2x2_ASAP7_75t_SL \i57/i472  (.A(n7[3]),
    .B(n7[1]),
    .Y(\i57/n35 ));
 AND2x4_ASAP7_75t_SL \i57/i473  (.A(n7[7]),
    .B(\i57/n21 ),
    .Y(\i57/n34 ));
 AND2x2_ASAP7_75t_SL \i57/i474  (.A(n7[7]),
    .B(n7[6]),
    .Y(\i57/n33 ));
 AND2x4_ASAP7_75t_L \i57/i475  (.A(\i57/n22 ),
    .B(\i57/n19 ),
    .Y(\i57/n32 ));
 INVx1_ASAP7_75t_SL \i57/i476  (.A(\i57/n30 ),
    .Y(\i57/n31 ));
 NAND2xp5_ASAP7_75t_SL \i57/i477  (.A(n7[3]),
    .B(\i57/n22 ),
    .Y(\i57/n25 ));
 NOR2xp33_ASAP7_75t_SL \i57/i478  (.A(\i57/n19 ),
    .B(n7[2]),
    .Y(\i57/n24 ));
 OR2x2_ASAP7_75t_SL \i57/i479  (.A(\i57/n19 ),
    .B(n7[1]),
    .Y(\i57/n30 ));
 NOR3xp33_ASAP7_75t_SL \i57/i48  (.A(\i57/n339 ),
    .B(\i57/n512 ),
    .C(\i57/n374 ),
    .Y(\i57/n459 ));
 AND2x2_ASAP7_75t_SL \i57/i480  (.A(n7[2]),
    .B(\i57/n19 ),
    .Y(\i57/n29 ));
 AND2x2_ASAP7_75t_SL \i57/i481  (.A(n7[1]),
    .B(\i57/n23 ),
    .Y(\i57/n28 ));
 AND2x2_ASAP7_75t_SL \i57/i482  (.A(n7[5]),
    .B(n7[4]),
    .Y(\i57/n27 ));
 OR2x2_ASAP7_75t_SL \i57/i483  (.A(n7[7]),
    .B(n7[6]),
    .Y(\i57/n26 ));
 INVx3_ASAP7_75t_SL \i57/i484  (.A(n7[7]),
    .Y(\i57/n5 ));
 INVx2_ASAP7_75t_SL \i57/i485  (.A(n7[3]),
    .Y(\i57/n23 ));
 INVx4_ASAP7_75t_SL \i57/i486  (.A(n7[2]),
    .Y(\i57/n22 ));
 INVx1_ASAP7_75t_SL \i57/i487  (.A(n7[6]),
    .Y(\i57/n21 ));
 INVx2_ASAP7_75t_SL \i57/i488  (.A(n7[4]),
    .Y(\i57/n20 ));
 INVx3_ASAP7_75t_SL \i57/i489  (.A(n7[0]),
    .Y(\i57/n19 ));
 NAND2xp67_ASAP7_75t_SL \i57/i49  (.A(\i57/n555 ),
    .B(\i57/n425 ),
    .Y(\i57/n457 ));
 OR2x2_ASAP7_75t_SL \i57/i490  (.A(\i57/n128 ),
    .B(\i57/n232 ),
    .Y(\i57/n4 ));
 AND2x2_ASAP7_75t_SL \i57/i491  (.A(\i57/n22 ),
    .B(\i57/n23 ),
    .Y(\i57/n484 ));
 AOI222xp33_ASAP7_75t_R \i57/i492  (.A1(\i57/n63 ),
    .A2(\i57/n91 ),
    .B1(\i57/n85 ),
    .B2(\i57/n486 ),
    .C1(\i57/n74 ),
    .C2(\i57/n63 ),
    .Y(\i57/n487 ));
 AND2x4_ASAP7_75t_SL \i57/i493  (.A(\i57/n485 ),
    .B(\i57/n484 ),
    .Y(\i57/n486 ));
 AND2x2_ASAP7_75t_SL \i57/i494  (.A(n7[1]),
    .B(n7[0]),
    .Y(\i57/n485 ));
 INVx3_ASAP7_75t_SL \i57/i495  (.A(\i57/n486 ),
    .Y(\i57/n488 ));
 AOI211xp5_ASAP7_75t_SL \i57/i496  (.A1(\i57/n181 ),
    .A2(\i57/n486 ),
    .B(\i57/n279 ),
    .C(\i57/n326 ),
    .Y(\i57/n489 ));
 AOI222xp33_ASAP7_75t_SL \i57/i497  (.A1(\i57/n91 ),
    .A2(\i57/n526 ),
    .B1(\i57/n45 ),
    .B2(\i57/n53 ),
    .C1(\i57/n62 ),
    .C2(\i57/n486 ),
    .Y(\i57/n490 ));
 AOI22xp5_ASAP7_75t_SL \i57/i498  (.A1(\i57/n486 ),
    .A2(\i57/n124 ),
    .B1(\i57/n47 ),
    .B2(\i57/n88 ),
    .Y(\i57/n491 ));
 AOI221x1_ASAP7_75t_SL \i57/i499  (.A1(\i57/n7 ),
    .A2(\i57/n486 ),
    .B1(\i57/n6 ),
    .B2(\i57/n10 ),
    .C(\i57/n162 ),
    .Y(\i57/n492 ));
 AND2x4_ASAP7_75t_SL \i57/i5  (.A(\i57/n481 ),
    .B(\i57/n473 ),
    .Y(n6[3]));
 NAND2xp5_ASAP7_75t_SL \i57/i50  (.A(\i57/n368 ),
    .B(\i57/n398 ),
    .Y(\i57/n456 ));
 AOI22xp5_ASAP7_75t_SL \i57/i500  (.A1(\i57/n486 ),
    .A2(\i57/n65 ),
    .B1(\i57/n54 ),
    .B2(\i57/n62 ),
    .Y(\i57/n493 ));
 NAND2xp5_ASAP7_75t_SL \i57/i501  (.A(\i57/n486 ),
    .B(\i57/n74 ),
    .Y(\i57/n494 ));
 NAND2xp5_ASAP7_75t_SL \i57/i502  (.A(\i57/n486 ),
    .B(\i57/n91 ),
    .Y(\i57/n495 ));
 NAND2xp5_ASAP7_75t_SL \i57/i503  (.A(\i57/n486 ),
    .B(\i57/n83 ),
    .Y(\i57/n496 ));
 NAND2xp5_ASAP7_75t_SL \i57/i504  (.A(\i57/n486 ),
    .B(\i57/n43 ),
    .Y(\i57/n497 ));
 NOR2xp33_ASAP7_75t_SL \i57/i505  (.A(\i57/n486 ),
    .B(\i57/n49 ),
    .Y(\i57/n498 ));
 NAND2xp5_ASAP7_75t_SL \i57/i506  (.A(\i57/n76 ),
    .B(\i57/n486 ),
    .Y(\i57/n499 ));
 NOR2xp33_ASAP7_75t_L \i57/i507  (.A(\i57/n486 ),
    .B(\i57/n69 ),
    .Y(\i57/n500 ));
 NAND2xp5_ASAP7_75t_SL \i57/i508  (.A(\i57/n486 ),
    .B(\i57/n53 ),
    .Y(\i57/n501 ));
 NAND2xp5_ASAP7_75t_SL \i57/i509  (.A(\i57/n486 ),
    .B(\i57/n81 ),
    .Y(\i57/n502 ));
 INVx1_ASAP7_75t_SL \i57/i51  (.A(\i57/n540 ),
    .Y(\i57/n444 ));
 NAND2xp5_ASAP7_75t_SL \i57/i510  (.A(\i57/n486 ),
    .B(\i57/n62 ),
    .Y(\i57/n503 ));
 AND2x2_ASAP7_75t_SL \i57/i511  (.A(n7[3]),
    .B(\i57/n1 ),
    .Y(\i57/n504 ));
 AOI22xp5_ASAP7_75t_SL \i57/i512  (.A1(\i57/n486 ),
    .A2(\i57/n43 ),
    .B1(\i57/n56 ),
    .B2(\i57/n506 ),
    .Y(\i57/n507 ));
 AND2x4_ASAP7_75t_SL \i57/i513  (.A(\i57/n505 ),
    .B(\i57/n504 ),
    .Y(\i57/n506 ));
 NOR2xp33_ASAP7_75t_SL \i57/i514  (.A(\i57/n22 ),
    .B(n7[0]),
    .Y(\i57/n505 ));
 INVx3_ASAP7_75t_SL \i57/i515  (.A(\i57/n506 ),
    .Y(\i57/n508 ));
 AOI222xp33_ASAP7_75t_SL \i57/i516  (.A1(\i57/n526 ),
    .A2(\i57/n76 ),
    .B1(\i57/n6 ),
    .B2(\i57/n83 ),
    .C1(\i57/n506 ),
    .C2(\i57/n81 ),
    .Y(\i57/n509 ));
 OAI21xp33_ASAP7_75t_SL \i57/i517  (.A1(\i57/n506 ),
    .A2(\i57/n47 ),
    .B(\i57/n85 ),
    .Y(\i57/n510 ));
 AOI22xp33_ASAP7_75t_SL \i57/i518  (.A1(\i57/n65 ),
    .A2(\i57/n6 ),
    .B1(\i57/n506 ),
    .B2(\i57/n53 ),
    .Y(\i57/n511 ));
 AO22x1_ASAP7_75t_SL \i57/i519  (.A1(\i57/n62 ),
    .A2(\i57/n69 ),
    .B1(\i57/n83 ),
    .B2(\i57/n506 ),
    .Y(\i57/n512 ));
 INVxp67_ASAP7_75t_SL \i57/i52  (.A(\i57/n442 ),
    .Y(\i57/n443 ));
 AOI22xp5_ASAP7_75t_SL \i57/i520  (.A1(\i57/n88 ),
    .A2(\i57/n526 ),
    .B1(\i57/n43 ),
    .B2(\i57/n506 ),
    .Y(\i57/n513 ));
 AOI22xp5_ASAP7_75t_SL \i57/i521  (.A1(\i57/n51 ),
    .A2(\i57/n67 ),
    .B1(\i57/n506 ),
    .B2(\i57/n7 ),
    .Y(\i57/n514 ));
 NOR2xp33_ASAP7_75t_L \i57/i522  (.A(\i57/n506 ),
    .B(\i57/n63 ),
    .Y(\i57/n515 ));
 NOR2xp33_ASAP7_75t_SL \i57/i523  (.A(\i57/n67 ),
    .B(\i57/n506 ),
    .Y(\i57/n516 ));
 NAND2xp5_ASAP7_75t_SL \i57/i524  (.A(\i57/n74 ),
    .B(\i57/n506 ),
    .Y(\i57/n517 ));
 NAND2xp5_ASAP7_75t_SL \i57/i525  (.A(\i57/n56 ),
    .B(\i57/n506 ),
    .Y(\i57/n518 ));
 NAND2xp5_ASAP7_75t_SL \i57/i526  (.A(\i57/n51 ),
    .B(\i57/n506 ),
    .Y(\i57/n519 ));
 NAND2xp5_ASAP7_75t_SL \i57/i527  (.A(\i57/n62 ),
    .B(\i57/n506 ),
    .Y(\i57/n520 ));
 OAI22x1_ASAP7_75t_SL \i57/i528  (.A1(\i57/n3 ),
    .A2(\i57/n2 ),
    .B1(\i57/n84 ),
    .B2(\i57/n508 ),
    .Y(\i57/n521 ));
 OAI21xp5_ASAP7_75t_SL \i57/i529  (.A1(\i57/n55 ),
    .A2(\i57/n82 ),
    .B(\i57/n523 ),
    .Y(\i57/n524 ));
 NAND3xp33_ASAP7_75t_L \i57/i53  (.A(\i57/n381 ),
    .B(\i57/n347 ),
    .C(\i57/n392 ),
    .Y(\i57/n441 ));
 NOR2x1_ASAP7_75t_SL \i57/i530  (.A(\i57/n522 ),
    .B(\i57/n521 ),
    .Y(\i57/n523 ));
 OAI22xp5_ASAP7_75t_SL \i57/i531  (.A1(\i57/n48 ),
    .A2(\i57/n89 ),
    .B1(\i57/n86 ),
    .B2(\i57/n488 ),
    .Y(\i57/n522 ));
 NAND5xp2_ASAP7_75t_SL \i57/i532  (.A(\i57/n363 ),
    .B(\i57/n335 ),
    .C(\i57/n311 ),
    .D(\i57/n309 ),
    .E(\i57/n523 ),
    .Y(\i57/n525 ));
 INVx5_ASAP7_75t_SL \i57/i533  (.A(\i57/n60 ),
    .Y(\i57/n7 ));
 AND2x4_ASAP7_75t_SL \i57/i534  (.A(\i57/n32 ),
    .B(\i57/n28 ),
    .Y(\i57/n526 ));
 OAI211xp5_ASAP7_75t_SL \i57/i535  (.A1(\i57/n89 ),
    .A2(\i57/n156 ),
    .B(\i57/n527 ),
    .C(\i57/n182 ),
    .Y(\i57/n528 ));
 NAND2xp5_ASAP7_75t_SL \i57/i536  (.A(\i57/n7 ),
    .B(\i57/n526 ),
    .Y(\i57/n527 ));
 NAND4xp25_ASAP7_75t_SL \i57/i537  (.A(\i57/n527 ),
    .B(\i57/n115 ),
    .C(\i57/n204 ),
    .D(\i57/n146 ),
    .Y(\i57/n529 ));
 INVx2_ASAP7_75t_SL \i57/i538  (.A(\i57/n63 ),
    .Y(\i57/n530 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i57/i539  (.A1(\i57/n77 ),
    .A2(\i57/n531 ),
    .B(\i57/n7 ),
    .C(\i57/n72 ),
    .Y(\i57/n532 ));
 NAND3xp33_ASAP7_75t_L \i57/i54  (.A(\i57/n389 ),
    .B(\i57/n185 ),
    .C(\i57/n18 ),
    .Y(\i57/n440 ));
 NAND2x1_ASAP7_75t_SL \i57/i540  (.A(\i57/n44 ),
    .B(\i57/n530 ),
    .Y(\i57/n531 ));
 OAI31xp33_ASAP7_75t_SL \i57/i541  (.A1(\i57/n531 ),
    .A2(\i57/n72 ),
    .A3(\i57/n6 ),
    .B(\i57/n83 ),
    .Y(\i57/n533 ));
 NAND2xp5_ASAP7_75t_SL \i57/i542  (.A(\i57/n87 ),
    .B(\i57/n531 ),
    .Y(\i57/n534 ));
 OAI22xp5_ASAP7_75t_SL \i57/i543  (.A1(\i57/n92 ),
    .A2(\i57/n90 ),
    .B1(\i57/n46 ),
    .B2(\i57/n61 ),
    .Y(\i57/n535 ));
 AND2x2_ASAP7_75t_SL \i57/i544  (.A(\i57/n47 ),
    .B(\i57/n91 ),
    .Y(\i57/n536 ));
 NAND3xp33_ASAP7_75t_SL \i57/i545  (.A(\i57/n538 ),
    .B(\i57/n353 ),
    .C(\i57/n331 ),
    .Y(\i57/n539 ));
 NOR3xp33_ASAP7_75t_SL \i57/i546  (.A(\i57/n535 ),
    .B(\i57/n537 ),
    .C(\i57/n536 ),
    .Y(\i57/n538 ));
 OAI22xp5_ASAP7_75t_SL \i57/i547  (.A1(\i57/n42 ),
    .A2(\i57/n66 ),
    .B1(\i57/n530 ),
    .B2(\i57/n61 ),
    .Y(\i57/n537 ));
 NAND4xp25_ASAP7_75t_SL \i57/i548  (.A(\i57/n392 ),
    .B(\i57/n538 ),
    .C(\i57/n395 ),
    .D(\i57/n321 ),
    .Y(\i57/n540 ));
 NAND2xp5_ASAP7_75t_SL \i57/i549  (.A(\i57/n538 ),
    .B(\i57/n395 ),
    .Y(\i57/n541 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i57/i55  (.A1(\i57/n60 ),
    .A2(\i57/n52 ),
    .B(\i57/n532 ),
    .C(\i57/n400 ),
    .Y(\i57/n439 ));
 AND2x2_ASAP7_75t_SL \i57/i550  (.A(\i57/n0 ),
    .B(\i57/n20 ),
    .Y(\i57/n542 ));
 INVx3_ASAP7_75t_SL \i57/i551  (.A(\i57/n26 ),
    .Y(\i57/n543 ));
 AOI22xp5_ASAP7_75t_SL \i57/i552  (.A1(\i57/n544 ),
    .A2(\i57/n69 ),
    .B1(\i57/n83 ),
    .B2(\i57/n506 ),
    .Y(\i57/n545 ));
 AND2x4_ASAP7_75t_SL \i57/i553  (.A(\i57/n542 ),
    .B(\i57/n543 ),
    .Y(\i57/n544 ));
 O2A1O1Ixp33_ASAP7_75t_R \i57/i554  (.A1(\i57/n506 ),
    .A2(\i57/n45 ),
    .B(\i57/n544 ),
    .C(\i57/n229 ),
    .Y(\i57/n546 ));
 AOI22x1_ASAP7_75t_L \i57/i555  (.A1(\i57/n54 ),
    .A2(\i57/n544 ),
    .B1(\i57/n56 ),
    .B2(\i57/n526 ),
    .Y(\i57/n547 ));
 AOI22xp5_ASAP7_75t_SL \i57/i556  (.A1(\i57/n93 ),
    .A2(\i57/n544 ),
    .B1(\i57/n51 ),
    .B2(\i57/n72 ),
    .Y(\i57/n548 ));
 NAND2xp5_ASAP7_75t_SL \i57/i557  (.A(\i57/n63 ),
    .B(\i57/n544 ),
    .Y(\i57/n549 ));
 NAND2xp5_ASAP7_75t_SL \i57/i558  (.A(\i57/n79 ),
    .B(\i57/n544 ),
    .Y(\i57/n550 ));
 NAND2xp5_ASAP7_75t_SL \i57/i559  (.A(\i57/n544 ),
    .B(\i57/n45 ),
    .Y(\i57/n551 ));
 NAND2xp33_ASAP7_75t_SL \i57/i56  (.A(\i57/n406 ),
    .B(\i57/n399 ),
    .Y(\i57/n438 ));
 AOI221xp5_ASAP7_75t_SL \i57/i560  (.A1(\i57/n49 ),
    .A2(\i57/n544 ),
    .B1(\i57/n45 ),
    .B2(\i57/n43 ),
    .C(\i57/n244 ),
    .Y(\i57/n552 ));
 OAI31xp33_ASAP7_75t_SL \i57/i561  (.A1(\i57/n43 ),
    .A2(\i57/n51 ),
    .A3(\i57/n544 ),
    .B(\i57/n72 ),
    .Y(\i57/n553 ));
 NAND2xp5_ASAP7_75t_SL \i57/i562  (.A(\i57/n72 ),
    .B(\i57/n544 ),
    .Y(\i57/n554 ));
 AOI211xp5_ASAP7_75t_SL \i57/i563  (.A1(\i57/n544 ),
    .A2(\i57/n47 ),
    .B(\i57/n257 ),
    .C(\i57/n264 ),
    .Y(\i57/n555 ));
 AND4x1_ASAP7_75t_SL \i57/i564  (.A(\i57/n422 ),
    .B(\i57/n185 ),
    .C(\i57/n18 ),
    .D(\i57/n415 ),
    .Y(\i57/n556 ));
 AND3x1_ASAP7_75t_SL \i57/i565  (.A(\i57/n527 ),
    .B(\i57/n146 ),
    .C(\i57/n204 ),
    .Y(\i57/n557 ));
 AND4x1_ASAP7_75t_SL \i57/i566  (.A(\i57/n198 ),
    .B(\i57/n196 ),
    .C(\i57/n145 ),
    .D(\i57/n549 ),
    .Y(\i57/n558 ));
 NOR2xp33_ASAP7_75t_SL \i57/i57  (.A(\i57/n384 ),
    .B(\i57/n403 ),
    .Y(\i57/n437 ));
 NAND5xp2_ASAP7_75t_SL \i57/i58  (.A(\i57/n342 ),
    .B(\i57/n303 ),
    .C(\i57/n293 ),
    .D(\i57/n553 ),
    .E(\i57/n322 ),
    .Y(\i57/n436 ));
 NOR3xp33_ASAP7_75t_SL \i57/i59  (.A(\i57/n355 ),
    .B(\i57/n268 ),
    .C(\i57/n328 ),
    .Y(\i57/n435 ));
 AND3x4_ASAP7_75t_SL \i57/i6  (.A(\i57/n556 ),
    .B(\i57/n475 ),
    .C(\i57/n472 ),
    .Y(n6[4]));
 NAND2xp33_ASAP7_75t_SL \i57/i60  (.A(\i57/n383 ),
    .B(\i57/n406 ),
    .Y(\i57/n434 ));
 NAND4xp25_ASAP7_75t_SL \i57/i61  (.A(\i57/n393 ),
    .B(\i57/n369 ),
    .C(\i57/n299 ),
    .D(\i57/n317 ),
    .Y(\i57/n433 ));
 NOR3xp33_ASAP7_75t_SL \i57/i62  (.A(\i57/n405 ),
    .B(\i57/n366 ),
    .C(\i57/n388 ),
    .Y(\i57/n432 ));
 NAND5xp2_ASAP7_75t_SL \i57/i63  (.A(\i57/n373 ),
    .B(\i57/n343 ),
    .C(\i57/n338 ),
    .D(\i57/n218 ),
    .E(\i57/n306 ),
    .Y(\i57/n431 ));
 NOR4xp25_ASAP7_75t_SL \i57/i64  (.A(\i57/n360 ),
    .B(\i57/n361 ),
    .C(\i57/n220 ),
    .D(\i57/n188 ),
    .Y(\i57/n430 ));
 NAND2xp33_ASAP7_75t_SL \i57/i65  (.A(\i57/n410 ),
    .B(\i57/n387 ),
    .Y(\i57/n429 ));
 NOR3x1_ASAP7_75t_SL \i57/i66  (.A(\i57/n524 ),
    .B(\i57/n341 ),
    .C(\i57/n378 ),
    .Y(\i57/n442 ));
 INVxp67_ASAP7_75t_SL \i57/i67  (.A(\i57/n427 ),
    .Y(\i57/n428 ));
 INVx1_ASAP7_75t_SL \i57/i68  (.A(\i57/n423 ),
    .Y(\i57/n424 ));
 INVxp67_ASAP7_75t_SL \i57/i69  (.A(\i57/n421 ),
    .Y(\i57/n422 ));
 AND5x2_ASAP7_75t_SL \i57/i7  (.A(\i57/n442 ),
    .B(\i57/n463 ),
    .C(\i57/n432 ),
    .D(\i57/n464 ),
    .E(\i57/n462 ),
    .Y(n6[1]));
 INVx1_ASAP7_75t_SL \i57/i70  (.A(\i57/n419 ),
    .Y(\i57/n420 ));
 NOR3xp33_ASAP7_75t_SL \i57/i71  (.A(\i57/n382 ),
    .B(\i57/n17 ),
    .C(\i57/n234 ),
    .Y(\i57/n418 ));
 NAND3xp33_ASAP7_75t_SL \i57/i72  (.A(\i57/n266 ),
    .B(\i57/n533 ),
    .C(\i57/n552 ),
    .Y(\i57/n417 ));
 NAND2xp5_ASAP7_75t_SL \i57/i73  (.A(\i57/n370 ),
    .B(\i57/n385 ),
    .Y(\i57/n416 ));
 NOR2xp33_ASAP7_75t_SL \i57/i74  (.A(\i57/n394 ),
    .B(\i57/n362 ),
    .Y(\i57/n415 ));
 NOR2xp33_ASAP7_75t_SL \i57/i75  (.A(\i57/n354 ),
    .B(\i57/n298 ),
    .Y(\i57/n414 ));
 NOR5xp2_ASAP7_75t_SL \i57/i76  (.A(\i57/n288 ),
    .B(\i57/n512 ),
    .C(\i57/n220 ),
    .D(\i57/n261 ),
    .E(\i57/n259 ),
    .Y(\i57/n413 ));
 NOR2xp33_ASAP7_75t_SL \i57/i77  (.A(\i57/n340 ),
    .B(\i57/n364 ),
    .Y(\i57/n412 ));
 AOI211xp5_ASAP7_75t_SL \i57/i78  (.A1(\i57/n327 ),
    .A2(\i57/n112 ),
    .B(\i57/n281 ),
    .C(\i57/n235 ),
    .Y(\i57/n411 ));
 NAND2xp5_ASAP7_75t_SL \i57/i79  (.A(\i57/n292 ),
    .B(\i57/n386 ),
    .Y(\i57/n427 ));
 NOR2xp33_ASAP7_75t_SL \i57/i8  (.A(\i57/n454 ),
    .B(\i57/n482 ),
    .Y(\i57/n483 ));
 NAND3xp33_ASAP7_75t_SL \i57/i80  (.A(\i57/n367 ),
    .B(\i57/n348 ),
    .C(\i57/n320 ),
    .Y(\i57/n426 ));
 NOR2x1_ASAP7_75t_SL \i57/i81  (.A(\i57/n375 ),
    .B(\i57/n302 ),
    .Y(\i57/n425 ));
 AND3x1_ASAP7_75t_SL \i57/i82  (.A(\i57/n534 ),
    .B(\i57/n492 ),
    .C(\i57/n491 ),
    .Y(\i57/n423 ));
 NAND3xp33_ASAP7_75t_SL \i57/i83  (.A(\i57/n299 ),
    .B(\i57/n297 ),
    .C(\i57/n558 ),
    .Y(\i57/n421 ));
 NOR3x1_ASAP7_75t_SL \i57/i84  (.A(\i57/n301 ),
    .B(\i57/n324 ),
    .C(\i57/n231 ),
    .Y(\i57/n419 ));
 INVxp33_ASAP7_75t_SL \i57/i85  (.A(\i57/n407 ),
    .Y(\i57/n408 ));
 OAI211xp5_ASAP7_75t_SL \i57/i86  (.A1(\i57/n508 ),
    .A2(\i57/n180 ),
    .B(\i57/n316 ),
    .C(\i57/n251 ),
    .Y(\i57/n404 ));
 NAND4xp25_ASAP7_75t_SL \i57/i87  (.A(\i57/n289 ),
    .B(\i57/n325 ),
    .C(\i57/n291 ),
    .D(\i57/n249 ),
    .Y(\i57/n403 ));
 NOR3xp33_ASAP7_75t_SL \i57/i88  (.A(\i57/n380 ),
    .B(\i57/n307 ),
    .C(\i57/n4 ),
    .Y(\i57/n402 ));
 NAND4xp25_ASAP7_75t_SL \i57/i89  (.A(\i57/n348 ),
    .B(\i57/n547 ),
    .C(\i57/n313 ),
    .D(\i57/n507 ),
    .Y(\i57/n401 ));
 AND4x2_ASAP7_75t_SL \i57/i9  (.A(\i57/n472 ),
    .B(\i57/n480 ),
    .C(\i57/n479 ),
    .D(\i57/n430 ),
    .Y(n6[5]));
 NOR3xp33_ASAP7_75t_SL \i57/i90  (.A(\i57/n315 ),
    .B(\i57/n269 ),
    .C(\i57/n273 ),
    .Y(\i57/n400 ));
 NOR4xp25_ASAP7_75t_SL \i57/i91  (.A(\i57/n377 ),
    .B(\i57/n339 ),
    .C(\i57/n226 ),
    .D(\i57/n521 ),
    .Y(\i57/n399 ));
 NOR3xp33_ASAP7_75t_SL \i57/i92  (.A(\i57/n308 ),
    .B(\i57/n253 ),
    .C(\i57/n280 ),
    .Y(\i57/n410 ));
 NOR2xp33_ASAP7_75t_SL \i57/i93  (.A(\i57/n388 ),
    .B(\i57/n529 ),
    .Y(\i57/n398 ));
 NOR2xp33_ASAP7_75t_SL \i57/i94  (.A(\i57/n376 ),
    .B(\i57/n358 ),
    .Y(\i57/n397 ));
 NAND5xp2_ASAP7_75t_SL \i57/i95  (.A(\i57/n295 ),
    .B(\i57/n490 ),
    .C(\i57/n217 ),
    .D(\i57/n225 ),
    .E(\i57/n218 ),
    .Y(\i57/n409 ));
 NOR3xp33_ASAP7_75t_SL \i57/i96  (.A(\i57/n349 ),
    .B(\i57/n224 ),
    .C(\i57/n107 ),
    .Y(\i57/n407 ));
 NOR2xp33_ASAP7_75t_L \i57/i97  (.A(\i57/n351 ),
    .B(\i57/n334 ),
    .Y(\i57/n406 ));
 NOR2xp33_ASAP7_75t_R \i57/i98  (.A(\i57/n341 ),
    .B(\i57/n524 ),
    .Y(\i57/n396 ));
 NAND2xp5_ASAP7_75t_SL \i57/i99  (.A(\i57/n357 ),
    .B(\i57/n391 ),
    .Y(\i57/n405 ));
 OAI22xp5_ASAP7_75t_SL i570 (.A1(n761),
    .A2(n779),
    .B1(n780),
    .B2(n760),
    .Y(n902));
 XOR2xp5_ASAP7_75t_SL i571 (.A(n334),
    .B(n589),
    .Y(n901));
 AOI22xp5_ASAP7_75t_SL i572 (.A1(n760),
    .A2(n1176),
    .B1(n789),
    .B2(n761),
    .Y(n900));
 AOI22xp5_ASAP7_75t_SL i573 (.A1(n869),
    .A2(n800),
    .B1(n868),
    .B2(n801),
    .Y(n899));
 XOR2xp5_ASAP7_75t_SL i574 (.A(n314),
    .B(n328),
    .Y(n898));
 AOI22xp5_ASAP7_75t_SL i575 (.A1(n1153),
    .A2(n522),
    .B1(n521),
    .B2(n227),
    .Y(n897));
 AOI22xp5_ASAP7_75t_SL i576 (.A1(n526),
    .A2(n493),
    .B1(n525),
    .B2(n492),
    .Y(n896));
 XOR2xp5_ASAP7_75t_SL i577 (.A(n304),
    .B(n295),
    .Y(n895));
 AOI22xp5_ASAP7_75t_SL i578 (.A1(n1155),
    .A2(n536),
    .B1(n535),
    .B2(n226),
    .Y(n894));
 OAI22xp5_ASAP7_75t_SL i579 (.A1(n1211),
    .A2(n504),
    .B1(n505),
    .B2(n479),
    .Y(n893));
 INVx1_ASAP7_75t_SL \i58/i0  (.A(n5[5]),
    .Y(\i58/n0 ));
 INVx2_ASAP7_75t_SL \i58/i1  (.A(\i58/n57 ),
    .Y(\i58/n1 ));
 AND4x2_ASAP7_75t_SL \i58/i10  (.A(\i58/n459 ),
    .B(\i58/n460 ),
    .C(\i58/n456 ),
    .D(\i58/n457 ),
    .Y(n4[7]));
 NOR2xp33_ASAP7_75t_SL \i58/i100  (.A(\i58/n536 ),
    .B(\i58/n358 ),
    .Y(\i58/n385 ));
 NAND2xp5_ASAP7_75t_SL \i58/i101  (.A(\i58/n344 ),
    .B(\i58/n380 ),
    .Y(\i58/n393 ));
 INVxp33_ASAP7_75t_SL \i58/i102  (.A(\i58/n382 ),
    .Y(\i58/n383 ));
 INVxp67_ASAP7_75t_SL \i58/i103  (.A(\i58/n378 ),
    .Y(\i58/n379 ));
 NOR3xp33_ASAP7_75t_SL \i58/i104  (.A(\i58/n513 ),
    .B(\i58/n205 ),
    .C(\i58/n86 ),
    .Y(\i58/n374 ));
 OAI211xp5_ASAP7_75t_SL \i58/i105  (.A1(\i58/n62 ),
    .A2(\i58/n165 ),
    .B(\i58/n501 ),
    .C(\i58/n285 ),
    .Y(\i58/n373 ));
 NOR2xp33_ASAP7_75t_SL \i58/i106  (.A(\i58/n324 ),
    .B(\i58/n18 ),
    .Y(\i58/n372 ));
 OAI21xp5_ASAP7_75t_SL \i58/i107  (.A1(\i58/n54 ),
    .A2(\i58/n72 ),
    .B(\i58/n326 ),
    .Y(\i58/n371 ));
 NOR4xp25_ASAP7_75t_SL \i58/i108  (.A(\i58/n230 ),
    .B(\i58/n231 ),
    .C(\i58/n196 ),
    .D(\i58/n221 ),
    .Y(\i58/n370 ));
 NAND2xp33_ASAP7_75t_SL \i58/i109  (.A(\i58/n556 ),
    .B(\i58/n328 ),
    .Y(\i58/n369 ));
 NAND4xp25_ASAP7_75t_SL \i58/i11  (.A(\i58/n450 ),
    .B(\i58/n387 ),
    .C(\i58/n376 ),
    .D(\i58/n481 ),
    .Y(\i58/n474 ));
 NOR3xp33_ASAP7_75t_SL \i58/i110  (.A(\i58/n524 ),
    .B(\i58/n120 ),
    .C(\i58/n175 ),
    .Y(\i58/n368 ));
 NAND2xp5_ASAP7_75t_SL \i58/i111  (.A(\i58/n216 ),
    .B(\i58/n260 ),
    .Y(\i58/n367 ));
 NOR2xp33_ASAP7_75t_L \i58/i112  (.A(\i58/n270 ),
    .B(\i58/n292 ),
    .Y(\i58/n384 ));
 OAI211xp5_ASAP7_75t_SL \i58/i113  (.A1(\i58/n45 ),
    .A2(\i58/n54 ),
    .B(\i58/n219 ),
    .C(\i58/n208 ),
    .Y(\i58/n366 ));
 NAND3xp33_ASAP7_75t_L \i58/i114  (.A(\i58/n247 ),
    .B(\i58/n545 ),
    .C(\i58/n294 ),
    .Y(\i58/n365 ));
 NAND2xp5_ASAP7_75t_SL \i58/i115  (.A(\i58/n515 ),
    .B(\i58/n219 ),
    .Y(\i58/n364 ));
 NAND2xp5_ASAP7_75t_L \i58/i116  (.A(\i58/n502 ),
    .B(\i58/n512 ),
    .Y(\i58/n363 ));
 NOR3xp33_ASAP7_75t_SL \i58/i117  (.A(\i58/n289 ),
    .B(\i58/n197 ),
    .C(\i58/n213 ),
    .Y(\i58/n362 ));
 NOR3xp33_ASAP7_75t_SL \i58/i118  (.A(\i58/n17 ),
    .B(\i58/n184 ),
    .C(\i58/n170 ),
    .Y(\i58/n361 ));
 NOR4xp25_ASAP7_75t_SL \i58/i119  (.A(\i58/n17 ),
    .B(\i58/n198 ),
    .C(\i58/n188 ),
    .D(\i58/n89 ),
    .Y(\i58/n360 ));
 NOR3xp33_ASAP7_75t_SL \i58/i12  (.A(\i58/n433 ),
    .B(\i58/n463 ),
    .C(\i58/n446 ),
    .Y(\i58/n473 ));
 AOI211xp5_ASAP7_75t_SL \i58/i120  (.A1(\i58/n105 ),
    .A2(\i58/n68 ),
    .B(\i58/n226 ),
    .C(\i58/n217 ),
    .Y(\i58/n382 ));
 NOR3xp33_ASAP7_75t_SL \i58/i121  (.A(\i58/n252 ),
    .B(\i58/n120 ),
    .C(\i58/n234 ),
    .Y(\i58/n381 ));
 NOR2xp33_ASAP7_75t_L \i58/i122  (.A(\i58/n213 ),
    .B(\i58/n333 ),
    .Y(\i58/n359 ));
 NOR2xp33_ASAP7_75t_SL \i58/i123  (.A(\i58/n258 ),
    .B(\i58/n321 ),
    .Y(\i58/n380 ));
 NOR2xp33_ASAP7_75t_SL \i58/i124  (.A(\i58/n264 ),
    .B(\i58/n327 ),
    .Y(\i58/n378 ));
 NAND2xp5_ASAP7_75t_SL \i58/i125  (.A(\i58/n208 ),
    .B(\i58/n500 ),
    .Y(\i58/n377 ));
 NOR2xp67_ASAP7_75t_SL \i58/i126  (.A(\i58/n307 ),
    .B(\i58/n329 ),
    .Y(\i58/n376 ));
 NOR3x1_ASAP7_75t_SL \i58/i127  (.A(\i58/n523 ),
    .B(\i58/n513 ),
    .C(\i58/n527 ),
    .Y(\i58/n375 ));
 INVx1_ASAP7_75t_SL \i58/i128  (.A(\i58/n354 ),
    .Y(\i58/n355 ));
 NOR2xp33_ASAP7_75t_SL \i58/i129  (.A(\i58/n521 ),
    .B(\i58/n302 ),
    .Y(\i58/n352 ));
 AND2x2_ASAP7_75t_SL \i58/i13  (.A(\i58/n468 ),
    .B(\i58/n469 ),
    .Y(n4[2]));
 NAND5xp2_ASAP7_75t_SL \i58/i130  (.A(\i58/n87 ),
    .B(\i58/n189 ),
    .C(\i58/n154 ),
    .D(\i58/n156 ),
    .E(\i58/n182 ),
    .Y(\i58/n351 ));
 NOR2xp33_ASAP7_75t_SL \i58/i131  (.A(\i58/n303 ),
    .B(\i58/n537 ),
    .Y(\i58/n350 ));
 OAI211xp5_ASAP7_75t_SL \i58/i132  (.A1(\i58/n45 ),
    .A2(\i58/n168 ),
    .B(\i58/n480 ),
    .C(\i58/n251 ),
    .Y(\i58/n349 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i58/i133  (.A1(\i58/n69 ),
    .A2(\i58/n183 ),
    .B(\i58/n6 ),
    .C(\i58/n244 ),
    .Y(\i58/n348 ));
 NAND3xp33_ASAP7_75t_SL \i58/i134  (.A(\i58/n547 ),
    .B(\i58/n236 ),
    .C(\i58/n227 ),
    .Y(\i58/n347 ));
 OAI21xp5_ASAP7_75t_SL \i58/i135  (.A1(\i58/n53 ),
    .A2(\i58/n76 ),
    .B(\i58/n331 ),
    .Y(\i58/n358 ));
 NOR3xp33_ASAP7_75t_SL \i58/i136  (.A(\i58/n261 ),
    .B(\i58/n212 ),
    .C(\i58/n218 ),
    .Y(\i58/n346 ));
 NAND3xp33_ASAP7_75t_L \i58/i137  (.A(\i58/n504 ),
    .B(\i58/n208 ),
    .C(\i58/n296 ),
    .Y(\i58/n345 ));
 NOR3xp33_ASAP7_75t_SL \i58/i138  (.A(\i58/n273 ),
    .B(\i58/n249 ),
    .C(\i58/n212 ),
    .Y(\i58/n344 ));
 AOI211xp5_ASAP7_75t_SL \i58/i139  (.A1(\i58/n534 ),
    .A2(\i58/n75 ),
    .B(\i58/n315 ),
    .C(\i58/n121 ),
    .Y(\i58/n343 ));
 NOR3xp33_ASAP7_75t_SL \i58/i14  (.A(\i58/n447 ),
    .B(\i58/n393 ),
    .C(\i58/n451 ),
    .Y(\i58/n472 ));
 OAI221xp5_ASAP7_75t_SL \i58/i140  (.A1(\i58/n165 ),
    .A2(\i58/n45 ),
    .B1(\i58/n108 ),
    .B2(\i58/n514 ),
    .C(\i58/n174 ),
    .Y(\i58/n342 ));
 AOI211xp5_ASAP7_75t_SL \i58/i141  (.A1(\i58/n532 ),
    .A2(\i58/n44 ),
    .B(\i58/n246 ),
    .C(\i58/n253 ),
    .Y(\i58/n341 ));
 NAND2xp33_ASAP7_75t_SL \i58/i142  (.A(\i58/n271 ),
    .B(\i58/n268 ),
    .Y(\i58/n340 ));
 NOR2xp33_ASAP7_75t_SL \i58/i143  (.A(\i58/n314 ),
    .B(\i58/n279 ),
    .Y(\i58/n339 ));
 NAND4xp25_ASAP7_75t_SL \i58/i144  (.A(\i58/n15 ),
    .B(\i58/n107 ),
    .C(\i58/n553 ),
    .D(\i58/n139 ),
    .Y(\i58/n338 ));
 O2A1O1Ixp33_ASAP7_75t_R \i58/i145  (.A1(\i58/n71 ),
    .A2(\i58/n11 ),
    .B(\i58/n1 ),
    .C(\i58/n66 ),
    .Y(\i58/n337 ));
 OAI221xp5_ASAP7_75t_SL \i58/i146  (.A1(\i58/n237 ),
    .A2(\i58/n84 ),
    .B1(\i58/n10 ),
    .B2(\i58/n78 ),
    .C(\i58/n548 ),
    .Y(\i58/n336 ));
 NAND4xp25_ASAP7_75t_SL \i58/i147  (.A(\i58/n543 ),
    .B(\i58/n204 ),
    .C(\i58/n176 ),
    .D(\i58/n190 ),
    .Y(\i58/n335 ));
 NOR2xp67_ASAP7_75t_SL \i58/i148  (.A(\i58/n281 ),
    .B(\i58/n290 ),
    .Y(\i58/n357 ));
 NAND2xp33_ASAP7_75t_L \i58/i149  (.A(\i58/n320 ),
    .B(\i58/n222 ),
    .Y(\i58/n334 ));
 NOR3xp33_ASAP7_75t_SL \i58/i15  (.A(\i58/n425 ),
    .B(\i58/n430 ),
    .C(\i58/n408 ),
    .Y(\i58/n471 ));
 NOR2x1_ASAP7_75t_SL \i58/i150  (.A(\i58/n299 ),
    .B(\i58/n317 ),
    .Y(\i58/n356 ));
 NAND2xp5_ASAP7_75t_SL \i58/i151  (.A(\i58/n263 ),
    .B(\i58/n210 ),
    .Y(\i58/n354 ));
 NOR3xp33_ASAP7_75t_SL \i58/i152  (.A(\i58/n221 ),
    .B(\i58/n202 ),
    .C(\i58/n195 ),
    .Y(\i58/n353 ));
 NOR2xp67_ASAP7_75t_SL \i58/i153  (.A(\i58/n262 ),
    .B(\i58/n269 ),
    .Y(\i58/n19 ));
 INVxp67_ASAP7_75t_SL \i58/i154  (.A(\i58/n329 ),
    .Y(\i58/n330 ));
 INVxp33_ASAP7_75t_SL \i58/i155  (.A(\i58/n327 ),
    .Y(\i58/n328 ));
 INVx1_ASAP7_75t_SL \i58/i156  (.A(\i58/n536 ),
    .Y(\i58/n325 ));
 INVxp67_ASAP7_75t_SL \i58/i157  (.A(\i58/n321 ),
    .Y(\i58/n322 ));
 INVxp67_ASAP7_75t_SL \i58/i158  (.A(\i58/n18 ),
    .Y(\i58/n320 ));
 INVxp67_ASAP7_75t_SL \i58/i159  (.A(\i58/n318 ),
    .Y(\i58/n319 ));
 NOR3xp33_ASAP7_75t_SL \i58/i16  (.A(\i58/n436 ),
    .B(\i58/n438 ),
    .C(\i58/n420 ),
    .Y(\i58/n470 ));
 NAND2xp5_ASAP7_75t_SL \i58/i160  (.A(\i58/n545 ),
    .B(\i58/n542 ),
    .Y(\i58/n317 ));
 AOI21xp5_ASAP7_75t_SL \i58/i161  (.A1(\i58/n172 ),
    .A2(\i58/n85 ),
    .B(\i58/n249 ),
    .Y(\i58/n316 ));
 OAI22xp5_ASAP7_75t_SL \i58/i162  (.A1(\i58/n103 ),
    .A2(\i58/n134 ),
    .B1(\i58/n80 ),
    .B2(\i58/n118 ),
    .Y(\i58/n315 ));
 NAND4xp25_ASAP7_75t_SL \i58/i163  (.A(\i58/n178 ),
    .B(\i58/n507 ),
    .C(\i58/n129 ),
    .D(\i58/n491 ),
    .Y(\i58/n314 ));
 NAND3xp33_ASAP7_75t_SL \i58/i164  (.A(\i58/n126 ),
    .B(\i58/n138 ),
    .C(\i58/n7 ),
    .Y(\i58/n313 ));
 NAND3xp33_ASAP7_75t_SL \i58/i165  (.A(\i58/n164 ),
    .B(\i58/n177 ),
    .C(\i58/n47 ),
    .Y(\i58/n312 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i58/i166  (.A1(\i58/n48 ),
    .A2(\i58/n42 ),
    .B(\i58/n532 ),
    .C(\i58/n217 ),
    .Y(\i58/n311 ));
 OAI31xp33_ASAP7_75t_SL \i58/i167  (.A1(\i58/n11 ),
    .A2(\i58/n66 ),
    .A3(\i58/n511 ),
    .B(\i58/n77 ),
    .Y(\i58/n310 ));
 NOR2xp33_ASAP7_75t_SL \i58/i168  (.A(\i58/n527 ),
    .B(\i58/n228 ),
    .Y(\i58/n309 ));
 OAI21xp5_ASAP7_75t_SL \i58/i169  (.A1(\i58/n80 ),
    .A2(\i58/n146 ),
    .B(\i58/n506 ),
    .Y(\i58/n308 ));
 NOR4xp25_ASAP7_75t_SL \i58/i17  (.A(\i58/n417 ),
    .B(\i58/n405 ),
    .C(\i58/n409 ),
    .D(\i58/n419 ),
    .Y(\i58/n469 ));
 NAND4xp25_ASAP7_75t_SL \i58/i170  (.A(\i58/n193 ),
    .B(\i58/n140 ),
    .C(\i58/n127 ),
    .D(\i58/n549 ),
    .Y(\i58/n307 ));
 AOI211xp5_ASAP7_75t_SL \i58/i171  (.A1(\i58/n42 ),
    .A2(\i58/n1 ),
    .B(\i58/n137 ),
    .C(\i58/n131 ),
    .Y(\i58/n306 ));
 NOR2xp33_ASAP7_75t_L \i58/i172  (.A(\i58/n201 ),
    .B(\i58/n242 ),
    .Y(\i58/n305 ));
 NOR2xp33_ASAP7_75t_L \i58/i173  (.A(\i58/n200 ),
    .B(\i58/n220 ),
    .Y(\i58/n304 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i58/i174  (.A1(\i58/n62 ),
    .A2(\i58/n5 ),
    .B(\i58/n49 ),
    .C(\i58/n245 ),
    .Y(\i58/n303 ));
 NAND3xp33_ASAP7_75t_SL \i58/i175  (.A(\i58/n502 ),
    .B(\i58/n176 ),
    .C(\i58/n493 ),
    .Y(\i58/n302 ));
 NOR3xp33_ASAP7_75t_SL \i58/i176  (.A(\i58/n225 ),
    .B(\i58/n143 ),
    .C(\i58/n191 ),
    .Y(\i58/n301 ));
 NAND4xp25_ASAP7_75t_SL \i58/i177  (.A(\i58/n486 ),
    .B(\i58/n113 ),
    .C(\i58/n14 ),
    .D(\i58/n16 ),
    .Y(\i58/n300 ));
 OAI211xp5_ASAP7_75t_SL \i58/i178  (.A1(\i58/n55 ),
    .A2(\i58/n546 ),
    .B(\i58/n96 ),
    .C(\i58/n488 ),
    .Y(\i58/n299 ));
 OAI31xp33_ASAP7_75t_SL \i58/i179  (.A1(\i58/n41 ),
    .A2(\i58/n50 ),
    .A3(\i58/n532 ),
    .B(\i58/n66 ),
    .Y(\i58/n298 ));
 NOR5xp2_ASAP7_75t_SL \i58/i18  (.A(\i58/n445 ),
    .B(\i58/n414 ),
    .C(\i58/n447 ),
    .D(\i58/n397 ),
    .E(\i58/n379 ),
    .Y(\i58/n468 ));
 AOI221xp5_ASAP7_75t_SL \i58/i180  (.A1(\i58/n157 ),
    .A2(\i58/n56 ),
    .B1(\i58/n52 ),
    .B2(\i58/n85 ),
    .C(\i58/n142 ),
    .Y(\i58/n297 ));
 NOR2xp33_ASAP7_75t_SL \i58/i181  (.A(\i58/n125 ),
    .B(\i58/n526 ),
    .Y(\i58/n296 ));
 OAI221xp5_ASAP7_75t_SL \i58/i182  (.A1(\i58/n5 ),
    .A2(\i58/n40 ),
    .B1(\i58/n51 ),
    .B2(\i58/n498 ),
    .C(\i58/n485 ),
    .Y(\i58/n333 ));
 AOI222xp33_ASAP7_75t_SL \i58/i183  (.A1(\i58/n511 ),
    .A2(\i58/n533 ),
    .B1(\i58/n71 ),
    .B2(\i58/n68 ),
    .C1(\i58/n61 ),
    .C2(\i58/n75 ),
    .Y(\i58/n332 ));
 NOR2x1_ASAP7_75t_SL \i58/i184  (.A(\i58/n525 ),
    .B(\i58/n211 ),
    .Y(\i58/n331 ));
 NAND2xp5_ASAP7_75t_SL \i58/i185  (.A(\i58/n239 ),
    .B(\i58/n199 ),
    .Y(\i58/n329 ));
 OAI221xp5_ASAP7_75t_SL \i58/i186  (.A1(\i58/n546 ),
    .A2(\i58/n53 ),
    .B1(\i58/n60 ),
    .B2(\i58/n54 ),
    .C(\i58/n7 ),
    .Y(\i58/n327 ));
 OAI21xp5_ASAP7_75t_SL \i58/i187  (.A1(\i58/n56 ),
    .A2(\i58/n117 ),
    .B(\i58/n166 ),
    .Y(\i58/n326 ));
 NOR2xp33_ASAP7_75t_SL \i58/i188  (.A(\i58/n120 ),
    .B(\i58/n252 ),
    .Y(\i58/n295 ));
 NOR2xp33_ASAP7_75t_SL \i58/i189  (.A(\i58/n195 ),
    .B(\i58/n221 ),
    .Y(\i58/n294 ));
 NOR3xp33_ASAP7_75t_SL \i58/i19  (.A(\i58/n386 ),
    .B(\i58/n448 ),
    .C(\i58/n461 ),
    .Y(\i58/n467 ));
 NAND2xp5_ASAP7_75t_SL \i58/i190  (.A(\i58/n206 ),
    .B(\i58/n207 ),
    .Y(\i58/n324 ));
 NAND2xp5_ASAP7_75t_SL \i58/i191  (.A(\i58/n229 ),
    .B(\i58/n245 ),
    .Y(\i58/n323 ));
 OAI221xp5_ASAP7_75t_SL \i58/i192  (.A1(\i58/n47 ),
    .A2(\i58/n82 ),
    .B1(\i58/n64 ),
    .B2(\i58/n80 ),
    .C(\i58/n133 ),
    .Y(\i58/n321 ));
 NAND2x1_ASAP7_75t_SL \i58/i193  (.A(\i58/n235 ),
    .B(\i58/n504 ),
    .Y(\i58/n18 ));
 NAND3xp33_ASAP7_75t_SL \i58/i194  (.A(\i58/n132 ),
    .B(\i58/n128 ),
    .C(\i58/n124 ),
    .Y(\i58/n17 ));
 NOR2xp33_ASAP7_75t_SL \i58/i195  (.A(\i58/n253 ),
    .B(\i58/n246 ),
    .Y(\i58/n293 ));
 OAI211xp5_ASAP7_75t_SL \i58/i196  (.A1(\i58/n74 ),
    .A2(\i58/n65 ),
    .B(\i58/n194 ),
    .C(\i58/n12 ),
    .Y(\i58/n318 ));
 INVxp67_ASAP7_75t_SL \i58/i197  (.A(\i58/n290 ),
    .Y(\i58/n291 ));
 INVxp67_ASAP7_75t_SL \i58/i198  (.A(\i58/n516 ),
    .Y(\i58/n289 ));
 INVxp67_ASAP7_75t_SL \i58/i199  (.A(\i58/n287 ),
    .Y(\i58/n288 ));
 INVx1_ASAP7_75t_SL \i58/i2  (.A(\i58/n532 ),
    .Y(\i58/n2 ));
 NOR3xp33_ASAP7_75t_SL \i58/i20  (.A(\i58/n427 ),
    .B(\i58/n414 ),
    .C(\i58/n452 ),
    .Y(\i58/n466 ));
 INVx2_ASAP7_75t_SL \i58/i200  (.A(\i58/n285 ),
    .Y(\i58/n286 ));
 INVx1_ASAP7_75t_SL \i58/i201  (.A(\i58/n283 ),
    .Y(\i58/n284 ));
 OAI22xp5_ASAP7_75t_SL \i58/i202  (.A1(\i58/n60 ),
    .A2(\i58/n115 ),
    .B1(\i58/n69 ),
    .B2(\i58/n65 ),
    .Y(\i58/n281 ));
 AOI21xp5_ASAP7_75t_SL \i58/i203  (.A1(\i58/n101 ),
    .A2(\i58/n70 ),
    .B(\i58/n121 ),
    .Y(\i58/n280 ));
 OAI22xp5_ASAP7_75t_SL \i58/i204  (.A1(\i58/n54 ),
    .A2(\i58/n98 ),
    .B1(\i58/n53 ),
    .B2(\i58/n180 ),
    .Y(\i58/n279 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i58/i205  (.A1(\i58/n534 ),
    .A2(\i58/n63 ),
    .B(\i58/n68 ),
    .C(\i58/n91 ),
    .Y(\i58/n278 ));
 AOI21xp5_ASAP7_75t_SL \i58/i206  (.A1(\i58/n167 ),
    .A2(\i58/n534 ),
    .B(\i58/n232 ),
    .Y(\i58/n277 ));
 AOI22xp5_ASAP7_75t_SL \i58/i207  (.A1(\i58/n50 ),
    .A2(\i58/n102 ),
    .B1(\i58/n73 ),
    .B2(\i58/n160 ),
    .Y(\i58/n276 ));
 AOI211xp5_ASAP7_75t_SL \i58/i208  (.A1(\i58/n50 ),
    .A2(\i58/n531 ),
    .B(\i58/n121 ),
    .C(\i58/n93 ),
    .Y(\i58/n275 ));
 OAI22xp5_ASAP7_75t_SL \i58/i209  (.A1(\i58/n62 ),
    .A2(\i58/n155 ),
    .B1(\i58/n6 ),
    .B2(\i58/n551 ),
    .Y(\i58/n274 ));
 AND4x1_ASAP7_75t_SL \i58/i21  (.A(\i58/n443 ),
    .B(\i58/n449 ),
    .C(\i58/n431 ),
    .D(\i58/n416 ),
    .Y(\i58/n465 ));
 OAI22xp5_ASAP7_75t_SL \i58/i210  (.A1(\i58/n57 ),
    .A2(\i58/n148 ),
    .B1(\i58/n53 ),
    .B2(\i58/n69 ),
    .Y(\i58/n273 ));
 AOI221xp5_ASAP7_75t_SL \i58/i211  (.A1(\i58/n46 ),
    .A2(\i58/n532 ),
    .B1(\i58/n42 ),
    .B2(\i58/n41 ),
    .C(\i58/n233 ),
    .Y(\i58/n272 ));
 AND4x1_ASAP7_75t_SL \i58/i212  (.A(\i58/n127 ),
    .B(\i58/n9 ),
    .C(\i58/n13 ),
    .D(\i58/n133 ),
    .Y(\i58/n271 ));
 NAND4xp25_ASAP7_75t_SL \i58/i213  (.A(\i58/n122 ),
    .B(\i58/n505 ),
    .C(\i58/n110 ),
    .D(\i58/n487 ),
    .Y(\i58/n270 ));
 NAND4xp25_ASAP7_75t_SL \i58/i214  (.A(\i58/n132 ),
    .B(\i58/n507 ),
    .C(\i58/n186 ),
    .D(\i58/n128 ),
    .Y(\i58/n269 ));
 AOI22xp5_ASAP7_75t_SL \i58/i215  (.A1(\i58/n520 ),
    .A2(\i58/n97 ),
    .B1(\i58/n75 ),
    .B2(\i58/n111 ),
    .Y(\i58/n268 ));
 OAI211xp5_ASAP7_75t_SL \i58/i216  (.A1(\i58/n67 ),
    .A2(\i58/n177 ),
    .B(\i58/n88 ),
    .C(\i58/n135 ),
    .Y(\i58/n267 ));
 NAND4xp25_ASAP7_75t_SL \i58/i217  (.A(\i58/n13 ),
    .B(\i58/n149 ),
    .C(\i58/n161 ),
    .D(\i58/n550 ),
    .Y(\i58/n266 ));
 OAI22xp5_ASAP7_75t_SL \i58/i218  (.A1(\i58/n78 ),
    .A2(\i58/n152 ),
    .B1(\i58/n6 ),
    .B2(\i58/n112 ),
    .Y(\i58/n265 ));
 OAI22xp5_ASAP7_75t_SL \i58/i219  (.A1(\i58/n2 ),
    .A2(\i58/n497 ),
    .B1(\i58/n72 ),
    .B2(\i58/n40 ),
    .Y(\i58/n264 ));
 NAND3xp33_ASAP7_75t_SL \i58/i22  (.A(\i58/n401 ),
    .B(\i58/n376 ),
    .C(\i58/n398 ),
    .Y(\i58/n463 ));
 AOI211x1_ASAP7_75t_SL \i58/i220  (.A1(\i58/n162 ),
    .A2(\i58/n85 ),
    .B(\i58/n181 ),
    .C(\i58/n179 ),
    .Y(\i58/n263 ));
 NAND4xp25_ASAP7_75t_SL \i58/i221  (.A(\i58/n169 ),
    .B(\i58/n554 ),
    .C(\i58/n490 ),
    .D(\i58/n124 ),
    .Y(\i58/n262 ));
 OAI22xp5_ASAP7_75t_SL \i58/i222  (.A1(\i58/n498 ),
    .A2(\i58/n95 ),
    .B1(\i58/n80 ),
    .B2(\i58/n6 ),
    .Y(\i58/n261 ));
 AOI222xp33_ASAP7_75t_SL \i58/i223  (.A1(\i58/n56 ),
    .A2(\i58/n94 ),
    .B1(\i58/n534 ),
    .B2(\i58/n77 ),
    .C1(\i58/n66 ),
    .C2(\i58/n41 ),
    .Y(\i58/n260 ));
 OAI221xp5_ASAP7_75t_R \i58/i224  (.A1(\i58/n489 ),
    .A2(\i58/n76 ),
    .B1(\i58/n69 ),
    .B2(\i58/n84 ),
    .C(\i58/n153 ),
    .Y(\i58/n259 ));
 OAI221xp5_ASAP7_75t_SL \i58/i225  (.A1(\i58/n498 ),
    .A2(\i58/n78 ),
    .B1(\i58/n76 ),
    .B2(\i58/n45 ),
    .C(\i58/n144 ),
    .Y(\i58/n258 ));
 OAI221xp5_ASAP7_75t_SL \i58/i226  (.A1(\i58/n10 ),
    .A2(\i58/n40 ),
    .B1(\i58/n2 ),
    .B2(\i58/n55 ),
    .C(\i58/n492 ),
    .Y(\i58/n257 ));
 OAI211xp5_ASAP7_75t_SL \i58/i227  (.A1(\i58/n55 ),
    .A2(\i58/n134 ),
    .B(\i58/n130 ),
    .C(\i58/n92 ),
    .Y(\i58/n256 ));
 AOI221xp5_ASAP7_75t_SL \i58/i228  (.A1(\i58/n192 ),
    .A2(\i58/n59 ),
    .B1(\i58/n83 ),
    .B2(\i58/n534 ),
    .C(\i58/n123 ),
    .Y(\i58/n255 ));
 AOI22xp33_ASAP7_75t_SL \i58/i229  (.A1(\i58/n50 ),
    .A2(\i58/n192 ),
    .B1(\i58/n70 ),
    .B2(\i58/n511 ),
    .Y(\i58/n254 ));
 NOR2xp33_ASAP7_75t_SL \i58/i23  (.A(\i58/n435 ),
    .B(\i58/n432 ),
    .Y(\i58/n462 ));
 OAI221xp5_ASAP7_75t_SL \i58/i230  (.A1(\i58/n498 ),
    .A2(\i58/n69 ),
    .B1(\i58/n65 ),
    .B2(\i58/n82 ),
    .C(\i58/n552 ),
    .Y(\i58/n292 ));
 OAI221xp5_ASAP7_75t_SL \i58/i231  (.A1(\i58/n49 ),
    .A2(\i58/n43 ),
    .B1(\i58/n78 ),
    .B2(\i58/n514 ),
    .C(\i58/n100 ),
    .Y(\i58/n290 ));
 OAI21xp5_ASAP7_75t_L \i58/i232  (.A1(\i58/n180 ),
    .A2(\i58/n514 ),
    .B(\i58/n106 ),
    .Y(\i58/n287 ));
 AOI221x1_ASAP7_75t_SL \i58/i233  (.A1(\i58/n1 ),
    .A2(\i58/n511 ),
    .B1(\i58/n71 ),
    .B2(\i58/n158 ),
    .C(\i58/n150 ),
    .Y(\i58/n285 ));
 OAI221xp5_ASAP7_75t_SL \i58/i234  (.A1(\i58/n151 ),
    .A2(\i58/n546 ),
    .B1(\i58/n80 ),
    .B2(\i58/n45 ),
    .C(\i58/n173 ),
    .Y(\i58/n283 ));
 AOI22xp5_ASAP7_75t_SL \i58/i235  (.A1(\i58/n71 ),
    .A2(\i58/n163 ),
    .B1(\i58/n52 ),
    .B2(\i58/n73 ),
    .Y(\i58/n282 ));
 INVxp67_ASAP7_75t_SL \i58/i236  (.A(\i58/n250 ),
    .Y(\i58/n251 ));
 INVxp67_ASAP7_75t_SL \i58/i237  (.A(\i58/n542 ),
    .Y(\i58/n248 ));
 INVxp67_ASAP7_75t_SL \i58/i238  (.A(\i58/n246 ),
    .Y(\i58/n247 ));
 INVx1_ASAP7_75t_SL \i58/i239  (.A(\i58/n243 ),
    .Y(\i58/n244 ));
 NAND2xp33_ASAP7_75t_SL \i58/i24  (.A(\i58/n437 ),
    .B(\i58/n426 ),
    .Y(\i58/n461 ));
 INVxp67_ASAP7_75t_SL \i58/i240  (.A(\i58/n241 ),
    .Y(\i58/n242 ));
 INVxp67_ASAP7_75t_SL \i58/i241  (.A(\i58/n503 ),
    .Y(\i58/n238 ));
 NOR2xp33_ASAP7_75t_SL \i58/i242  (.A(\i58/n530 ),
    .B(\i58/n167 ),
    .Y(\i58/n237 ));
 OAI21xp5_ASAP7_75t_SL \i58/i243  (.A1(\i58/n48 ),
    .A2(\i58/n44 ),
    .B(\i58/n79 ),
    .Y(\i58/n236 ));
 AOI22xp5_ASAP7_75t_SL \i58/i244  (.A1(\i58/n50 ),
    .A2(\i58/n511 ),
    .B1(\i58/n83 ),
    .B2(\i58/n56 ),
    .Y(\i58/n235 ));
 OAI21xp5_ASAP7_75t_SL \i58/i245  (.A1(\i58/n546 ),
    .A2(\i58/n43 ),
    .B(\i58/n135 ),
    .Y(\i58/n234 ));
 AOI21xp33_ASAP7_75t_SL \i58/i246  (.A1(\i58/n64 ),
    .A2(\i58/n514 ),
    .B(\i58/n164 ),
    .Y(\i58/n233 ));
 OAI21xp5_ASAP7_75t_SL \i58/i247  (.A1(\i58/n2 ),
    .A2(\i58/n62 ),
    .B(\i58/n174 ),
    .Y(\i58/n253 ));
 NAND2xp5_ASAP7_75t_L \i58/i248  (.A(\i58/n136 ),
    .B(\i58/n145 ),
    .Y(\i58/n232 ));
 OAI21xp33_ASAP7_75t_SL \i58/i249  (.A1(\i58/n58 ),
    .A2(\i58/n62 ),
    .B(\i58/n186 ),
    .Y(\i58/n231 ));
 NOR2xp33_ASAP7_75t_SL \i58/i25  (.A(\i58/n415 ),
    .B(\i58/n440 ),
    .Y(\i58/n460 ));
 AOI21xp5_ASAP7_75t_SL \i58/i250  (.A1(\i58/n5 ),
    .A2(\i58/n72 ),
    .B(\i58/n78 ),
    .Y(\i58/n252 ));
 AOI21xp33_ASAP7_75t_SL \i58/i251  (.A1(\i58/n72 ),
    .A2(\i58/n479 ),
    .B(\i58/n164 ),
    .Y(\i58/n230 ));
 AOI22xp5_ASAP7_75t_SL \i58/i252  (.A1(\i58/n531 ),
    .A2(\i58/n81 ),
    .B1(\i58/n77 ),
    .B2(\i58/n73 ),
    .Y(\i58/n229 ));
 OAI21xp33_ASAP7_75t_SL \i58/i253  (.A1(\i58/n57 ),
    .A2(\i58/n62 ),
    .B(\i58/n129 ),
    .Y(\i58/n228 ));
 NOR2xp33_ASAP7_75t_SL \i58/i254  (.A(\i58/n141 ),
    .B(\i58/n170 ),
    .Y(\i58/n227 ));
 OAI22xp5_ASAP7_75t_SL \i58/i255  (.A1(\i58/n82 ),
    .A2(\i58/n514 ),
    .B1(\i58/n74 ),
    .B2(\i58/n5 ),
    .Y(\i58/n226 ));
 OAI21xp5_ASAP7_75t_SL \i58/i256  (.A1(\i58/n53 ),
    .A2(\i58/n51 ),
    .B(\i58/n185 ),
    .Y(\i58/n225 ));
 OAI21xp5_ASAP7_75t_SL \i58/i257  (.A1(\i58/n53 ),
    .A2(\i58/n57 ),
    .B(\i58/n9 ),
    .Y(\i58/n250 ));
 OAI21xp5_ASAP7_75t_SL \i58/i258  (.A1(\i58/n80 ),
    .A2(\i58/n498 ),
    .B(\i58/n189 ),
    .Y(\i58/n249 ));
 OAI22xp5_ASAP7_75t_SL \i58/i259  (.A1(\i58/n64 ),
    .A2(\i58/n58 ),
    .B1(\i58/n76 ),
    .B2(\i58/n498 ),
    .Y(\i58/n246 ));
 NOR2xp33_ASAP7_75t_SL \i58/i26  (.A(\i58/n448 ),
    .B(\i58/n442 ),
    .Y(\i58/n459 ));
 AOI22xp5_ASAP7_75t_SL \i58/i260  (.A1(\i58/n71 ),
    .A2(\i58/n59 ),
    .B1(\i58/n70 ),
    .B2(\i58/n73 ),
    .Y(\i58/n245 ));
 OAI22xp5_ASAP7_75t_SL \i58/i261  (.A1(\i58/n54 ),
    .A2(\i58/n514 ),
    .B1(\i58/n67 ),
    .B2(\i58/n6 ),
    .Y(\i58/n224 ));
 OAI21xp5_ASAP7_75t_SL \i58/i262  (.A1(\i58/n53 ),
    .A2(\i58/n40 ),
    .B(\i58/n14 ),
    .Y(\i58/n243 ));
 NAND2xp5_ASAP7_75t_SL \i58/i263  (.A(\i58/n44 ),
    .B(\i58/n8 ),
    .Y(\i58/n241 ));
 NAND2xp5_ASAP7_75t_SL \i58/i264  (.A(\i58/n81 ),
    .B(\i58/n11 ),
    .Y(\i58/n240 ));
 NAND2xp5_ASAP7_75t_SL \i58/i265  (.A(\i58/n85 ),
    .B(\i58/n163 ),
    .Y(\i58/n239 ));
 INVxp67_ASAP7_75t_SL \i58/i266  (.A(\i58/n222 ),
    .Y(\i58/n223 ));
 INVxp67_ASAP7_75t_SL \i58/i267  (.A(\i58/n528 ),
    .Y(\i58/n216 ));
 INVxp67_ASAP7_75t_SL \i58/i268  (.A(\i58/n214 ),
    .Y(\i58/n215 ));
 INVx1_ASAP7_75t_SL \i58/i269  (.A(\i58/n209 ),
    .Y(\i58/n210 ));
 AND2x2_ASAP7_75t_SL \i58/i27  (.A(\i58/n406 ),
    .B(\i58/n439 ),
    .Y(\i58/n464 ));
 OAI21xp5_ASAP7_75t_SL \i58/i270  (.A1(\i58/n44 ),
    .A2(\i58/n42 ),
    .B(\i58/n52 ),
    .Y(\i58/n206 ));
 AOI21xp33_ASAP7_75t_SL \i58/i271  (.A1(\i58/n62 ),
    .A2(\i58/n72 ),
    .B(\i58/n40 ),
    .Y(\i58/n205 ));
 AOI22xp5_ASAP7_75t_SL \i58/i272  (.A1(\i58/n85 ),
    .A2(\i58/n532 ),
    .B1(\i58/n50 ),
    .B2(\i58/n66 ),
    .Y(\i58/n204 ));
 AOI22xp5_ASAP7_75t_SL \i58/i273  (.A1(\i58/n56 ),
    .A2(\i58/n59 ),
    .B1(\i58/n73 ),
    .B2(\i58/n520 ),
    .Y(\i58/n203 ));
 AOI22xp5_ASAP7_75t_SL \i58/i274  (.A1(\i58/n85 ),
    .A2(\i58/n59 ),
    .B1(\i58/n81 ),
    .B2(\i58/n44 ),
    .Y(\i58/n222 ));
 OAI22xp5_ASAP7_75t_SL \i58/i275  (.A1(\i58/n40 ),
    .A2(\i58/n62 ),
    .B1(\i58/n60 ),
    .B2(\i58/n58 ),
    .Y(\i58/n202 ));
 OAI22xp5_ASAP7_75t_SL \i58/i276  (.A1(\i58/n76 ),
    .A2(\i58/n55 ),
    .B1(\i58/n53 ),
    .B2(\i58/n78 ),
    .Y(\i58/n201 ));
 OAI21xp5_ASAP7_75t_SL \i58/i277  (.A1(\i58/n82 ),
    .A2(\i58/n5 ),
    .B(\i58/n114 ),
    .Y(\i58/n200 ));
 AOI22xp5_ASAP7_75t_SL \i58/i278  (.A1(\i58/n520 ),
    .A2(\i58/n534 ),
    .B1(\i58/n41 ),
    .B2(\i58/n48 ),
    .Y(\i58/n199 ));
 OAI22xp5_ASAP7_75t_SL \i58/i279  (.A1(\i58/n84 ),
    .A2(\i58/n82 ),
    .B1(\i58/n43 ),
    .B2(\i58/n58 ),
    .Y(\i58/n221 ));
 NOR2xp33_ASAP7_75t_SL \i58/i28  (.A(\i58/n447 ),
    .B(\i58/n429 ),
    .Y(\i58/n457 ));
 OAI22xp5_ASAP7_75t_SL \i58/i280  (.A1(\i58/n69 ),
    .A2(\i58/n62 ),
    .B1(\i58/n40 ),
    .B2(\i58/n64 ),
    .Y(\i58/n220 ));
 NAND2xp5_ASAP7_75t_SL \i58/i281  (.A(\i58/n194 ),
    .B(\i58/n12 ),
    .Y(\i58/n198 ));
 AOI22xp5_ASAP7_75t_SL \i58/i282  (.A1(\i58/n50 ),
    .A2(\i58/n63 ),
    .B1(\i58/n48 ),
    .B2(\i58/n1 ),
    .Y(\i58/n219 ));
 NAND2xp5_ASAP7_75t_SL \i58/i283  (.A(\i58/n193 ),
    .B(\i58/n140 ),
    .Y(\i58/n197 ));
 OAI22xp5_ASAP7_75t_SL \i58/i284  (.A1(\i58/n53 ),
    .A2(\i58/n82 ),
    .B1(\i58/n67 ),
    .B2(\i58/n65 ),
    .Y(\i58/n218 ));
 OAI22xp33_ASAP7_75t_SL \i58/i285  (.A1(\i58/n78 ),
    .A2(\i58/n479 ),
    .B1(\i58/n60 ),
    .B2(\i58/n67 ),
    .Y(\i58/n196 ));
 OAI22xp5_ASAP7_75t_SL \i58/i286  (.A1(\i58/n62 ),
    .A2(\i58/n67 ),
    .B1(\i58/n43 ),
    .B2(\i58/n40 ),
    .Y(\i58/n217 ));
 AOI22xp5_ASAP7_75t_SL \i58/i287  (.A1(\i58/n63 ),
    .A2(\i58/n83 ),
    .B1(\i58/n85 ),
    .B2(\i58/n75 ),
    .Y(\i58/n214 ));
 OAI22xp5_ASAP7_75t_SL \i58/i288  (.A1(\i58/n76 ),
    .A2(\i58/n5 ),
    .B1(\i58/n65 ),
    .B2(\i58/n54 ),
    .Y(\i58/n213 ));
 OAI22xp5_ASAP7_75t_SL \i58/i289  (.A1(\i58/n479 ),
    .A2(\i58/n49 ),
    .B1(\i58/n6 ),
    .B2(\i58/n40 ),
    .Y(\i58/n212 ));
 NOR2xp33_ASAP7_75t_SL \i58/i29  (.A(\i58/n428 ),
    .B(\i58/n423 ),
    .Y(\i58/n456 ));
 OAI22x1_ASAP7_75t_SL \i58/i290  (.A1(\i58/n2 ),
    .A2(\i58/n514 ),
    .B1(\i58/n47 ),
    .B2(\i58/n78 ),
    .Y(\i58/n211 ));
 AO22x1_ASAP7_75t_SL \i58/i291  (.A1(\i58/n52 ),
    .A2(\i58/n63 ),
    .B1(\i58/n73 ),
    .B2(\i58/n83 ),
    .Y(\i58/n209 ));
 AOI22xp5_ASAP7_75t_SL \i58/i292  (.A1(\i58/n42 ),
    .A2(\i58/n59 ),
    .B1(\i58/n75 ),
    .B2(\i58/n73 ),
    .Y(\i58/n208 ));
 AOI22xp5_ASAP7_75t_SL \i58/i293  (.A1(\i58/n534 ),
    .A2(\i58/n79 ),
    .B1(\i58/n68 ),
    .B2(\i58/n56 ),
    .Y(\i58/n207 ));
 INVxp67_ASAP7_75t_SL \i58/i294  (.A(\i58/n12 ),
    .Y(\i58/n191 ));
 INVxp67_ASAP7_75t_SL \i58/i295  (.A(\i58/n187 ),
    .Y(\i58/n188 ));
 INVxp67_ASAP7_75t_SL \i58/i296  (.A(\i58/n554 ),
    .Y(\i58/n184 ));
 INVxp67_ASAP7_75t_SL \i58/i297  (.A(\i58/n530 ),
    .Y(\i58/n183 ));
 INVxp67_ASAP7_75t_SL \i58/i298  (.A(\i58/n181 ),
    .Y(\i58/n182 ));
 INVxp67_ASAP7_75t_SL \i58/i299  (.A(\i58/n486 ),
    .Y(\i58/n175 ));
 AND3x2_ASAP7_75t_SL \i58/i3  (.A(\i58/n462 ),
    .B(\i58/n475 ),
    .C(\i58/n458 ),
    .Y(n4[6]));
 NOR2xp33_ASAP7_75t_SL \i58/i30  (.A(\i58/n422 ),
    .B(\i58/n441 ),
    .Y(\i58/n455 ));
 INVx1_ASAP7_75t_SL \i58/i300  (.A(\i58/n171 ),
    .Y(\i58/n172 ));
 INVxp67_ASAP7_75t_SL \i58/i301  (.A(\i58/n169 ),
    .Y(\i58/n170 ));
 INVxp67_ASAP7_75t_SL \i58/i302  (.A(\i58/n167 ),
    .Y(\i58/n168 ));
 INVx1_ASAP7_75t_SL \i58/i303  (.A(\i58/n165 ),
    .Y(\i58/n166 ));
 NAND2xp5_ASAP7_75t_L \i58/i304  (.A(\i58/n80 ),
    .B(\i58/n69 ),
    .Y(\i58/n162 ));
 NAND2xp5_ASAP7_75t_SL \i58/i305  (.A(\i58/n532 ),
    .B(\i58/n42 ),
    .Y(\i58/n161 ));
 NAND2xp33_ASAP7_75t_L \i58/i306  (.A(\i58/n82 ),
    .B(\i58/n74 ),
    .Y(\i58/n160 ));
 NOR2xp33_ASAP7_75t_L \i58/i307  (.A(\i58/n48 ),
    .B(\i58/n61 ),
    .Y(\i58/n159 ));
 AND2x2_ASAP7_75t_SL \i58/i308  (.A(\i58/n44 ),
    .B(\i58/n83 ),
    .Y(\i58/n195 ));
 NAND2xp5_ASAP7_75t_SL \i58/i309  (.A(\i58/n51 ),
    .B(\i58/n2 ),
    .Y(\i58/n158 ));
 AND4x1_ASAP7_75t_SL \i58/i31  (.A(\i58/n411 ),
    .B(\i58/n407 ),
    .C(\i58/n368 ),
    .D(\i58/n361 ),
    .Y(\i58/n454 ));
 NAND2xp5_ASAP7_75t_SL \i58/i310  (.A(\i58/n58 ),
    .B(\i58/n2 ),
    .Y(\i58/n157 ));
 NAND2xp5_ASAP7_75t_SL \i58/i311  (.A(\i58/n66 ),
    .B(\i58/n532 ),
    .Y(\i58/n156 ));
 NOR2xp33_ASAP7_75t_SL \i58/i312  (.A(\i58/n75 ),
    .B(\i58/n79 ),
    .Y(\i58/n155 ));
 NAND2xp5_ASAP7_75t_SL \i58/i313  (.A(\i58/n46 ),
    .B(\i58/n83 ),
    .Y(\i58/n194 ));
 NAND2xp5_ASAP7_75t_SL \i58/i314  (.A(\i58/n56 ),
    .B(\i58/n520 ),
    .Y(\i58/n154 ));
 NAND2xp5_ASAP7_75t_SL \i58/i315  (.A(\i58/n61 ),
    .B(\i58/n52 ),
    .Y(\i58/n153 ));
 NOR2xp33_ASAP7_75t_SL \i58/i316  (.A(\i58/n531 ),
    .B(\i58/n42 ),
    .Y(\i58/n152 ));
 NOR2xp33_ASAP7_75t_SL \i58/i317  (.A(\i58/n63 ),
    .B(\i58/n48 ),
    .Y(\i58/n151 ));
 NOR2xp67_ASAP7_75t_SL \i58/i318  (.A(\i58/n76 ),
    .B(\i58/n65 ),
    .Y(\i58/n150 ));
 NAND2xp5_ASAP7_75t_SL \i58/i319  (.A(\i58/n79 ),
    .B(\i58/n46 ),
    .Y(\i58/n149 ));
 NOR3xp33_ASAP7_75t_SL \i58/i32  (.A(\i58/n404 ),
    .B(\i58/n336 ),
    .C(\i58/n392 ),
    .Y(\i58/n453 ));
 NOR2xp33_ASAP7_75t_SL \i58/i320  (.A(\i58/n63 ),
    .B(\i58/n66 ),
    .Y(\i58/n148 ));
 NOR2xp33_ASAP7_75t_SL \i58/i321  (.A(\i58/n44 ),
    .B(\i58/n63 ),
    .Y(\i58/n147 ));
 NOR2xp33_ASAP7_75t_SL \i58/i322  (.A(\i58/n71 ),
    .B(\i58/n66 ),
    .Y(\i58/n146 ));
 NAND2xp5_ASAP7_75t_SL \i58/i323  (.A(\i58/n68 ),
    .B(\i58/n48 ),
    .Y(\i58/n193 ));
 NAND2xp5_ASAP7_75t_SL \i58/i324  (.A(\i58/n73 ),
    .B(\i58/n59 ),
    .Y(\i58/n145 ));
 NAND2xp5_ASAP7_75t_SL \i58/i325  (.A(\i58/n531 ),
    .B(\i58/n68 ),
    .Y(\i58/n144 ));
 NAND2xp5_ASAP7_75t_SL \i58/i326  (.A(\i58/n61 ),
    .B(\i58/n532 ),
    .Y(\i58/n16 ));
 NOR2xp33_ASAP7_75t_SL \i58/i327  (.A(\i58/n67 ),
    .B(\i58/n6 ),
    .Y(\i58/n143 ));
 NAND2xp5_ASAP7_75t_SL \i58/i328  (.A(\i58/n1 ),
    .B(\i58/n534 ),
    .Y(\i58/n15 ));
 NAND2xp33_ASAP7_75t_SL \i58/i329  (.A(\i58/n43 ),
    .B(\i58/n72 ),
    .Y(\i58/n192 ));
 NAND2xp33_ASAP7_75t_SL \i58/i33  (.A(\i58/n19 ),
    .B(\i58/n424 ),
    .Y(\i58/n452 ));
 NAND2xp5_ASAP7_75t_SL \i58/i330  (.A(\i58/n533 ),
    .B(\i58/n63 ),
    .Y(\i58/n14 ));
 NAND2xp5_ASAP7_75t_SL \i58/i331  (.A(\i58/n73 ),
    .B(\i58/n1 ),
    .Y(\i58/n13 ));
 NOR2xp33_ASAP7_75t_SL \i58/i332  (.A(\i58/n72 ),
    .B(\i58/n69 ),
    .Y(\i58/n142 ));
 NAND2xp5_ASAP7_75t_SL \i58/i333  (.A(\i58/n77 ),
    .B(\i58/n63 ),
    .Y(\i58/n12 ));
 NAND2xp5_ASAP7_75t_SL \i58/i334  (.A(\i58/n85 ),
    .B(\i58/n77 ),
    .Y(\i58/n190 ));
 NAND2xp5_ASAP7_75t_SL \i58/i335  (.A(\i58/n85 ),
    .B(\i58/n533 ),
    .Y(\i58/n189 ));
 NAND2xp5_ASAP7_75t_L \i58/i336  (.A(\i58/n79 ),
    .B(\i58/n85 ),
    .Y(\i58/n187 ));
 NAND2xp5_ASAP7_75t_SL \i58/i337  (.A(\i58/n71 ),
    .B(\i58/n77 ),
    .Y(\i58/n186 ));
 NAND2xp5_ASAP7_75t_SL \i58/i338  (.A(\i58/n75 ),
    .B(\i58/n71 ),
    .Y(\i58/n185 ));
 AND2x2_ASAP7_75t_SL \i58/i339  (.A(\i58/n83 ),
    .B(\i58/n71 ),
    .Y(\i58/n181 ));
 AND3x1_ASAP7_75t_SL \i58/i34  (.A(\i58/n410 ),
    .B(\i58/n3 ),
    .C(\i58/n403 ),
    .Y(\i58/n458 ));
 NOR2x1_ASAP7_75t_SL \i58/i340  (.A(\i58/n68 ),
    .B(\i58/n52 ),
    .Y(\i58/n180 ));
 AND2x2_ASAP7_75t_SL \i58/i341  (.A(\i58/n520 ),
    .B(\i58/n66 ),
    .Y(\i58/n179 ));
 NAND2xp5_ASAP7_75t_SL \i58/i342  (.A(\i58/n68 ),
    .B(\i58/n46 ),
    .Y(\i58/n178 ));
 NOR2xp33_ASAP7_75t_L \i58/i343  (.A(\i58/n44 ),
    .B(\i58/n61 ),
    .Y(\i58/n177 ));
 NAND2xp5_ASAP7_75t_SL \i58/i344  (.A(\i58/n73 ),
    .B(\i58/n532 ),
    .Y(\i58/n176 ));
 NAND2xp5_ASAP7_75t_SL \i58/i345  (.A(\i58/n61 ),
    .B(\i58/n41 ),
    .Y(\i58/n174 ));
 NAND2xp5_ASAP7_75t_SL \i58/i346  (.A(\i58/n61 ),
    .B(\i58/n79 ),
    .Y(\i58/n173 ));
 NOR2xp33_ASAP7_75t_SL \i58/i347  (.A(\i58/n49 ),
    .B(\i58/n60 ),
    .Y(\i58/n141 ));
 NOR2xp33_ASAP7_75t_L \i58/i348  (.A(\i58/n41 ),
    .B(\i58/n68 ),
    .Y(\i58/n171 ));
 NAND2xp5_ASAP7_75t_SL \i58/i349  (.A(\i58/n85 ),
    .B(\i58/n1 ),
    .Y(\i58/n169 ));
 INVxp67_ASAP7_75t_SL \i58/i35  (.A(\i58/n450 ),
    .Y(\i58/n451 ));
 NAND2xp5_ASAP7_75t_L \i58/i350  (.A(\i58/n2 ),
    .B(\i58/n74 ),
    .Y(\i58/n167 ));
 NOR2xp33_ASAP7_75t_L \i58/i351  (.A(\i58/n81 ),
    .B(\i58/n75 ),
    .Y(\i58/n165 ));
 NOR2xp33_ASAP7_75t_L \i58/i352  (.A(\i58/n81 ),
    .B(\i58/n68 ),
    .Y(\i58/n164 ));
 NAND2xp5_ASAP7_75t_SL \i58/i353  (.A(\i58/n49 ),
    .B(\i58/n546 ),
    .Y(\i58/n163 ));
 NAND2xp67_ASAP7_75t_SL \i58/i354  (.A(\i58/n5 ),
    .B(\i58/n60 ),
    .Y(\i58/n11 ));
 INVxp67_ASAP7_75t_SL \i58/i355  (.A(\i58/n136 ),
    .Y(\i58/n137 ));
 INVxp67_ASAP7_75t_SL \i58/i356  (.A(\i58/n130 ),
    .Y(\i58/n131 ));
 INVxp67_ASAP7_75t_SL \i58/i357  (.A(\i58/n125 ),
    .Y(\i58/n126 ));
 INVxp67_ASAP7_75t_SL \i58/i358  (.A(\i58/n122 ),
    .Y(\i58/n123 ));
 INVxp67_ASAP7_75t_SL \i58/i359  (.A(\i58/n7 ),
    .Y(\i58/n119 ));
 INVxp67_ASAP7_75t_SL \i58/i36  (.A(\i58/n448 ),
    .Y(\i58/n449 ));
 NOR2xp33_ASAP7_75t_SL \i58/i360  (.A(\i58/n44 ),
    .B(\i58/n56 ),
    .Y(\i58/n118 ));
 NOR2xp33_ASAP7_75t_SL \i58/i361  (.A(\i58/n80 ),
    .B(\i58/n47 ),
    .Y(\i58/n117 ));
 NAND2xp33_ASAP7_75t_SL \i58/i362  (.A(\i58/n54 ),
    .B(\i58/n74 ),
    .Y(\i58/n116 ));
 NOR2xp33_ASAP7_75t_R \i58/i363  (.A(\i58/n77 ),
    .B(\i58/n1 ),
    .Y(\i58/n115 ));
 NAND2xp5_ASAP7_75t_SL \i58/i364  (.A(\i58/n44 ),
    .B(\i58/n79 ),
    .Y(\i58/n114 ));
 NAND2xp5_ASAP7_75t_SL \i58/i365  (.A(\i58/n81 ),
    .B(\i58/n42 ),
    .Y(\i58/n113 ));
 NOR2xp33_ASAP7_75t_SL \i58/i366  (.A(\i58/n81 ),
    .B(\i58/n52 ),
    .Y(\i58/n112 ));
 NAND2xp33_ASAP7_75t_L \i58/i367  (.A(\i58/n514 ),
    .B(\i58/n55 ),
    .Y(\i58/n111 ));
 NAND2xp5_ASAP7_75t_SL \i58/i368  (.A(\i58/n70 ),
    .B(\i58/n71 ),
    .Y(\i58/n110 ));
 NAND2xp33_ASAP7_75t_SL \i58/i369  (.A(\i58/n57 ),
    .B(\i58/n54 ),
    .Y(\i58/n109 ));
 NAND3xp33_ASAP7_75t_SL \i58/i37  (.A(\i58/n400 ),
    .B(\i58/n352 ),
    .C(\i58/n360 ),
    .Y(\i58/n446 ));
 NOR2xp33_ASAP7_75t_SL \i58/i370  (.A(\i58/n1 ),
    .B(\i58/n41 ),
    .Y(\i58/n108 ));
 NAND2xp5_ASAP7_75t_SL \i58/i371  (.A(\i58/n71 ),
    .B(\i58/n533 ),
    .Y(\i58/n107 ));
 NAND2xp5_ASAP7_75t_SL \i58/i372  (.A(\i58/n1 ),
    .B(\i58/n56 ),
    .Y(\i58/n106 ));
 NAND2xp33_ASAP7_75t_SL \i58/i373  (.A(\i58/n43 ),
    .B(\i58/n64 ),
    .Y(\i58/n105 ));
 NAND2xp33_ASAP7_75t_SL \i58/i374  (.A(\i58/n69 ),
    .B(\i58/n65 ),
    .Y(\i58/n104 ));
 NOR2xp33_ASAP7_75t_SL \i58/i375  (.A(\i58/n46 ),
    .B(\i58/n534 ),
    .Y(\i58/n103 ));
 NAND2xp33_ASAP7_75t_L \i58/i376  (.A(\i58/n45 ),
    .B(\i58/n53 ),
    .Y(\i58/n102 ));
 NAND2xp5_ASAP7_75t_SL \i58/i377  (.A(\i58/n46 ),
    .B(\i58/n59 ),
    .Y(\i58/n140 ));
 NAND2xp33_ASAP7_75t_SL \i58/i378  (.A(\i58/n47 ),
    .B(\i58/n45 ),
    .Y(\i58/n101 ));
 NAND2xp5_ASAP7_75t_SL \i58/i379  (.A(\i58/n52 ),
    .B(\i58/n66 ),
    .Y(\i58/n100 ));
 NAND3xp33_ASAP7_75t_SL \i58/i38  (.A(\i58/n353 ),
    .B(\i58/n339 ),
    .C(\i58/n316 ),
    .Y(\i58/n445 ));
 NAND2xp5_ASAP7_75t_SL \i58/i380  (.A(\i58/n46 ),
    .B(\i58/n50 ),
    .Y(\i58/n139 ));
 NOR2xp33_ASAP7_75t_SL \i58/i381  (.A(\i58/n49 ),
    .B(\i58/n64 ),
    .Y(\i58/n99 ));
 NOR2xp33_ASAP7_75t_SL \i58/i382  (.A(\i58/n56 ),
    .B(\i58/n42 ),
    .Y(\i58/n98 ));
 NAND2xp33_ASAP7_75t_SL \i58/i383  (.A(\i58/n47 ),
    .B(\i58/n498 ),
    .Y(\i58/n97 ));
 NAND2xp5_ASAP7_75t_SL \i58/i384  (.A(\i58/n533 ),
    .B(\i58/n48 ),
    .Y(\i58/n96 ));
 NOR2xp33_ASAP7_75t_SL \i58/i385  (.A(\i58/n533 ),
    .B(\i58/n41 ),
    .Y(\i58/n95 ));
 NAND2xp5_ASAP7_75t_L \i58/i386  (.A(\i58/n54 ),
    .B(\i58/n69 ),
    .Y(\i58/n94 ));
 NOR2xp33_ASAP7_75t_SL \i58/i387  (.A(\i58/n71 ),
    .B(\i58/n534 ),
    .Y(\i58/n10 ));
 NAND2xp5_ASAP7_75t_SL \i58/i388  (.A(\i58/n52 ),
    .B(\i58/n534 ),
    .Y(\i58/n138 ));
 NOR2xp33_ASAP7_75t_SL \i58/i389  (.A(\i58/n54 ),
    .B(\i58/n64 ),
    .Y(\i58/n93 ));
 NAND2xp5_ASAP7_75t_L \i58/i39  (.A(\i58/n558 ),
    .B(\i58/n380 ),
    .Y(\i58/n444 ));
 NAND2xp5_ASAP7_75t_SL \i58/i390  (.A(\i58/n50 ),
    .B(\i58/n511 ),
    .Y(\i58/n92 ));
 NOR2xp33_ASAP7_75t_SL \i58/i391  (.A(\i58/n74 ),
    .B(\i58/n5 ),
    .Y(\i58/n91 ));
 NAND2xp5_ASAP7_75t_SL \i58/i392  (.A(\i58/n77 ),
    .B(\i58/n44 ),
    .Y(\i58/n136 ));
 NOR2xp33_ASAP7_75t_SL \i58/i393  (.A(\i58/n76 ),
    .B(\i58/n498 ),
    .Y(\i58/n90 ));
 NAND2xp5_ASAP7_75t_SL \i58/i394  (.A(\i58/n531 ),
    .B(\i58/n75 ),
    .Y(\i58/n135 ));
 NAND2xp5_ASAP7_75t_SL \i58/i395  (.A(\i58/n59 ),
    .B(\i58/n66 ),
    .Y(\i58/n9 ));
 NAND2x1p5_ASAP7_75t_SL \i58/i396  (.A(\i58/n74 ),
    .B(\i58/n69 ),
    .Y(\i58/n8 ));
 NOR2xp33_ASAP7_75t_L \i58/i397  (.A(\i58/n1 ),
    .B(\i58/n70 ),
    .Y(\i58/n134 ));
 NAND2xp5_ASAP7_75t_SL \i58/i398  (.A(\i58/n70 ),
    .B(\i58/n42 ),
    .Y(\i58/n133 ));
 NAND2xp5_ASAP7_75t_SL \i58/i399  (.A(\i58/n533 ),
    .B(\i58/n42 ),
    .Y(\i58/n132 ));
 AND2x4_ASAP7_75t_SL \i58/i4  (.A(\i58/n473 ),
    .B(\i58/n465 ),
    .Y(n4[3]));
 NOR2xp33_ASAP7_75t_SL \i58/i40  (.A(\i58/n408 ),
    .B(\i58/n334 ),
    .Y(\i58/n443 ));
 NOR2xp33_ASAP7_75t_SL \i58/i400  (.A(\i58/n53 ),
    .B(\i58/n58 ),
    .Y(\i58/n89 ));
 NAND2xp5_ASAP7_75t_SL \i58/i401  (.A(\i58/n531 ),
    .B(\i58/n81 ),
    .Y(\i58/n88 ));
 NAND2xp5_ASAP7_75t_SL \i58/i402  (.A(\i58/n41 ),
    .B(\i58/n511 ),
    .Y(\i58/n87 ));
 NAND2xp5_ASAP7_75t_SL \i58/i403  (.A(\i58/n50 ),
    .B(\i58/n48 ),
    .Y(\i58/n130 ));
 NAND2xp5_ASAP7_75t_SL \i58/i404  (.A(\i58/n59 ),
    .B(\i58/n48 ),
    .Y(\i58/n129 ));
 NOR2xp33_ASAP7_75t_SL \i58/i405  (.A(\i58/n47 ),
    .B(\i58/n51 ),
    .Y(\i58/n86 ));
 NAND2xp5_ASAP7_75t_SL \i58/i406  (.A(\i58/n41 ),
    .B(\i58/n56 ),
    .Y(\i58/n128 ));
 NAND2xp5_ASAP7_75t_SL \i58/i407  (.A(\i58/n52 ),
    .B(\i58/n56 ),
    .Y(\i58/n127 ));
 AND2x2_ASAP7_75t_SL \i58/i408  (.A(\i58/n533 ),
    .B(\i58/n44 ),
    .Y(\i58/n125 ));
 NAND4xp25_ASAP7_75t_SL \i58/i409  (.A(\i58/n509 ),
    .B(\i58/n495 ),
    .C(\i58/n29 ),
    .D(\i58/n30 ),
    .Y(\i58/n124 ));
 NAND2xp33_ASAP7_75t_L \i58/i41  (.A(\i58/n385 ),
    .B(\i58/n402 ),
    .Y(\i58/n442 ));
 NAND2xp5_ASAP7_75t_SL \i58/i410  (.A(\i58/n46 ),
    .B(\i58/n41 ),
    .Y(\i58/n122 ));
 AND2x2_ASAP7_75t_SL \i58/i411  (.A(\i58/n52 ),
    .B(\i58/n44 ),
    .Y(\i58/n121 ));
 AND2x2_ASAP7_75t_SL \i58/i412  (.A(\i58/n50 ),
    .B(\i58/n56 ),
    .Y(\i58/n120 ));
 NAND2xp5_ASAP7_75t_SL \i58/i413  (.A(\i58/n79 ),
    .B(\i58/n56 ),
    .Y(\i58/n7 ));
 INVx2_ASAP7_75t_SL \i58/i414  (.A(\i58/n85 ),
    .Y(\i58/n84 ));
 INVx2_ASAP7_75t_SL \i58/i415  (.A(\i58/n83 ),
    .Y(\i58/n82 ));
 INVx4_ASAP7_75t_SL \i58/i416  (.A(\i58/n81 ),
    .Y(\i58/n80 ));
 INVx3_ASAP7_75t_SL \i58/i417  (.A(\i58/n79 ),
    .Y(\i58/n78 ));
 INVx3_ASAP7_75t_SL \i58/i418  (.A(\i58/n77 ),
    .Y(\i58/n76 ));
 INVx3_ASAP7_75t_SL \i58/i419  (.A(\i58/n75 ),
    .Y(\i58/n74 ));
 NAND3xp33_ASAP7_75t_SL \i58/i42  (.A(\i58/n413 ),
    .B(\i58/n255 ),
    .C(\i58/n282 ),
    .Y(\i58/n441 ));
 INVx2_ASAP7_75t_SL \i58/i420  (.A(\i58/n73 ),
    .Y(\i58/n72 ));
 INVx3_ASAP7_75t_SL \i58/i421  (.A(\i58/n70 ),
    .Y(\i58/n69 ));
 INVx2_ASAP7_75t_SL \i58/i422  (.A(\i58/n68 ),
    .Y(\i58/n67 ));
 INVx2_ASAP7_75t_SL \i58/i423  (.A(\i58/n66 ),
    .Y(\i58/n65 ));
 INVx2_ASAP7_75t_SL \i58/i424  (.A(\i58/n534 ),
    .Y(\i58/n64 ));
 INVx3_ASAP7_75t_SL \i58/i425  (.A(\i58/n63 ),
    .Y(\i58/n62 ));
 AND2x4_ASAP7_75t_SL \i58/i426  (.A(\i58/n476 ),
    .B(\i58/n34 ),
    .Y(\i58/n85 ));
 AND2x4_ASAP7_75t_SL \i58/i427  (.A(\i58/n38 ),
    .B(\i58/n29 ),
    .Y(\i58/n83 ));
 AND2x4_ASAP7_75t_SL \i58/i428  (.A(\i58/n39 ),
    .B(\i58/n35 ),
    .Y(\i58/n81 ));
 AND2x4_ASAP7_75t_SL \i58/i429  (.A(\i58/n540 ),
    .B(\i58/n30 ),
    .Y(\i58/n79 ));
 NAND2xp33_ASAP7_75t_SL \i58/i43  (.A(\i58/n395 ),
    .B(\i58/n399 ),
    .Y(\i58/n440 ));
 AND2x4_ASAP7_75t_SL \i58/i430  (.A(\i58/n35 ),
    .B(\i58/n38 ),
    .Y(\i58/n77 ));
 AND2x4_ASAP7_75t_SL \i58/i431  (.A(\i58/n36 ),
    .B(\i58/n30 ),
    .Y(\i58/n75 ));
 AND2x4_ASAP7_75t_SL \i58/i432  (.A(\i58/n494 ),
    .B(\i58/n37 ),
    .Y(\i58/n73 ));
 AND2x2_ASAP7_75t_SL \i58/i433  (.A(\i58/n494 ),
    .B(\i58/n31 ),
    .Y(\i58/n71 ));
 NAND2x1_ASAP7_75t_SL \i58/i434  (.A(\i58/n494 ),
    .B(\i58/n31 ),
    .Y(\i58/n6 ));
 AND2x4_ASAP7_75t_SL \i58/i435  (.A(\i58/n35 ),
    .B(\i58/n539 ),
    .Y(\i58/n70 ));
 AND2x4_ASAP7_75t_SL \i58/i436  (.A(\i58/n35 ),
    .B(\i58/n30 ),
    .Y(\i58/n68 ));
 AND2x4_ASAP7_75t_SL \i58/i437  (.A(\i58/n494 ),
    .B(\i58/n510 ),
    .Y(\i58/n66 ));
 AND2x4_ASAP7_75t_SL \i58/i438  (.A(\i58/n509 ),
    .B(\i58/n495 ),
    .Y(\i58/n63 ));
 INVx2_ASAP7_75t_SL \i58/i439  (.A(\i58/n61 ),
    .Y(\i58/n60 ));
 NOR2xp33_ASAP7_75t_SL \i58/i44  (.A(\i58/n397 ),
    .B(\i58/n396 ),
    .Y(\i58/n439 ));
 INVx2_ASAP7_75t_SL \i58/i440  (.A(\i58/n59 ),
    .Y(\i58/n58 ));
 INVx2_ASAP7_75t_SL \i58/i441  (.A(\i58/n56 ),
    .Y(\i58/n55 ));
 INVx2_ASAP7_75t_SL \i58/i442  (.A(\i58/n52 ),
    .Y(\i58/n51 ));
 INVx3_ASAP7_75t_SL \i58/i443  (.A(\i58/n50 ),
    .Y(\i58/n49 ));
 INVx3_ASAP7_75t_SL \i58/i444  (.A(\i58/n48 ),
    .Y(\i58/n47 ));
 INVx4_ASAP7_75t_SL \i58/i445  (.A(\i58/n46 ),
    .Y(\i58/n45 ));
 INVx2_ASAP7_75t_SL \i58/i446  (.A(\i58/n44 ),
    .Y(\i58/n43 ));
 INVx5_ASAP7_75t_SL \i58/i447  (.A(\i58/n42 ),
    .Y(\i58/n5 ));
 INVx3_ASAP7_75t_SL \i58/i448  (.A(\i58/n41 ),
    .Y(\i58/n40 ));
 AND2x4_ASAP7_75t_SL \i58/i449  (.A(\i58/n27 ),
    .B(\i58/n37 ),
    .Y(\i58/n61 ));
 NAND4xp25_ASAP7_75t_SL \i58/i45  (.A(\i58/n375 ),
    .B(\i58/n311 ),
    .C(\i58/n238 ),
    .D(\i58/n275 ),
    .Y(\i58/n438 ));
 AND2x4_ASAP7_75t_SL \i58/i450  (.A(\i58/n30 ),
    .B(\i58/n29 ),
    .Y(\i58/n59 ));
 NAND2x1p5_ASAP7_75t_SL \i58/i451  (.A(\i58/n36 ),
    .B(\i58/n539 ),
    .Y(\i58/n57 ));
 AND2x4_ASAP7_75t_SL \i58/i452  (.A(\i58/n32 ),
    .B(\i58/n31 ),
    .Y(\i58/n56 ));
 NAND2xp5_ASAP7_75t_SL \i58/i453  (.A(\i58/n540 ),
    .B(\i58/n38 ),
    .Y(\i58/n54 ));
 OR2x6_ASAP7_75t_SL \i58/i454  (.A(\i58/n33 ),
    .B(\i58/n28 ),
    .Y(\i58/n53 ));
 AND2x4_ASAP7_75t_SL \i58/i455  (.A(\i58/n39 ),
    .B(\i58/n540 ),
    .Y(\i58/n52 ));
 AND2x4_ASAP7_75t_SL \i58/i456  (.A(\i58/n38 ),
    .B(\i58/n36 ),
    .Y(\i58/n50 ));
 AND2x4_ASAP7_75t_SL \i58/i457  (.A(\i58/n26 ),
    .B(\i58/n510 ),
    .Y(\i58/n48 ));
 AND2x4_ASAP7_75t_SL \i58/i458  (.A(\i58/n37 ),
    .B(\i58/n32 ),
    .Y(\i58/n46 ));
 AND2x4_ASAP7_75t_SL \i58/i459  (.A(\i58/n37 ),
    .B(\i58/n509 ),
    .Y(\i58/n44 ));
 NOR2xp33_ASAP7_75t_SL \i58/i46  (.A(\i58/n412 ),
    .B(\i58/n538 ),
    .Y(\i58/n437 ));
 AND2x4_ASAP7_75t_SL \i58/i460  (.A(\i58/n495 ),
    .B(\i58/n32 ),
    .Y(\i58/n42 ));
 AND2x4_ASAP7_75t_SL \i58/i461  (.A(\i58/n39 ),
    .B(\i58/n36 ),
    .Y(\i58/n41 ));
 AND2x2_ASAP7_75t_SL \i58/i462  (.A(n5[5]),
    .B(\i58/n22 ),
    .Y(\i58/n39 ));
 AND2x2_ASAP7_75t_SL \i58/i463  (.A(n5[4]),
    .B(\i58/n0 ),
    .Y(\i58/n38 ));
 AND2x2_ASAP7_75t_SL \i58/i464  (.A(n5[3]),
    .B(n5[1]),
    .Y(\i58/n37 ));
 AND2x4_ASAP7_75t_SL \i58/i465  (.A(n5[7]),
    .B(\i58/n23 ),
    .Y(\i58/n36 ));
 AND2x2_ASAP7_75t_SL \i58/i466  (.A(n5[7]),
    .B(n5[6]),
    .Y(\i58/n35 ));
 INVx1_ASAP7_75t_SL \i58/i467  (.A(\i58/n33 ),
    .Y(\i58/n34 ));
 INVx3_ASAP7_75t_SL \i58/i468  (.A(\i58/n517 ),
    .Y(\i58/n29 ));
 NAND2xp5_ASAP7_75t_R \i58/i469  (.A(n5[3]),
    .B(\i58/n24 ),
    .Y(\i58/n28 ));
 NAND3xp33_ASAP7_75t_SL \i58/i47  (.A(\i58/n356 ),
    .B(\i58/n346 ),
    .C(\i58/n282 ),
    .Y(\i58/n436 ));
 NOR2xp33_ASAP7_75t_SL \i58/i470  (.A(\i58/n20 ),
    .B(n5[2]),
    .Y(\i58/n27 ));
 NOR2xp33_ASAP7_75t_SL \i58/i471  (.A(\i58/n24 ),
    .B(n5[0]),
    .Y(\i58/n26 ));
 OR2x2_ASAP7_75t_SL \i58/i472  (.A(\i58/n20 ),
    .B(n5[1]),
    .Y(\i58/n33 ));
 AND2x2_ASAP7_75t_SL \i58/i473  (.A(n5[2]),
    .B(\i58/n20 ),
    .Y(\i58/n32 ));
 AND2x2_ASAP7_75t_SL \i58/i474  (.A(n5[1]),
    .B(\i58/n25 ),
    .Y(\i58/n31 ));
 AND2x2_ASAP7_75t_SL \i58/i475  (.A(n5[5]),
    .B(n5[4]),
    .Y(\i58/n30 ));
 INVx3_ASAP7_75t_SL \i58/i476  (.A(n5[7]),
    .Y(\i58/n4 ));
 INVx2_ASAP7_75t_SL \i58/i477  (.A(n5[3]),
    .Y(\i58/n25 ));
 INVx4_ASAP7_75t_SL \i58/i478  (.A(n5[2]),
    .Y(\i58/n24 ));
 INVx1_ASAP7_75t_SL \i58/i479  (.A(n5[6]),
    .Y(\i58/n23 ));
 NAND3xp33_ASAP7_75t_SL \i58/i48  (.A(\i58/n375 ),
    .B(\i58/n357 ),
    .C(\i58/n343 ),
    .Y(\i58/n435 ));
 INVx2_ASAP7_75t_SL \i58/i480  (.A(n5[4]),
    .Y(\i58/n22 ));
 INVx2_ASAP7_75t_SL \i58/i481  (.A(n5[1]),
    .Y(\i58/n21 ));
 INVx3_ASAP7_75t_SL \i58/i482  (.A(n5[0]),
    .Y(\i58/n20 ));
 AND2x2_ASAP7_75t_SL \i58/i483  (.A(\i58/n555 ),
    .B(\i58/n19 ),
    .Y(\i58/n3 ));
 AND2x2_ASAP7_75t_SL \i58/i484  (.A(\i58/n25 ),
    .B(\i58/n24 ),
    .Y(\i58/n476 ));
 INVx3_ASAP7_75t_SL \i58/i485  (.A(\i58/n478 ),
    .Y(\i58/n479 ));
 AND2x6_ASAP7_75t_SL \i58/i486  (.A(\i58/n477 ),
    .B(\i58/n476 ),
    .Y(\i58/n478 ));
 AND2x2_ASAP7_75t_SL \i58/i487  (.A(n5[1]),
    .B(n5[0]),
    .Y(\i58/n477 ));
 AOI222xp33_ASAP7_75t_R \i58/i488  (.A1(\i58/n61 ),
    .A2(\i58/n83 ),
    .B1(\i58/n79 ),
    .B2(\i58/n478 ),
    .C1(\i58/n68 ),
    .C2(\i58/n61 ),
    .Y(\i58/n480 ));
 AOI211xp5_ASAP7_75t_SL \i58/i489  (.A1(\i58/n172 ),
    .A2(\i58/n478 ),
    .B(\i58/n265 ),
    .C(\i58/n522 ),
    .Y(\i58/n481 ));
 NOR3xp33_ASAP7_75t_SL \i58/i49  (.A(\i58/n323 ),
    .B(\i58/n503 ),
    .C(\i58/n363 ),
    .Y(\i58/n450 ));
 AOI222xp33_ASAP7_75t_SL \i58/i490  (.A1(\i58/n83 ),
    .A2(\i58/n534 ),
    .B1(\i58/n42 ),
    .B2(\i58/n52 ),
    .C1(\i58/n59 ),
    .C2(\i58/n478 ),
    .Y(\i58/n482 ));
 AOI22xp5_ASAP7_75t_SL \i58/i491  (.A1(\i58/n478 ),
    .A2(\i58/n116 ),
    .B1(\i58/n44 ),
    .B2(\i58/n520 ),
    .Y(\i58/n483 ));
 AOI22xp5_ASAP7_75t_SL \i58/i492  (.A1(\i58/n478 ),
    .A2(\i58/n41 ),
    .B1(\i58/n533 ),
    .B2(\i58/n48 ),
    .Y(\i58/n484 ));
 NAND2xp5_ASAP7_75t_SL \i58/i493  (.A(\i58/n478 ),
    .B(\i58/n68 ),
    .Y(\i58/n485 ));
 NAND2xp5_ASAP7_75t_SL \i58/i494  (.A(\i58/n478 ),
    .B(\i58/n83 ),
    .Y(\i58/n486 ));
 NAND2xp5_ASAP7_75t_SL \i58/i495  (.A(\i58/n478 ),
    .B(\i58/n77 ),
    .Y(\i58/n487 ));
 NAND2xp5_ASAP7_75t_SL \i58/i496  (.A(\i58/n478 ),
    .B(\i58/n41 ),
    .Y(\i58/n488 ));
 NOR2xp33_ASAP7_75t_SL \i58/i497  (.A(\i58/n478 ),
    .B(\i58/n46 ),
    .Y(\i58/n489 ));
 NAND2xp5_ASAP7_75t_SL \i58/i498  (.A(\i58/n70 ),
    .B(\i58/n478 ),
    .Y(\i58/n490 ));
 NAND2xp5_ASAP7_75t_SL \i58/i499  (.A(\i58/n478 ),
    .B(\i58/n52 ),
    .Y(\i58/n491 ));
 AND3x4_ASAP7_75t_SL \i58/i5  (.A(\i58/n458 ),
    .B(\i58/n467 ),
    .C(\i58/n464 ),
    .Y(n4[4]));
 NAND2xp5_ASAP7_75t_SL \i58/i50  (.A(\i58/n341 ),
    .B(\i58/n413 ),
    .Y(\i58/n448 ));
 NAND2xp5_ASAP7_75t_SL \i58/i500  (.A(\i58/n478 ),
    .B(\i58/n75 ),
    .Y(\i58/n492 ));
 NAND2xp5_ASAP7_75t_SL \i58/i501  (.A(\i58/n478 ),
    .B(\i58/n59 ),
    .Y(\i58/n493 ));
 AND2x2_ASAP7_75t_SL \i58/i502  (.A(n5[2]),
    .B(n5[0]),
    .Y(\i58/n494 ));
 AND2x2_ASAP7_75t_SL \i58/i503  (.A(\i58/n25 ),
    .B(\i58/n21 ),
    .Y(\i58/n495 ));
 NOR2xp33_ASAP7_75t_L \i58/i504  (.A(\i58/n478 ),
    .B(\i58/n496 ),
    .Y(\i58/n497 ));
 AND2x4_ASAP7_75t_SL \i58/i505  (.A(\i58/n494 ),
    .B(\i58/n495 ),
    .Y(\i58/n496 ));
 INVx3_ASAP7_75t_SL \i58/i506  (.A(\i58/n496 ),
    .Y(\i58/n498 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i58/i507  (.A1(\i58/n61 ),
    .A2(\i58/n496 ),
    .B(\i58/n533 ),
    .C(\i58/n119 ),
    .Y(\i58/n499 ));
 AOI222xp33_ASAP7_75t_SL \i58/i508  (.A1(\i58/n109 ),
    .A2(\i58/n46 ),
    .B1(\i58/n63 ),
    .B2(\i58/n79 ),
    .C1(\i58/n496 ),
    .C2(\i58/n83 ),
    .Y(\i58/n500 ));
 AOI22xp5_ASAP7_75t_SL \i58/i509  (.A1(\i58/n532 ),
    .A2(\i58/n496 ),
    .B1(\i58/n77 ),
    .B2(\i58/n48 ),
    .Y(\i58/n501 ));
 NAND2xp5_ASAP7_75t_SL \i58/i51  (.A(\i58/n356 ),
    .B(\i58/n388 ),
    .Y(\i58/n447 ));
 OAI21xp5_ASAP7_75t_SL \i58/i510  (.A1(\i58/n71 ),
    .A2(\i58/n496 ),
    .B(\i58/n1 ),
    .Y(\i58/n502 ));
 AO22x1_ASAP7_75t_SL \i58/i511  (.A1(\i58/n59 ),
    .A2(\i58/n496 ),
    .B1(\i58/n77 ),
    .B2(\i58/n48 ),
    .Y(\i58/n503 ));
 AOI22xp5_ASAP7_75t_SL \i58/i512  (.A1(\i58/n59 ),
    .A2(\i58/n511 ),
    .B1(\i58/n41 ),
    .B2(\i58/n496 ),
    .Y(\i58/n504 ));
 NAND2xp5_ASAP7_75t_SL \i58/i513  (.A(\i58/n68 ),
    .B(\i58/n496 ),
    .Y(\i58/n505 ));
 NAND2xp5_ASAP7_75t_SL \i58/i514  (.A(\i58/n75 ),
    .B(\i58/n496 ),
    .Y(\i58/n506 ));
 NAND2xp5_ASAP7_75t_SL \i58/i515  (.A(\i58/n50 ),
    .B(\i58/n496 ),
    .Y(\i58/n507 ));
 AOI22xp33_ASAP7_75t_SL \i58/i516  (.A1(\i58/n41 ),
    .A2(\i58/n511 ),
    .B1(\i58/n531 ),
    .B2(\i58/n533 ),
    .Y(\i58/n508 ));
 AND2x4_ASAP7_75t_L \i58/i517  (.A(\i58/n24 ),
    .B(\i58/n20 ),
    .Y(\i58/n509 ));
 AND2x2_ASAP7_75t_SL \i58/i518  (.A(n5[3]),
    .B(\i58/n21 ),
    .Y(\i58/n510 ));
 AOI222xp33_ASAP7_75t_SL \i58/i519  (.A1(\i58/n511 ),
    .A2(\i58/n81 ),
    .B1(\i58/n61 ),
    .B2(\i58/n70 ),
    .C1(\i58/n46 ),
    .C2(\i58/n52 ),
    .Y(\i58/n512 ));
 INVx1_ASAP7_75t_SL \i58/i52  (.A(\i58/n433 ),
    .Y(\i58/n434 ));
 AND2x4_ASAP7_75t_SL \i58/i520  (.A(\i58/n509 ),
    .B(\i58/n510 ),
    .Y(\i58/n511 ));
 AO22x1_ASAP7_75t_SL \i58/i521  (.A1(\i58/n520 ),
    .A2(\i58/n511 ),
    .B1(\i58/n50 ),
    .B2(\i58/n61 ),
    .Y(\i58/n513 ));
 AOI222xp33_ASAP7_75t_SL \i58/i522  (.A1(\i58/n534 ),
    .A2(\i58/n70 ),
    .B1(\i58/n511 ),
    .B2(\i58/n77 ),
    .C1(\i58/n48 ),
    .C2(\i58/n75 ),
    .Y(\i58/n515 ));
 INVx4_ASAP7_75t_SL \i58/i523  (.A(\i58/n511 ),
    .Y(\i58/n514 ));
 AOI221x1_ASAP7_75t_SL \i58/i524  (.A1(\i58/n1 ),
    .A2(\i58/n478 ),
    .B1(\i58/n511 ),
    .B2(\i58/n8 ),
    .C(\i58/n529 ),
    .Y(\i58/n516 ));
 OR2x2_ASAP7_75t_SL \i58/i525  (.A(n5[7]),
    .B(n5[6]),
    .Y(\i58/n517 ));
 INVx3_ASAP7_75t_SL \i58/i526  (.A(\i58/n519 ),
    .Y(\i58/n520 ));
 OR2x6_ASAP7_75t_SL \i58/i527  (.A(\i58/n517 ),
    .B(\i58/n518 ),
    .Y(\i58/n519 ));
 INVx2_ASAP7_75t_SL \i58/i528  (.A(\i58/n39 ),
    .Y(\i58/n518 ));
 OAI211xp5_ASAP7_75t_SL \i58/i529  (.A1(\i58/n519 ),
    .A2(\i58/n147 ),
    .B(\i58/n15 ),
    .C(\i58/n173 ),
    .Y(\i58/n521 ));
 INVxp67_ASAP7_75t_SL \i58/i53  (.A(\i58/n431 ),
    .Y(\i58/n432 ));
 OAI211xp5_ASAP7_75t_SL \i58/i530  (.A1(\i58/n498 ),
    .A2(\i58/n519 ),
    .B(\i58/n178 ),
    .C(\i58/n190 ),
    .Y(\i58/n522 ));
 OAI222xp33_ASAP7_75t_SL \i58/i531  (.A1(\i58/n67 ),
    .A2(\i58/n72 ),
    .B1(\i58/n5 ),
    .B2(\i58/n519 ),
    .C1(\i58/n40 ),
    .C2(\i58/n84 ),
    .Y(\i58/n523 ));
 OAI22xp5_ASAP7_75t_SL \i58/i532  (.A1(\i58/n519 ),
    .A2(\i58/n159 ),
    .B1(\i58/n80 ),
    .B2(\i58/n62 ),
    .Y(\i58/n524 ));
 OAI22xp5_ASAP7_75t_SL \i58/i533  (.A1(\i58/n45 ),
    .A2(\i58/n519 ),
    .B1(\i58/n80 ),
    .B2(\i58/n479 ),
    .Y(\i58/n525 ));
 OAI22xp5_ASAP7_75t_SL \i58/i534  (.A1(\i58/n519 ),
    .A2(\i58/n62 ),
    .B1(\i58/n67 ),
    .B2(\i58/n5 ),
    .Y(\i58/n526 ));
 OAI22xp5_ASAP7_75t_SL \i58/i535  (.A1(\i58/n49 ),
    .A2(\i58/n5 ),
    .B1(\i58/n479 ),
    .B2(\i58/n519 ),
    .Y(\i58/n527 ));
 OAI22xp5_ASAP7_75t_SL \i58/i536  (.A1(\i58/n53 ),
    .A2(\i58/n519 ),
    .B1(\i58/n84 ),
    .B2(\i58/n67 ),
    .Y(\i58/n528 ));
 NOR2xp67_ASAP7_75t_L \i58/i537  (.A(\i58/n519 ),
    .B(\i58/n6 ),
    .Y(\i58/n529 ));
 NAND2xp33_ASAP7_75t_SL \i58/i538  (.A(\i58/n49 ),
    .B(\i58/n519 ),
    .Y(\i58/n530 ));
 INVx2_ASAP7_75t_SL \i58/i539  (.A(\i58/n53 ),
    .Y(\i58/n531 ));
 NAND3xp33_ASAP7_75t_L \i58/i54  (.A(\i58/n370 ),
    .B(\i58/n330 ),
    .C(\i58/n381 ),
    .Y(\i58/n430 ));
 AND2x4_ASAP7_75t_SL \i58/i540  (.A(\i58/n539 ),
    .B(\i58/n29 ),
    .Y(\i58/n532 ));
 AND4x1_ASAP7_75t_SL \i58/i541  (.A(n5[6]),
    .B(\i58/n0 ),
    .C(\i58/n4 ),
    .D(n5[4]),
    .Y(\i58/n533 ));
 AND2x4_ASAP7_75t_SL \i58/i542  (.A(\i58/n509 ),
    .B(\i58/n31 ),
    .Y(\i58/n534 ));
 NAND2xp5_ASAP7_75t_SL \i58/i543  (.A(\i58/n203 ),
    .B(\i58/n535 ),
    .Y(\i58/n536 ));
 AOI22xp5_ASAP7_75t_SL \i58/i544  (.A1(\i58/n531 ),
    .A2(\i58/n532 ),
    .B1(\i58/n533 ),
    .B2(\i58/n534 ),
    .Y(\i58/n535 ));
 NAND2xp33_ASAP7_75t_SL \i58/i545  (.A(\i58/n240 ),
    .B(\i58/n535 ),
    .Y(\i58/n537 ));
 NAND4xp25_ASAP7_75t_SL \i58/i546  (.A(\i58/n332 ),
    .B(\i58/n535 ),
    .C(\i58/n297 ),
    .D(\i58/n484 ),
    .Y(\i58/n538 ));
 AND2x2_ASAP7_75t_SL \i58/i547  (.A(\i58/n0 ),
    .B(\i58/n22 ),
    .Y(\i58/n539 ));
 AND2x2_ASAP7_75t_SL \i58/i548  (.A(n5[6]),
    .B(\i58/n4 ),
    .Y(\i58/n540 ));
 AOI22xp33_ASAP7_75t_SL \i58/i549  (.A1(\i58/n541 ),
    .A2(\i58/n511 ),
    .B1(\i58/n48 ),
    .B2(\i58/n52 ),
    .Y(\i58/n542 ));
 NAND3xp33_ASAP7_75t_L \i58/i55  (.A(\i58/n378 ),
    .B(\i58/n555 ),
    .C(\i58/n19 ),
    .Y(\i58/n429 ));
 AND2x4_ASAP7_75t_SL \i58/i550  (.A(\i58/n539 ),
    .B(\i58/n540 ),
    .Y(\i58/n541 ));
 AOI22xp5_ASAP7_75t_SL \i58/i551  (.A1(\i58/n1 ),
    .A2(\i58/n44 ),
    .B1(\i58/n541 ),
    .B2(\i58/n496 ),
    .Y(\i58/n543 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i58/i552  (.A1(\i58/n66 ),
    .A2(\i58/n496 ),
    .B(\i58/n541 ),
    .C(\i58/n528 ),
    .Y(\i58/n544 ));
 AOI22xp5_ASAP7_75t_SL \i58/i553  (.A1(\i58/n478 ),
    .A2(\i58/n541 ),
    .B1(\i58/n531 ),
    .B2(\i58/n59 ),
    .Y(\i58/n545 ));
 INVx2_ASAP7_75t_SL \i58/i554  (.A(\i58/n541 ),
    .Y(\i58/n546 ));
 AOI221xp5_ASAP7_75t_SL \i58/i555  (.A1(\i58/n163 ),
    .A2(\i58/n73 ),
    .B1(\i58/n541 ),
    .B2(\i58/n63 ),
    .C(\i58/n90 ),
    .Y(\i58/n547 ));
 AOI22xp33_ASAP7_75t_SL \i58/i556  (.A1(\i58/n83 ),
    .A2(\i58/n66 ),
    .B1(\i58/n73 ),
    .B2(\i58/n541 ),
    .Y(\i58/n548 ));
 NAND2xp5_ASAP7_75t_SL \i58/i557  (.A(\i58/n61 ),
    .B(\i58/n541 ),
    .Y(\i58/n549 ));
 NAND2xp5_ASAP7_75t_SL \i58/i558  (.A(\i58/n66 ),
    .B(\i58/n541 ),
    .Y(\i58/n550 ));
 NOR2xp33_ASAP7_75t_SL \i58/i559  (.A(\i58/n79 ),
    .B(\i58/n541 ),
    .Y(\i58/n551 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i58/i56  (.A1(\i58/n57 ),
    .A2(\i58/n51 ),
    .B(\i58/n337 ),
    .C(\i58/n390 ),
    .Y(\i58/n428 ));
 NAND2xp5_ASAP7_75t_SL \i58/i560  (.A(\i58/n73 ),
    .B(\i58/n541 ),
    .Y(\i58/n552 ));
 NAND2xp5_ASAP7_75t_SL \i58/i561  (.A(\i58/n541 ),
    .B(\i58/n42 ),
    .Y(\i58/n553 ));
 NAND2xp5_ASAP7_75t_SL \i58/i562  (.A(\i58/n534 ),
    .B(\i58/n541 ),
    .Y(\i58/n554 ));
 NAND2xp5_ASAP7_75t_SL \i58/i563  (.A(\i58/n46 ),
    .B(\i58/n541 ),
    .Y(\i58/n555 ));
 AND3x1_ASAP7_75t_SL \i58/i564  (.A(\i58/n15 ),
    .B(\i58/n139 ),
    .C(\i58/n553 ),
    .Y(\i58/n556 ));
 AND4x1_ASAP7_75t_SL \i58/i565  (.A(\i58/n187 ),
    .B(\i58/n185 ),
    .C(\i58/n138 ),
    .D(\i58/n16 ),
    .Y(\i58/n557 ));
 NOR4xp25_ASAP7_75t_SL \i58/i566  (.A(\i58/n369 ),
    .B(\i58/n292 ),
    .C(\i58/n120 ),
    .D(\i58/n220 ),
    .Y(\i58/n558 ));
 NAND2xp33_ASAP7_75t_SL \i58/i57  (.A(\i58/n394 ),
    .B(\i58/n389 ),
    .Y(\i58/n427 ));
 NOR2xp33_ASAP7_75t_SL \i58/i58  (.A(\i58/n373 ),
    .B(\i58/n391 ),
    .Y(\i58/n426 ));
 NAND5xp2_ASAP7_75t_SL \i58/i59  (.A(\i58/n325 ),
    .B(\i58/n288 ),
    .C(\i58/n278 ),
    .D(\i58/n298 ),
    .E(\i58/n306 ),
    .Y(\i58/n425 ));
 AND5x2_ASAP7_75t_SL \i58/i6  (.A(\i58/n454 ),
    .B(\i58/n431 ),
    .C(\i58/n421 ),
    .D(\i58/n455 ),
    .E(\i58/n453 ),
    .Y(n4[1]));
 NOR3xp33_ASAP7_75t_SL \i58/i60  (.A(\i58/n342 ),
    .B(\i58/n256 ),
    .C(\i58/n313 ),
    .Y(\i58/n424 ));
 NAND2xp33_ASAP7_75t_SL \i58/i61  (.A(\i58/n372 ),
    .B(\i58/n394 ),
    .Y(\i58/n423 ));
 NAND4xp25_ASAP7_75t_SL \i58/i62  (.A(\i58/n382 ),
    .B(\i58/n357 ),
    .C(\i58/n284 ),
    .D(\i58/n301 ),
    .Y(\i58/n422 ));
 NOR3xp33_ASAP7_75t_SL \i58/i63  (.A(\i58/n393 ),
    .B(\i58/n354 ),
    .C(\i58/n377 ),
    .Y(\i58/n421 ));
 NAND5xp2_ASAP7_75t_SL \i58/i64  (.A(\i58/n362 ),
    .B(\i58/n326 ),
    .C(\i58/n322 ),
    .D(\i58/n207 ),
    .E(\i58/n291 ),
    .Y(\i58/n420 ));
 NAND5xp2_ASAP7_75t_SL \i58/i65  (.A(\i58/n350 ),
    .B(\i58/n319 ),
    .C(\i58/n295 ),
    .D(\i58/n293 ),
    .E(\i58/n331 ),
    .Y(\i58/n419 ));
 NOR4xp25_ASAP7_75t_SL \i58/i66  (.A(\i58/n347 ),
    .B(\i58/n348 ),
    .C(\i58/n209 ),
    .D(\i58/n179 ),
    .Y(\i58/n418 ));
 NAND2xp33_ASAP7_75t_SL \i58/i67  (.A(\i58/n398 ),
    .B(\i58/n376 ),
    .Y(\i58/n417 ));
 NAND4xp25_ASAP7_75t_SL \i58/i68  (.A(\i58/n381 ),
    .B(\i58/n353 ),
    .C(\i58/n384 ),
    .D(\i58/n305 ),
    .Y(\i58/n433 ));
 NOR3x1_ASAP7_75t_SL \i58/i69  (.A(\i58/n358 ),
    .B(\i58/n536 ),
    .C(\i58/n367 ),
    .Y(\i58/n431 ));
 NOR2xp33_ASAP7_75t_SL \i58/i7  (.A(\i58/n444 ),
    .B(\i58/n474 ),
    .Y(\i58/n475 ));
 INVxp67_ASAP7_75t_SL \i58/i70  (.A(\i58/n415 ),
    .Y(\i58/n416 ));
 INVx1_ASAP7_75t_SL \i58/i71  (.A(\i58/n411 ),
    .Y(\i58/n412 ));
 INVxp67_ASAP7_75t_SL \i58/i72  (.A(\i58/n409 ),
    .Y(\i58/n410 ));
 INVxp67_ASAP7_75t_SL \i58/i73  (.A(\i58/n407 ),
    .Y(\i58/n408 ));
 NOR3xp33_ASAP7_75t_SL \i58/i74  (.A(\i58/n371 ),
    .B(\i58/n18 ),
    .C(\i58/n223 ),
    .Y(\i58/n406 ));
 NAND3xp33_ASAP7_75t_SL \i58/i75  (.A(\i58/n254 ),
    .B(\i58/n310 ),
    .C(\i58/n272 ),
    .Y(\i58/n405 ));
 NAND2xp5_ASAP7_75t_SL \i58/i76  (.A(\i58/n359 ),
    .B(\i58/n374 ),
    .Y(\i58/n404 ));
 NOR2xp33_ASAP7_75t_SL \i58/i77  (.A(\i58/n383 ),
    .B(\i58/n349 ),
    .Y(\i58/n403 ));
 NOR2xp33_ASAP7_75t_SL \i58/i78  (.A(\i58/n340 ),
    .B(\i58/n283 ),
    .Y(\i58/n402 ));
 NOR5xp2_ASAP7_75t_SL \i58/i79  (.A(\i58/n274 ),
    .B(\i58/n503 ),
    .C(\i58/n209 ),
    .D(\i58/n250 ),
    .E(\i58/n248 ),
    .Y(\i58/n401 ));
 AND4x2_ASAP7_75t_SL \i58/i8  (.A(\i58/n464 ),
    .B(\i58/n472 ),
    .C(\i58/n471 ),
    .D(\i58/n418 ),
    .Y(n4[5]));
 NOR2xp33_ASAP7_75t_SL \i58/i80  (.A(\i58/n324 ),
    .B(\i58/n351 ),
    .Y(\i58/n400 ));
 AOI211xp5_ASAP7_75t_SL \i58/i81  (.A1(\i58/n312 ),
    .A2(\i58/n104 ),
    .B(\i58/n267 ),
    .C(\i58/n224 ),
    .Y(\i58/n399 ));
 NAND2xp5_ASAP7_75t_SL \i58/i82  (.A(\i58/n277 ),
    .B(\i58/n375 ),
    .Y(\i58/n415 ));
 NAND3xp33_ASAP7_75t_SL \i58/i83  (.A(\i58/n355 ),
    .B(\i58/n332 ),
    .C(\i58/n304 ),
    .Y(\i58/n414 ));
 NOR2x1_ASAP7_75t_SL \i58/i84  (.A(\i58/n364 ),
    .B(\i58/n287 ),
    .Y(\i58/n413 ));
 AND3x1_ASAP7_75t_SL \i58/i85  (.A(\i58/n240 ),
    .B(\i58/n516 ),
    .C(\i58/n483 ),
    .Y(\i58/n411 ));
 NAND3xp33_ASAP7_75t_SL \i58/i86  (.A(\i58/n284 ),
    .B(\i58/n282 ),
    .C(\i58/n557 ),
    .Y(\i58/n409 ));
 NOR3x1_ASAP7_75t_SL \i58/i87  (.A(\i58/n286 ),
    .B(\i58/n308 ),
    .C(\i58/n218 ),
    .Y(\i58/n407 ));
 INVxp33_ASAP7_75t_SL \i58/i88  (.A(\i58/n395 ),
    .Y(\i58/n396 ));
 OAI211xp5_ASAP7_75t_SL \i58/i89  (.A1(\i58/n47 ),
    .A2(\i58/n171 ),
    .B(\i58/n499 ),
    .C(\i58/n241 ),
    .Y(\i58/n392 ));
 AND3x4_ASAP7_75t_SL \i58/i9  (.A(\i58/n466 ),
    .B(\i58/n470 ),
    .C(\i58/n434 ),
    .Y(n4[0]));
 NAND4xp25_ASAP7_75t_SL \i58/i90  (.A(\i58/n544 ),
    .B(\i58/n309 ),
    .C(\i58/n276 ),
    .D(\i58/n239 ),
    .Y(\i58/n391 ));
 NOR3xp33_ASAP7_75t_SL \i58/i91  (.A(\i58/n300 ),
    .B(\i58/n257 ),
    .C(\i58/n259 ),
    .Y(\i58/n390 ));
 NOR4xp25_ASAP7_75t_SL \i58/i92  (.A(\i58/n366 ),
    .B(\i58/n323 ),
    .C(\i58/n215 ),
    .D(\i58/n211 ),
    .Y(\i58/n389 ));
 NOR3xp33_ASAP7_75t_SL \i58/i93  (.A(\i58/n524 ),
    .B(\i58/n243 ),
    .C(\i58/n266 ),
    .Y(\i58/n398 ));
 NOR2xp67_ASAP7_75t_SL \i58/i94  (.A(\i58/n377 ),
    .B(\i58/n338 ),
    .Y(\i58/n388 ));
 NOR2xp33_ASAP7_75t_SL \i58/i95  (.A(\i58/n365 ),
    .B(\i58/n345 ),
    .Y(\i58/n387 ));
 NAND5xp2_ASAP7_75t_SL \i58/i96  (.A(\i58/n280 ),
    .B(\i58/n482 ),
    .C(\i58/n508 ),
    .D(\i58/n214 ),
    .E(\i58/n207 ),
    .Y(\i58/n397 ));
 NAND2xp5_ASAP7_75t_SL \i58/i97  (.A(\i58/n353 ),
    .B(\i58/n384 ),
    .Y(\i58/n386 ));
 NOR3xp33_ASAP7_75t_SL \i58/i98  (.A(\i58/n333 ),
    .B(\i58/n99 ),
    .C(\i58/n213 ),
    .Y(\i58/n395 ));
 NOR2xp33_ASAP7_75t_L \i58/i99  (.A(\i58/n335 ),
    .B(\i58/n318 ),
    .Y(\i58/n394 ));
 AOI22xp5_ASAP7_75t_SL i580 (.A1(n1153),
    .A2(n506),
    .B1(n507),
    .B2(n227),
    .Y(n892));
 AOI22xp5_ASAP7_75t_SL i581 (.A1(n767),
    .A2(n1153),
    .B1(n227),
    .B2(n768),
    .Y(n891));
 AOI22xp33_ASAP7_75t_SL i582 (.A1(n479),
    .A2(n1177),
    .B1(n769),
    .B2(n1211),
    .Y(n890));
 AOI22xp5_ASAP7_75t_SL i583 (.A1(n1155),
    .A2(n802),
    .B1(n803),
    .B2(n226),
    .Y(n889));
 AOI22xp5_ASAP7_75t_SL i584 (.A1(n795),
    .A2(n1155),
    .B1(n1168),
    .B2(n226),
    .Y(n888));
 AOI22xp5_ASAP7_75t_SL i585 (.A1(n781),
    .A2(n481),
    .B1(n782),
    .B2(n480),
    .Y(n887));
 AOI22xp5_ASAP7_75t_SL i586 (.A1(n481),
    .A2(n780),
    .B1(n480),
    .B2(n779),
    .Y(n886));
 AOI22xp5_ASAP7_75t_SL i587 (.A1(n125),
    .A2(n1176),
    .B1(n475),
    .B2(n789),
    .Y(n885));
 AOI22xp5_ASAP7_75t_SL i588 (.A1(n125),
    .A2(n799),
    .B1(n798),
    .B2(n475),
    .Y(n884));
 OAI22xp5_ASAP7_75t_SL i589 (.A1(n474),
    .A2(n779),
    .B1(n780),
    .B2(n124),
    .Y(n883));
 INVx1_ASAP7_75t_SL \i59/i0  (.A(n3[5]),
    .Y(\i59/n0 ));
 INVx2_ASAP7_75t_SL \i59/i1  (.A(\i59/n59 ),
    .Y(\i59/n1 ));
 AND4x2_ASAP7_75t_SL \i59/i10  (.A(\i59/n468 ),
    .B(\i59/n469 ),
    .C(\i59/n466 ),
    .D(\i59/n467 ),
    .Y(n2[7]));
 NOR3xp33_ASAP7_75t_SL \i59/i100  (.A(\i59/n89 ),
    .B(\i59/n217 ),
    .C(\i59/n255 ),
    .Y(\i59/n387 ));
 OAI211xp5_ASAP7_75t_SL \i59/i101  (.A1(\i59/n64 ),
    .A2(\i59/n176 ),
    .B(\i59/n528 ),
    .C(\i59/n542 ),
    .Y(\i59/n386 ));
 NOR2xp33_ASAP7_75t_SL \i59/i102  (.A(\i59/n341 ),
    .B(\i59/n13 ),
    .Y(\i59/n385 ));
 OAI21xp5_ASAP7_75t_SL \i59/i103  (.A1(\i59/n54 ),
    .A2(\i59/n76 ),
    .B(\i59/n344 ),
    .Y(\i59/n384 ));
 NOR4xp25_ASAP7_75t_SL \i59/i104  (.A(\i59/n241 ),
    .B(\i59/n242 ),
    .C(\i59/n208 ),
    .D(\i59/n514 ),
    .Y(\i59/n383 ));
 NOR3xp33_ASAP7_75t_SL \i59/i105  (.A(\i59/n502 ),
    .B(\i59/n127 ),
    .C(\i59/n187 ),
    .Y(\i59/n382 ));
 NAND2xp5_ASAP7_75t_SL \i59/i106  (.A(\i59/n229 ),
    .B(\i59/n526 ),
    .Y(\i59/n381 ));
 NOR2xp33_ASAP7_75t_L \i59/i107  (.A(\i59/n284 ),
    .B(\i59/n306 ),
    .Y(\i59/n397 ));
 OAI211xp5_ASAP7_75t_SL \i59/i108  (.A1(\i59/n43 ),
    .A2(\i59/n54 ),
    .B(\i59/n232 ),
    .C(\i59/n221 ),
    .Y(\i59/n380 ));
 NAND3xp33_ASAP7_75t_L \i59/i109  (.A(\i59/n257 ),
    .B(\i59/n260 ),
    .C(\i59/n308 ),
    .Y(\i59/n379 ));
 NAND4xp25_ASAP7_75t_SL \i59/i11  (.A(\i59/n460 ),
    .B(\i59/n399 ),
    .C(\i59/n389 ),
    .D(\i59/n404 ),
    .Y(\i59/n483 ));
 NAND2xp5_ASAP7_75t_SL \i59/i110  (.A(\i59/n527 ),
    .B(\i59/n232 ),
    .Y(\i59/n378 ));
 NAND2xp5_ASAP7_75t_L \i59/i111  (.A(\i59/n550 ),
    .B(\i59/n270 ),
    .Y(\i59/n377 ));
 NOR3xp33_ASAP7_75t_SL \i59/i112  (.A(\i59/n303 ),
    .B(\i59/n209 ),
    .C(\i59/n226 ),
    .Y(\i59/n376 ));
 NOR3xp33_ASAP7_75t_SL \i59/i113  (.A(\i59/n12 ),
    .B(\i59/n197 ),
    .C(\i59/n181 ),
    .Y(\i59/n375 ));
 NOR4xp25_ASAP7_75t_SL \i59/i114  (.A(\i59/n12 ),
    .B(\i59/n210 ),
    .C(\i59/n199 ),
    .D(\i59/n92 ),
    .Y(\i59/n374 ));
 AOI211x1_ASAP7_75t_SL \i59/i115  (.A1(\i59/n109 ),
    .A2(\i59/n73 ),
    .B(\i59/n238 ),
    .C(\i59/n230 ),
    .Y(\i59/n395 ));
 NOR3xp33_ASAP7_75t_SL \i59/i116  (.A(\i59/n264 ),
    .B(\i59/n127 ),
    .C(\i59/n245 ),
    .Y(\i59/n394 ));
 NOR2xp33_ASAP7_75t_L \i59/i117  (.A(\i59/n226 ),
    .B(\i59/n350 ),
    .Y(\i59/n373 ));
 NOR2x1_ASAP7_75t_SL \i59/i118  (.A(\i59/n338 ),
    .B(\i59/n271 ),
    .Y(\i59/n393 ));
 NOR2xp33_ASAP7_75t_SL \i59/i119  (.A(\i59/n276 ),
    .B(\i59/n345 ),
    .Y(\i59/n391 ));
 NOR3xp33_ASAP7_75t_SL \i59/i12  (.A(\i59/n519 ),
    .B(\i59/n472 ),
    .C(\i59/n456 ),
    .Y(\i59/n482 ));
 NAND2xp5_ASAP7_75t_SL \i59/i120  (.A(\i59/n221 ),
    .B(\i59/n283 ),
    .Y(\i59/n390 ));
 NOR2xp67_ASAP7_75t_SL \i59/i121  (.A(\i59/n323 ),
    .B(\i59/n347 ),
    .Y(\i59/n389 ));
 NOR3x1_ASAP7_75t_SL \i59/i122  (.A(\i59/n503 ),
    .B(\i59/n255 ),
    .C(\i59/n500 ),
    .Y(\i59/n388 ));
 INVx1_ASAP7_75t_SL \i59/i123  (.A(\i59/n369 ),
    .Y(\i59/n370 ));
 NOR2xp33_ASAP7_75t_SL \i59/i124  (.A(\i59/n485 ),
    .B(\i59/n318 ),
    .Y(\i59/n368 ));
 NAND5xp2_ASAP7_75t_SL \i59/i125  (.A(\i59/n90 ),
    .B(\i59/n200 ),
    .C(\i59/n163 ),
    .D(\i59/n166 ),
    .E(\i59/n194 ),
    .Y(\i59/n367 ));
 NOR2xp33_ASAP7_75t_SL \i59/i126  (.A(\i59/n319 ),
    .B(\i59/n333 ),
    .Y(\i59/n366 ));
 OAI211xp5_ASAP7_75t_SL \i59/i127  (.A1(\i59/n43 ),
    .A2(\i59/n179 ),
    .B(\i59/n326 ),
    .C(\i59/n263 ),
    .Y(\i59/n365 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i59/i128  (.A1(\i59/n74 ),
    .A2(\i59/n195 ),
    .B(\i59/n4 ),
    .C(\i59/n254 ),
    .Y(\i59/n364 ));
 NAND3xp33_ASAP7_75t_SL \i59/i129  (.A(\i59/n513 ),
    .B(\i59/n247 ),
    .C(\i59/n239 ),
    .Y(\i59/n363 ));
 AND2x2_ASAP7_75t_SL \i59/i13  (.A(\i59/n477 ),
    .B(\i59/n478 ),
    .Y(n2[2]));
 NOR3xp33_ASAP7_75t_SL \i59/i130  (.A(\i59/n273 ),
    .B(\i59/n225 ),
    .C(\i59/n231 ),
    .Y(\i59/n362 ));
 NAND3xp33_ASAP7_75t_L \i59/i131  (.A(\i59/n224 ),
    .B(\i59/n221 ),
    .C(\i59/n310 ),
    .Y(\i59/n361 ));
 NOR3xp33_ASAP7_75t_SL \i59/i132  (.A(\i59/n287 ),
    .B(\i59/n261 ),
    .C(\i59/n225 ),
    .Y(\i59/n360 ));
 AOI211xp5_ASAP7_75t_SL \i59/i133  (.A1(\i59/n69 ),
    .A2(\i59/n79 ),
    .B(\i59/n331 ),
    .C(\i59/n128 ),
    .Y(\i59/n359 ));
 OAI221xp5_ASAP7_75t_SL \i59/i134  (.A1(\i59/n176 ),
    .A2(\i59/n43 ),
    .B1(\i59/n115 ),
    .B2(\i59/n58 ),
    .C(\i59/n185 ),
    .Y(\i59/n358 ));
 AOI211xp5_ASAP7_75t_SL \i59/i135  (.A1(\i59/n80 ),
    .A2(\i59/n42 ),
    .B(\i59/n256 ),
    .C(\i59/n265 ),
    .Y(\i59/n357 ));
 NAND2xp33_ASAP7_75t_SL \i59/i136  (.A(\i59/n285 ),
    .B(\i59/n281 ),
    .Y(\i59/n356 ));
 NOR2xp33_ASAP7_75t_SL \i59/i137  (.A(\i59/n330 ),
    .B(\i59/n294 ),
    .Y(\i59/n355 ));
 NAND4xp25_ASAP7_75t_SL \i59/i138  (.A(\i59/n547 ),
    .B(\i59/n10 ),
    .C(\i59/n203 ),
    .D(\i59/n146 ),
    .Y(\i59/n354 ));
 OAI221xp5_ASAP7_75t_SL \i59/i139  (.A1(\i59/n248 ),
    .A2(\i59/n86 ),
    .B1(\i59/n544 ),
    .B2(\i59/n487 ),
    .C(\i59/n206 ),
    .Y(\i59/n353 ));
 NOR3xp33_ASAP7_75t_SL \i59/i14  (.A(\i59/n457 ),
    .B(\i59/n406 ),
    .C(\i59/n461 ),
    .Y(\i59/n481 ));
 NAND4xp25_ASAP7_75t_SL \i59/i140  (.A(\i59/n211 ),
    .B(\i59/n216 ),
    .C(\i59/n189 ),
    .D(\i59/n532 ),
    .Y(\i59/n352 ));
 NOR2xp33_ASAP7_75t_SL \i59/i141  (.A(\i59/n296 ),
    .B(\i59/n304 ),
    .Y(\i59/n372 ));
 NAND2xp33_ASAP7_75t_L \i59/i142  (.A(\i59/n337 ),
    .B(\i59/n234 ),
    .Y(\i59/n351 ));
 NOR2xp33_ASAP7_75t_SL \i59/i143  (.A(\i59/n313 ),
    .B(\i59/n334 ),
    .Y(\i59/n371 ));
 NAND2xp5_ASAP7_75t_SL \i59/i144  (.A(\i59/n223 ),
    .B(\i59/n275 ),
    .Y(\i59/n369 ));
 NOR2xp67_ASAP7_75t_SL \i59/i145  (.A(\i59/n274 ),
    .B(\i59/n282 ),
    .Y(\i59/n14 ));
 INVxp67_ASAP7_75t_SL \i59/i146  (.A(\i59/n347 ),
    .Y(\i59/n348 ));
 INVxp33_ASAP7_75t_SL \i59/i147  (.A(\i59/n345 ),
    .Y(\i59/n346 ));
 INVx1_ASAP7_75t_SL \i59/i148  (.A(\i59/n342 ),
    .Y(\i59/n343 ));
 INVxp67_ASAP7_75t_SL \i59/i149  (.A(\i59/n338 ),
    .Y(\i59/n339 ));
 NOR3xp33_ASAP7_75t_SL \i59/i15  (.A(\i59/n437 ),
    .B(\i59/n442 ),
    .C(\i59/n421 ),
    .Y(\i59/n480 ));
 INVxp67_ASAP7_75t_SL \i59/i150  (.A(\i59/n13 ),
    .Y(\i59/n337 ));
 INVxp67_ASAP7_75t_SL \i59/i151  (.A(\i59/n335 ),
    .Y(\i59/n336 ));
 NAND2xp5_ASAP7_75t_SL \i59/i152  (.A(\i59/n260 ),
    .B(\i59/n258 ),
    .Y(\i59/n334 ));
 NAND2xp33_ASAP7_75t_SL \i59/i153  (.A(\i59/n508 ),
    .B(\i59/n250 ),
    .Y(\i59/n333 ));
 AOI21xp5_ASAP7_75t_SL \i59/i154  (.A1(\i59/n183 ),
    .A2(\i59/n87 ),
    .B(\i59/n261 ),
    .Y(\i59/n332 ));
 OAI22xp5_ASAP7_75t_SL \i59/i155  (.A1(\i59/n107 ),
    .A2(\i59/n142 ),
    .B1(\i59/n82 ),
    .B2(\i59/n125 ),
    .Y(\i59/n331 ));
 NAND4xp25_ASAP7_75t_SL \i59/i156  (.A(\i59/n191 ),
    .B(\i59/n137 ),
    .C(\i59/n136 ),
    .D(\i59/n112 ),
    .Y(\i59/n330 ));
 NAND3xp33_ASAP7_75t_SL \i59/i157  (.A(\i59/n133 ),
    .B(\i59/n145 ),
    .C(\i59/n5 ),
    .Y(\i59/n329 ));
 NAND3xp33_ASAP7_75t_SL \i59/i158  (.A(\i59/n175 ),
    .B(\i59/n190 ),
    .C(\i59/n486 ),
    .Y(\i59/n328 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i59/i159  (.A1(\i59/n45 ),
    .A2(\i59/n40 ),
    .B(\i59/n80 ),
    .C(\i59/n230 ),
    .Y(\i59/n327 ));
 NOR3xp33_ASAP7_75t_SL \i59/i16  (.A(\i59/n447 ),
    .B(\i59/n449 ),
    .C(\i59/n432 ),
    .Y(\i59/n479 ));
 AOI222xp33_ASAP7_75t_SL \i59/i160  (.A1(\i59/n62 ),
    .A2(\i59/n85 ),
    .B1(\i59/n81 ),
    .B2(\i59/n47 ),
    .C1(\i59/n73 ),
    .C2(\i59/n62 ),
    .Y(\i59/n326 ));
 NOR2xp33_ASAP7_75t_SL \i59/i161  (.A(\i59/n500 ),
    .B(\i59/n240 ),
    .Y(\i59/n325 ));
 OAI21xp5_ASAP7_75t_SL \i59/i162  (.A1(\i59/n82 ),
    .A2(\i59/n549 ),
    .B(\i59/n97 ),
    .Y(\i59/n324 ));
 NAND4xp25_ASAP7_75t_SL \i59/i163  (.A(\i59/n204 ),
    .B(\i59/n147 ),
    .C(\i59/n134 ),
    .D(\i59/n173 ),
    .Y(\i59/n323 ));
 AOI211xp5_ASAP7_75t_SL \i59/i164  (.A1(\i59/n40 ),
    .A2(\i59/n1 ),
    .B(\i59/n144 ),
    .C(\i59/n139 ),
    .Y(\i59/n322 ));
 NOR2xp33_ASAP7_75t_L \i59/i165  (.A(\i59/n214 ),
    .B(\i59/n252 ),
    .Y(\i59/n321 ));
 NOR2xp33_ASAP7_75t_L \i59/i166  (.A(\i59/n213 ),
    .B(\i59/n233 ),
    .Y(\i59/n320 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i59/i167  (.A1(\i59/n64 ),
    .A2(\i59/n39 ),
    .B(\i59/n509 ),
    .C(\i59/n545 ),
    .Y(\i59/n319 ));
 NAND3xp33_ASAP7_75t_SL \i59/i168  (.A(\i59/n550 ),
    .B(\i59/n189 ),
    .C(\i59/n88 ),
    .Y(\i59/n318 ));
 NOR3xp33_ASAP7_75t_SL \i59/i169  (.A(\i59/n237 ),
    .B(\i59/n150 ),
    .C(\i59/n201 ),
    .Y(\i59/n317 ));
 NOR4xp25_ASAP7_75t_SL \i59/i17  (.A(\i59/n430 ),
    .B(\i59/n418 ),
    .C(\i59/n422 ),
    .D(\i59/n493 ),
    .Y(\i59/n478 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i59/i170  (.A1(\i59/n62 ),
    .A2(\i59/n67 ),
    .B(\i59/n53 ),
    .C(\i59/n126 ),
    .Y(\i59/n316 ));
 NAND4xp25_ASAP7_75t_SL \i59/i171  (.A(\i59/n186 ),
    .B(\i59/n121 ),
    .C(\i59/n9 ),
    .D(\i59/n11 ),
    .Y(\i59/n315 ));
 AOI222xp33_ASAP7_75t_SL \i59/i172  (.A1(\i59/n85 ),
    .A2(\i59/n69 ),
    .B1(\i59/n40 ),
    .B2(\i59/n50 ),
    .C1(\i59/n61 ),
    .C2(\i59/n47 ),
    .Y(\i59/n314 ));
 OAI211xp5_ASAP7_75t_SL \i59/i173  (.A1(\i59/n55 ),
    .A2(\i59/n510 ),
    .B(\i59/n100 ),
    .C(\i59/n119 ),
    .Y(\i59/n313 ));
 OAI31xp33_ASAP7_75t_SL \i59/i174  (.A1(\i59/n38 ),
    .A2(\i59/n48 ),
    .A3(\i59/n80 ),
    .B(\i59/n71 ),
    .Y(\i59/n312 ));
 AOI221xp5_ASAP7_75t_SL \i59/i175  (.A1(\i59/n167 ),
    .A2(\i59/n56 ),
    .B1(\i59/n50 ),
    .B2(\i59/n87 ),
    .C(\i59/n149 ),
    .Y(\i59/n311 ));
 NOR2xp33_ASAP7_75t_SL \i59/i176  (.A(\i59/n132 ),
    .B(\i59/n501 ),
    .Y(\i59/n310 ));
 OAI221xp5_ASAP7_75t_SL \i59/i177  (.A1(\i59/n39 ),
    .A2(\i59/n37 ),
    .B1(\i59/n49 ),
    .B2(\i59/n66 ),
    .C(\i59/n155 ),
    .Y(\i59/n350 ));
 NAND2xp5_ASAP7_75t_SL \i59/i178  (.A(\i59/n512 ),
    .B(\i59/n212 ),
    .Y(\i59/n347 ));
 OAI221xp5_ASAP7_75t_SL \i59/i179  (.A1(\i59/n510 ),
    .A2(\i59/n52 ),
    .B1(\i59/n506 ),
    .B2(\i59/n54 ),
    .C(\i59/n5 ),
    .Y(\i59/n345 ));
 NOR5xp2_ASAP7_75t_SL \i59/i18  (.A(\i59/n518 ),
    .B(\i59/n427 ),
    .C(\i59/n457 ),
    .D(\i59/n410 ),
    .E(\i59/n392 ),
    .Y(\i59/n477 ));
 OAI21xp5_ASAP7_75t_SL \i59/i180  (.A1(\i59/n56 ),
    .A2(\i59/n124 ),
    .B(\i59/n177 ),
    .Y(\i59/n344 ));
 NOR2xp33_ASAP7_75t_SL \i59/i181  (.A(\i59/n127 ),
    .B(\i59/n264 ),
    .Y(\i59/n309 ));
 NAND2xp5_ASAP7_75t_SL \i59/i182  (.A(\i59/n215 ),
    .B(\i59/n250 ),
    .Y(\i59/n342 ));
 NOR2xp33_ASAP7_75t_SL \i59/i183  (.A(\i59/n515 ),
    .B(\i59/n514 ),
    .Y(\i59/n308 ));
 NAND2xp5_ASAP7_75t_SL \i59/i184  (.A(\i59/n218 ),
    .B(\i59/n220 ),
    .Y(\i59/n341 ));
 NAND2xp5_ASAP7_75t_SL \i59/i185  (.A(\i59/n529 ),
    .B(\i59/n545 ),
    .Y(\i59/n340 ));
 OAI221xp5_ASAP7_75t_SL \i59/i186  (.A1(\i59/n486 ),
    .A2(\i59/n84 ),
    .B1(\i59/n68 ),
    .B2(\i59/n82 ),
    .C(\i59/n141 ),
    .Y(\i59/n338 ));
 NAND2x1_ASAP7_75t_SL \i59/i187  (.A(\i59/n246 ),
    .B(\i59/n224 ),
    .Y(\i59/n13 ));
 NAND3xp33_ASAP7_75t_SL \i59/i188  (.A(\i59/n140 ),
    .B(\i59/n135 ),
    .C(\i59/n131 ),
    .Y(\i59/n12 ));
 NOR2xp33_ASAP7_75t_SL \i59/i189  (.A(\i59/n265 ),
    .B(\i59/n256 ),
    .Y(\i59/n307 ));
 NOR3xp33_ASAP7_75t_SL \i59/i19  (.A(\i59/n520 ),
    .B(\i59/n458 ),
    .C(\i59/n470 ),
    .Y(\i59/n476 ));
 OAI211xp5_ASAP7_75t_SL \i59/i190  (.A1(\i59/n78 ),
    .A2(\i59/n70 ),
    .B(\i59/n205 ),
    .C(\i59/n531 ),
    .Y(\i59/n335 ));
 INVxp67_ASAP7_75t_SL \i59/i191  (.A(\i59/n304 ),
    .Y(\i59/n305 ));
 INVxp67_ASAP7_75t_SL \i59/i192  (.A(\i59/n302 ),
    .Y(\i59/n303 ));
 INVxp67_ASAP7_75t_SL \i59/i193  (.A(\i59/n300 ),
    .Y(\i59/n301 ));
 INVx2_ASAP7_75t_SL \i59/i194  (.A(\i59/n542 ),
    .Y(\i59/n299 ));
 INVx1_ASAP7_75t_SL \i59/i195  (.A(\i59/n297 ),
    .Y(\i59/n298 ));
 OAI22xp5_ASAP7_75t_SL \i59/i196  (.A1(\i59/n506 ),
    .A2(\i59/n533 ),
    .B1(\i59/n74 ),
    .B2(\i59/n70 ),
    .Y(\i59/n296 ));
 AOI21xp5_ASAP7_75t_SL \i59/i197  (.A1(\i59/n105 ),
    .A2(\i59/n75 ),
    .B(\i59/n128 ),
    .Y(\i59/n295 ));
 OAI22xp5_ASAP7_75t_SL \i59/i198  (.A1(\i59/n54 ),
    .A2(\i59/n102 ),
    .B1(\i59/n52 ),
    .B2(\i59/n193 ),
    .Y(\i59/n294 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i59/i199  (.A1(\i59/n69 ),
    .A2(\i59/n65 ),
    .B(\i59/n73 ),
    .C(\i59/n94 ),
    .Y(\i59/n293 ));
 INVx3_ASAP7_75t_SL \i59/i2  (.A(\i59/n80 ),
    .Y(\i59/n2 ));
 NOR3xp33_ASAP7_75t_SL \i59/i20  (.A(\i59/n439 ),
    .B(\i59/n462 ),
    .C(\i59/n427 ),
    .Y(\i59/n475 ));
 AOI21xp5_ASAP7_75t_SL \i59/i200  (.A1(\i59/n178 ),
    .A2(\i59/n69 ),
    .B(\i59/n243 ),
    .Y(\i59/n292 ));
 AOI22xp5_ASAP7_75t_SL \i59/i201  (.A1(\i59/n48 ),
    .A2(\i59/n106 ),
    .B1(\i59/n77 ),
    .B2(\i59/n171 ),
    .Y(\i59/n291 ));
 AOI211xp5_ASAP7_75t_SL \i59/i202  (.A1(\i59/n48 ),
    .A2(\i59/n51 ),
    .B(\i59/n128 ),
    .C(\i59/n96 ),
    .Y(\i59/n290 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i59/i203  (.A1(\i59/n71 ),
    .A2(\i59/n67 ),
    .B(\i59/n63 ),
    .C(\i59/n499 ),
    .Y(\i59/n289 ));
 OAI22xp5_ASAP7_75t_SL \i59/i204  (.A1(\i59/n64 ),
    .A2(\i59/n165 ),
    .B1(\i59/n4 ),
    .B2(\i59/n164 ),
    .Y(\i59/n288 ));
 OAI22xp5_ASAP7_75t_SL \i59/i205  (.A1(\i59/n59 ),
    .A2(\i59/n157 ),
    .B1(\i59/n52 ),
    .B2(\i59/n74 ),
    .Y(\i59/n287 ));
 AOI221xp5_ASAP7_75t_SL \i59/i206  (.A1(\i59/n44 ),
    .A2(\i59/n80 ),
    .B1(\i59/n40 ),
    .B2(\i59/n38 ),
    .C(\i59/n244 ),
    .Y(\i59/n286 ));
 AND4x1_ASAP7_75t_SL \i59/i207  (.A(\i59/n134 ),
    .B(\i59/n7 ),
    .C(\i59/n8 ),
    .D(\i59/n141 ),
    .Y(\i59/n285 ));
 NAND4xp25_ASAP7_75t_SL \i59/i208  (.A(\i59/n129 ),
    .B(\i59/n152 ),
    .C(\i59/n546 ),
    .D(\i59/n534 ),
    .Y(\i59/n284 ));
 AOI222xp33_ASAP7_75t_SL \i59/i209  (.A1(\i59/n117 ),
    .A2(\i59/n44 ),
    .B1(\i59/n65 ),
    .B2(\i59/n81 ),
    .C1(\i59/n67 ),
    .C2(\i59/n85 ),
    .Y(\i59/n283 ));
 AND4x1_ASAP7_75t_SL \i59/i21  (.A(\i59/n454 ),
    .B(\i59/n459 ),
    .C(\i59/n443 ),
    .D(\i59/n429 ),
    .Y(\i59/n474 ));
 NAND4xp25_ASAP7_75t_SL \i59/i210  (.A(\i59/n140 ),
    .B(\i59/n137 ),
    .C(\i59/n539 ),
    .D(\i59/n135 ),
    .Y(\i59/n282 ));
 AOI22xp5_ASAP7_75t_SL \i59/i211  (.A1(\i59/n504 ),
    .A2(\i59/n101 ),
    .B1(\i59/n79 ),
    .B2(\i59/n118 ),
    .Y(\i59/n281 ));
 AOI22xp5_ASAP7_75t_SL \i59/i212  (.A1(\i59/n47 ),
    .A2(\i59/n123 ),
    .B1(\i59/n42 ),
    .B2(\i59/n504 ),
    .Y(\i59/n280 ));
 OAI211xp5_ASAP7_75t_SL \i59/i213  (.A1(\i59/n72 ),
    .A2(\i59/n190 ),
    .B(\i59/n91 ),
    .C(\i59/n143 ),
    .Y(\i59/n279 ));
 NAND4xp25_ASAP7_75t_SL \i59/i214  (.A(\i59/n8 ),
    .B(\i59/n158 ),
    .C(\i59/n172 ),
    .D(\i59/n170 ),
    .Y(\i59/n278 ));
 OAI22xp5_ASAP7_75t_SL \i59/i215  (.A1(\i59/n487 ),
    .A2(\i59/n161 ),
    .B1(\i59/n4 ),
    .B2(\i59/n120 ),
    .Y(\i59/n277 ));
 OAI22xp33_ASAP7_75t_SL \i59/i216  (.A1(\i59/n2 ),
    .A2(\i59/n113 ),
    .B1(\i59/n76 ),
    .B2(\i59/n37 ),
    .Y(\i59/n276 ));
 AOI211x1_ASAP7_75t_SL \i59/i217  (.A1(\i59/n174 ),
    .A2(\i59/n87 ),
    .B(\i59/n548 ),
    .C(\i59/n192 ),
    .Y(\i59/n275 ));
 NAND4xp25_ASAP7_75t_SL \i59/i218  (.A(\i59/n180 ),
    .B(\i59/n196 ),
    .C(\i59/n114 ),
    .D(\i59/n131 ),
    .Y(\i59/n274 ));
 OAI22xp5_ASAP7_75t_SL \i59/i219  (.A1(\i59/n66 ),
    .A2(\i59/n99 ),
    .B1(\i59/n82 ),
    .B2(\i59/n4 ),
    .Y(\i59/n273 ));
 NAND3xp33_ASAP7_75t_SL \i59/i22  (.A(\i59/n414 ),
    .B(\i59/n389 ),
    .C(\i59/n411 ),
    .Y(\i59/n472 ));
 OAI221xp5_ASAP7_75t_R \i59/i220  (.A1(\i59/n116 ),
    .A2(\i59/n525 ),
    .B1(\i59/n74 ),
    .B2(\i59/n86 ),
    .C(\i59/n162 ),
    .Y(\i59/n272 ));
 OAI221xp5_ASAP7_75t_SL \i59/i221  (.A1(\i59/n66 ),
    .A2(\i59/n487 ),
    .B1(\i59/n43 ),
    .B2(\i59/n525 ),
    .C(\i59/n151 ),
    .Y(\i59/n271 ));
 AOI222xp33_ASAP7_75t_SL \i59/i222  (.A1(\i59/n57 ),
    .A2(\i59/n83 ),
    .B1(\i59/n62 ),
    .B2(\i59/n75 ),
    .C1(\i59/n44 ),
    .C2(\i59/n50 ),
    .Y(\i59/n270 ));
 OAI221xp5_ASAP7_75t_SL \i59/i223  (.A1(\i59/n544 ),
    .A2(\i59/n37 ),
    .B1(\i59/n2 ),
    .B2(\i59/n55 ),
    .C(\i59/n110 ),
    .Y(\i59/n269 ));
 OAI211xp5_ASAP7_75t_SL \i59/i224  (.A1(\i59/n55 ),
    .A2(\i59/n142 ),
    .B(\i59/n138 ),
    .C(\i59/n95 ),
    .Y(\i59/n268 ));
 AOI221xp5_ASAP7_75t_SL \i59/i225  (.A1(\i59/n202 ),
    .A2(\i59/n61 ),
    .B1(\i59/n85 ),
    .B2(\i59/n69 ),
    .C(\i59/n130 ),
    .Y(\i59/n267 ));
 AOI22xp33_ASAP7_75t_SL \i59/i226  (.A1(\i59/n48 ),
    .A2(\i59/n202 ),
    .B1(\i59/n75 ),
    .B2(\i59/n57 ),
    .Y(\i59/n266 ));
 OAI221xp5_ASAP7_75t_SL \i59/i227  (.A1(\i59/n66 ),
    .A2(\i59/n74 ),
    .B1(\i59/n70 ),
    .B2(\i59/n84 ),
    .C(\i59/n154 ),
    .Y(\i59/n306 ));
 OAI221xp5_ASAP7_75t_SL \i59/i228  (.A1(\i59/n509 ),
    .A2(\i59/n41 ),
    .B1(\i59/n487 ),
    .B2(\i59/n58 ),
    .C(\i59/n104 ),
    .Y(\i59/n304 ));
 AOI221x1_ASAP7_75t_SL \i59/i229  (.A1(\i59/n1 ),
    .A2(\i59/n47 ),
    .B1(\i59/n57 ),
    .B2(\i59/n6 ),
    .C(\i59/n498 ),
    .Y(\i59/n302 ));
 NOR2xp33_ASAP7_75t_SL \i59/i23  (.A(\i59/n446 ),
    .B(\i59/n444 ),
    .Y(\i59/n471 ));
 OAI21xp5_ASAP7_75t_L \i59/i230  (.A1(\i59/n193 ),
    .A2(\i59/n58 ),
    .B(\i59/n111 ),
    .Y(\i59/n300 ));
 OAI221xp5_ASAP7_75t_SL \i59/i231  (.A1(\i59/n160 ),
    .A2(\i59/n510 ),
    .B1(\i59/n82 ),
    .B2(\i59/n43 ),
    .C(\i59/n184 ),
    .Y(\i59/n297 ));
 INVxp67_ASAP7_75t_SL \i59/i232  (.A(\i59/n262 ),
    .Y(\i59/n263 ));
 INVxp67_ASAP7_75t_SL \i59/i233  (.A(\i59/n258 ),
    .Y(\i59/n259 ));
 INVxp67_ASAP7_75t_SL \i59/i234  (.A(\i59/n256 ),
    .Y(\i59/n257 ));
 INVx1_ASAP7_75t_SL \i59/i235  (.A(\i59/n253 ),
    .Y(\i59/n254 ));
 INVxp67_ASAP7_75t_SL \i59/i236  (.A(\i59/n251 ),
    .Y(\i59/n252 ));
 INVxp67_ASAP7_75t_SL \i59/i237  (.A(\i59/n530 ),
    .Y(\i59/n249 ));
 NOR2xp33_ASAP7_75t_SL \i59/i238  (.A(\i59/n497 ),
    .B(\i59/n178 ),
    .Y(\i59/n248 ));
 OAI21xp5_ASAP7_75t_SL \i59/i239  (.A1(\i59/n45 ),
    .A2(\i59/n42 ),
    .B(\i59/n81 ),
    .Y(\i59/n247 ));
 NAND2xp5_ASAP7_75t_SL \i59/i24  (.A(\i59/n448 ),
    .B(\i59/n438 ),
    .Y(\i59/n470 ));
 AOI22xp5_ASAP7_75t_SL \i59/i240  (.A1(\i59/n48 ),
    .A2(\i59/n57 ),
    .B1(\i59/n85 ),
    .B2(\i59/n56 ),
    .Y(\i59/n246 ));
 OAI21xp5_ASAP7_75t_SL \i59/i241  (.A1(\i59/n510 ),
    .A2(\i59/n41 ),
    .B(\i59/n143 ),
    .Y(\i59/n245 ));
 AOI21xp33_ASAP7_75t_SL \i59/i242  (.A1(\i59/n68 ),
    .A2(\i59/n58 ),
    .B(\i59/n175 ),
    .Y(\i59/n244 ));
 OAI21xp5_ASAP7_75t_SL \i59/i243  (.A1(\i59/n2 ),
    .A2(\i59/n64 ),
    .B(\i59/n185 ),
    .Y(\i59/n265 ));
 NAND2xp5_ASAP7_75t_L \i59/i244  (.A(\i59/n535 ),
    .B(\i59/n153 ),
    .Y(\i59/n243 ));
 OAI21xp33_ASAP7_75t_SL \i59/i245  (.A1(\i59/n60 ),
    .A2(\i59/n64 ),
    .B(\i59/n539 ),
    .Y(\i59/n242 ));
 AOI21xp5_ASAP7_75t_SL \i59/i246  (.A1(\i59/n39 ),
    .A2(\i59/n76 ),
    .B(\i59/n487 ),
    .Y(\i59/n264 ));
 AOI21xp33_ASAP7_75t_SL \i59/i247  (.A1(\i59/n76 ),
    .A2(\i59/n46 ),
    .B(\i59/n175 ),
    .Y(\i59/n241 ));
 OAI21xp33_ASAP7_75t_SL \i59/i248  (.A1(\i59/n59 ),
    .A2(\i59/n64 ),
    .B(\i59/n136 ),
    .Y(\i59/n240 ));
 NOR2xp33_ASAP7_75t_SL \i59/i249  (.A(\i59/n148 ),
    .B(\i59/n181 ),
    .Y(\i59/n239 ));
 NOR2xp33_ASAP7_75t_SL \i59/i25  (.A(\i59/n428 ),
    .B(\i59/n451 ),
    .Y(\i59/n469 ));
 OAI22xp5_ASAP7_75t_SL \i59/i250  (.A1(\i59/n84 ),
    .A2(\i59/n58 ),
    .B1(\i59/n78 ),
    .B2(\i59/n39 ),
    .Y(\i59/n238 ));
 OAI21xp5_ASAP7_75t_SL \i59/i251  (.A1(\i59/n52 ),
    .A2(\i59/n49 ),
    .B(\i59/n543 ),
    .Y(\i59/n237 ));
 OAI21xp5_ASAP7_75t_SL \i59/i252  (.A1(\i59/n52 ),
    .A2(\i59/n59 ),
    .B(\i59/n7 ),
    .Y(\i59/n262 ));
 OAI21xp5_ASAP7_75t_SL \i59/i253  (.A1(\i59/n82 ),
    .A2(\i59/n66 ),
    .B(\i59/n200 ),
    .Y(\i59/n261 ));
 AOI22xp5_ASAP7_75t_SL \i59/i254  (.A1(\i59/n47 ),
    .A2(\i59/n63 ),
    .B1(\i59/n51 ),
    .B2(\i59/n61 ),
    .Y(\i59/n260 ));
 AOI22xp5_ASAP7_75t_SL \i59/i255  (.A1(\i59/n63 ),
    .A2(\i59/n57 ),
    .B1(\i59/n45 ),
    .B2(\i59/n50 ),
    .Y(\i59/n258 ));
 OAI22xp5_ASAP7_75t_SL \i59/i256  (.A1(\i59/n68 ),
    .A2(\i59/n60 ),
    .B1(\i59/n525 ),
    .B2(\i59/n66 ),
    .Y(\i59/n256 ));
 AO22x1_ASAP7_75t_SL \i59/i257  (.A1(\i59/n504 ),
    .A2(\i59/n57 ),
    .B1(\i59/n48 ),
    .B2(\i59/n62 ),
    .Y(\i59/n255 ));
 OAI22xp5_ASAP7_75t_SL \i59/i258  (.A1(\i59/n54 ),
    .A2(\i59/n58 ),
    .B1(\i59/n72 ),
    .B2(\i59/n4 ),
    .Y(\i59/n236 ));
 OAI21xp5_ASAP7_75t_SL \i59/i259  (.A1(\i59/n52 ),
    .A2(\i59/n37 ),
    .B(\i59/n9 ),
    .Y(\i59/n253 ));
 NOR2xp33_ASAP7_75t_SL \i59/i26  (.A(\i59/n453 ),
    .B(\i59/n458 ),
    .Y(\i59/n468 ));
 NAND2xp5_ASAP7_75t_SL \i59/i260  (.A(\i59/n42 ),
    .B(\i59/n6 ),
    .Y(\i59/n251 ));
 AOI22xp5_ASAP7_75t_SL \i59/i261  (.A1(\i59/n51 ),
    .A2(\i59/n80 ),
    .B1(\i59/n53 ),
    .B2(\i59/n69 ),
    .Y(\i59/n250 ));
 INVxp67_ASAP7_75t_SL \i59/i262  (.A(\i59/n234 ),
    .Y(\i59/n235 ));
 INVxp67_ASAP7_75t_SL \i59/i263  (.A(\i59/n499 ),
    .Y(\i59/n229 ));
 INVxp67_ASAP7_75t_SL \i59/i264  (.A(\i59/n227 ),
    .Y(\i59/n228 ));
 INVx1_ASAP7_75t_SL \i59/i265  (.A(\i59/n222 ),
    .Y(\i59/n223 ));
 AOI22xp33_ASAP7_75t_SL \i59/i266  (.A1(\i59/n38 ),
    .A2(\i59/n57 ),
    .B1(\i59/n51 ),
    .B2(\i59/n53 ),
    .Y(\i59/n219 ));
 OAI21xp5_ASAP7_75t_SL \i59/i267  (.A1(\i59/n42 ),
    .A2(\i59/n40 ),
    .B(\i59/n50 ),
    .Y(\i59/n218 ));
 AOI21xp33_ASAP7_75t_SL \i59/i268  (.A1(\i59/n64 ),
    .A2(\i59/n76 ),
    .B(\i59/n37 ),
    .Y(\i59/n217 ));
 AOI22xp5_ASAP7_75t_SL \i59/i269  (.A1(\i59/n87 ),
    .A2(\i59/n80 ),
    .B1(\i59/n48 ),
    .B2(\i59/n71 ),
    .Y(\i59/n216 ));
 AND2x2_ASAP7_75t_SL \i59/i27  (.A(\i59/n419 ),
    .B(\i59/n450 ),
    .Y(\i59/n473 ));
 AOI22xp5_ASAP7_75t_SL \i59/i270  (.A1(\i59/n56 ),
    .A2(\i59/n61 ),
    .B1(\i59/n77 ),
    .B2(\i59/n504 ),
    .Y(\i59/n215 ));
 AOI22xp5_ASAP7_75t_SL \i59/i271  (.A1(\i59/n87 ),
    .A2(\i59/n61 ),
    .B1(\i59/n83 ),
    .B2(\i59/n42 ),
    .Y(\i59/n234 ));
 OAI22xp5_ASAP7_75t_SL \i59/i272  (.A1(\i59/n525 ),
    .A2(\i59/n55 ),
    .B1(\i59/n52 ),
    .B2(\i59/n487 ),
    .Y(\i59/n214 ));
 OAI21xp5_ASAP7_75t_SL \i59/i273  (.A1(\i59/n84 ),
    .A2(\i59/n39 ),
    .B(\i59/n122 ),
    .Y(\i59/n213 ));
 AOI22xp5_ASAP7_75t_SL \i59/i274  (.A1(\i59/n504 ),
    .A2(\i59/n69 ),
    .B1(\i59/n38 ),
    .B2(\i59/n45 ),
    .Y(\i59/n212 ));
 AOI22xp5_ASAP7_75t_SL \i59/i275  (.A1(\i59/n1 ),
    .A2(\i59/n42 ),
    .B1(\i59/n63 ),
    .B2(\i59/n67 ),
    .Y(\i59/n211 ));
 OAI22xp5_ASAP7_75t_SL \i59/i276  (.A1(\i59/n74 ),
    .A2(\i59/n64 ),
    .B1(\i59/n37 ),
    .B2(\i59/n68 ),
    .Y(\i59/n233 ));
 NAND2xp5_ASAP7_75t_SL \i59/i277  (.A(\i59/n205 ),
    .B(\i59/n531 ),
    .Y(\i59/n210 ));
 AOI22xp5_ASAP7_75t_SL \i59/i278  (.A1(\i59/n48 ),
    .A2(\i59/n65 ),
    .B1(\i59/n45 ),
    .B2(\i59/n1 ),
    .Y(\i59/n232 ));
 NAND2xp5_ASAP7_75t_SL \i59/i279  (.A(\i59/n204 ),
    .B(\i59/n147 ),
    .Y(\i59/n209 ));
 NOR2xp33_ASAP7_75t_SL \i59/i28  (.A(\i59/n457 ),
    .B(\i59/n441 ),
    .Y(\i59/n467 ));
 OAI22xp5_ASAP7_75t_SL \i59/i280  (.A1(\i59/n52 ),
    .A2(\i59/n84 ),
    .B1(\i59/n72 ),
    .B2(\i59/n70 ),
    .Y(\i59/n231 ));
 OAI22xp33_ASAP7_75t_SL \i59/i281  (.A1(\i59/n487 ),
    .A2(\i59/n46 ),
    .B1(\i59/n506 ),
    .B2(\i59/n72 ),
    .Y(\i59/n208 ));
 OAI22xp5_ASAP7_75t_SL \i59/i282  (.A1(\i59/n64 ),
    .A2(\i59/n72 ),
    .B1(\i59/n41 ),
    .B2(\i59/n37 ),
    .Y(\i59/n230 ));
 AOI22xp5_ASAP7_75t_SL \i59/i283  (.A1(\i59/n65 ),
    .A2(\i59/n85 ),
    .B1(\i59/n87 ),
    .B2(\i59/n79 ),
    .Y(\i59/n227 ));
 OAI22xp5_ASAP7_75t_SL \i59/i284  (.A1(\i59/n525 ),
    .A2(\i59/n39 ),
    .B1(\i59/n70 ),
    .B2(\i59/n54 ),
    .Y(\i59/n226 ));
 OAI22xp5_ASAP7_75t_SL \i59/i285  (.A1(\i59/n46 ),
    .A2(\i59/n509 ),
    .B1(\i59/n4 ),
    .B2(\i59/n37 ),
    .Y(\i59/n225 ));
 AOI22xp5_ASAP7_75t_SL \i59/i286  (.A1(\i59/n61 ),
    .A2(\i59/n57 ),
    .B1(\i59/n38 ),
    .B2(\i59/n67 ),
    .Y(\i59/n224 ));
 AOI22xp5_ASAP7_75t_SL \i59/i287  (.A1(\i59/n47 ),
    .A2(\i59/n38 ),
    .B1(\i59/n53 ),
    .B2(\i59/n45 ),
    .Y(\i59/n207 ));
 AOI22xp33_ASAP7_75t_SL \i59/i288  (.A1(\i59/n85 ),
    .A2(\i59/n71 ),
    .B1(\i59/n77 ),
    .B2(\i59/n63 ),
    .Y(\i59/n206 ));
 AO22x1_ASAP7_75t_SL \i59/i289  (.A1(\i59/n50 ),
    .A2(\i59/n65 ),
    .B1(\i59/n77 ),
    .B2(\i59/n85 ),
    .Y(\i59/n222 ));
 NOR2xp33_ASAP7_75t_SL \i59/i29  (.A(\i59/n435 ),
    .B(\i59/n440 ),
    .Y(\i59/n466 ));
 AOI22xp5_ASAP7_75t_SL \i59/i290  (.A1(\i59/n40 ),
    .A2(\i59/n61 ),
    .B1(\i59/n79 ),
    .B2(\i59/n77 ),
    .Y(\i59/n221 ));
 AOI22xp5_ASAP7_75t_SL \i59/i291  (.A1(\i59/n69 ),
    .A2(\i59/n81 ),
    .B1(\i59/n73 ),
    .B2(\i59/n56 ),
    .Y(\i59/n220 ));
 INVxp67_ASAP7_75t_SL \i59/i292  (.A(\i59/n531 ),
    .Y(\i59/n201 ));
 INVxp67_ASAP7_75t_SL \i59/i293  (.A(\i59/n198 ),
    .Y(\i59/n199 ));
 INVxp67_ASAP7_75t_SL \i59/i294  (.A(\i59/n196 ),
    .Y(\i59/n197 ));
 INVxp67_ASAP7_75t_SL \i59/i295  (.A(\i59/n497 ),
    .Y(\i59/n195 ));
 INVxp67_ASAP7_75t_SL \i59/i296  (.A(\i59/n548 ),
    .Y(\i59/n194 ));
 INVxp67_ASAP7_75t_SL \i59/i297  (.A(\i59/n186 ),
    .Y(\i59/n187 ));
 INVx1_ASAP7_75t_SL \i59/i298  (.A(\i59/n182 ),
    .Y(\i59/n183 ));
 INVxp67_ASAP7_75t_SL \i59/i299  (.A(\i59/n180 ),
    .Y(\i59/n181 ));
 AND3x2_ASAP7_75t_SL \i59/i3  (.A(\i59/n471 ),
    .B(\i59/n484 ),
    .C(\i59/n551 ),
    .Y(n2[6]));
 NOR2xp33_ASAP7_75t_SL \i59/i30  (.A(\i59/n434 ),
    .B(\i59/n452 ),
    .Y(\i59/n465 ));
 INVxp67_ASAP7_75t_SL \i59/i300  (.A(\i59/n178 ),
    .Y(\i59/n179 ));
 INVx1_ASAP7_75t_SL \i59/i301  (.A(\i59/n176 ),
    .Y(\i59/n177 ));
 NAND2xp5_ASAP7_75t_L \i59/i302  (.A(\i59/n82 ),
    .B(\i59/n74 ),
    .Y(\i59/n174 ));
 NAND2xp5_ASAP7_75t_SL \i59/i303  (.A(\i59/n62 ),
    .B(\i59/n63 ),
    .Y(\i59/n173 ));
 NAND2xp5_ASAP7_75t_SL \i59/i304  (.A(\i59/n80 ),
    .B(\i59/n40 ),
    .Y(\i59/n172 ));
 NAND2xp33_ASAP7_75t_L \i59/i305  (.A(\i59/n84 ),
    .B(\i59/n78 ),
    .Y(\i59/n171 ));
 NAND2xp5_ASAP7_75t_SL \i59/i306  (.A(\i59/n71 ),
    .B(\i59/n63 ),
    .Y(\i59/n170 ));
 NOR2xp33_ASAP7_75t_L \i59/i307  (.A(\i59/n45 ),
    .B(\i59/n62 ),
    .Y(\i59/n169 ));
 NAND2xp5_ASAP7_75t_SL \i59/i308  (.A(\i59/n49 ),
    .B(\i59/n2 ),
    .Y(\i59/n168 ));
 NAND2xp5_ASAP7_75t_SL \i59/i309  (.A(\i59/n60 ),
    .B(\i59/n2 ),
    .Y(\i59/n167 ));
 AND4x1_ASAP7_75t_SL \i59/i31  (.A(\i59/n424 ),
    .B(\i59/n420 ),
    .C(\i59/n382 ),
    .D(\i59/n375 ),
    .Y(\i59/n464 ));
 NAND2xp5_ASAP7_75t_SL \i59/i310  (.A(\i59/n71 ),
    .B(\i59/n80 ),
    .Y(\i59/n166 ));
 NOR2xp33_ASAP7_75t_SL \i59/i311  (.A(\i59/n79 ),
    .B(\i59/n81 ),
    .Y(\i59/n165 ));
 NOR2xp33_ASAP7_75t_SL \i59/i312  (.A(\i59/n81 ),
    .B(\i59/n63 ),
    .Y(\i59/n164 ));
 NAND2xp5_ASAP7_75t_SL \i59/i313  (.A(\i59/n44 ),
    .B(\i59/n85 ),
    .Y(\i59/n205 ));
 NAND2xp5_ASAP7_75t_SL \i59/i314  (.A(\i59/n56 ),
    .B(\i59/n504 ),
    .Y(\i59/n163 ));
 NAND2xp5_ASAP7_75t_SL \i59/i315  (.A(\i59/n62 ),
    .B(\i59/n50 ),
    .Y(\i59/n162 ));
 NOR2xp33_ASAP7_75t_SL \i59/i316  (.A(\i59/n51 ),
    .B(\i59/n40 ),
    .Y(\i59/n161 ));
 NOR2xp33_ASAP7_75t_SL \i59/i317  (.A(\i59/n65 ),
    .B(\i59/n45 ),
    .Y(\i59/n160 ));
 NOR2xp67_ASAP7_75t_SL \i59/i318  (.A(\i59/n525 ),
    .B(\i59/n70 ),
    .Y(\i59/n159 ));
 NAND2xp5_ASAP7_75t_SL \i59/i319  (.A(\i59/n81 ),
    .B(\i59/n44 ),
    .Y(\i59/n158 ));
 NOR3xp33_ASAP7_75t_SL \i59/i32  (.A(\i59/n405 ),
    .B(\i59/n353 ),
    .C(\i59/n417 ),
    .Y(\i59/n463 ));
 NOR2xp33_ASAP7_75t_SL \i59/i320  (.A(\i59/n65 ),
    .B(\i59/n71 ),
    .Y(\i59/n157 ));
 NOR2xp33_ASAP7_75t_SL \i59/i321  (.A(\i59/n42 ),
    .B(\i59/n65 ),
    .Y(\i59/n156 ));
 NAND2xp5_ASAP7_75t_SL \i59/i322  (.A(\i59/n47 ),
    .B(\i59/n73 ),
    .Y(\i59/n155 ));
 NAND2xp5_ASAP7_75t_SL \i59/i323  (.A(\i59/n77 ),
    .B(\i59/n63 ),
    .Y(\i59/n154 ));
 NAND2xp5_ASAP7_75t_SL \i59/i324  (.A(\i59/n73 ),
    .B(\i59/n45 ),
    .Y(\i59/n204 ));
 NAND2xp5_ASAP7_75t_SL \i59/i325  (.A(\i59/n63 ),
    .B(\i59/n40 ),
    .Y(\i59/n203 ));
 NAND2xp5_ASAP7_75t_SL \i59/i326  (.A(\i59/n77 ),
    .B(\i59/n61 ),
    .Y(\i59/n153 ));
 NAND2xp5_ASAP7_75t_SL \i59/i327  (.A(\i59/n73 ),
    .B(\i59/n67 ),
    .Y(\i59/n152 ));
 NAND2xp5_ASAP7_75t_SL \i59/i328  (.A(\i59/n51 ),
    .B(\i59/n73 ),
    .Y(\i59/n151 ));
 NAND2xp5_ASAP7_75t_SL \i59/i329  (.A(\i59/n62 ),
    .B(\i59/n80 ),
    .Y(\i59/n11 ));
 NAND2xp33_ASAP7_75t_SL \i59/i33  (.A(\i59/n14 ),
    .B(\i59/n436 ),
    .Y(\i59/n462 ));
 NOR2xp33_ASAP7_75t_SL \i59/i330  (.A(\i59/n72 ),
    .B(\i59/n4 ),
    .Y(\i59/n150 ));
 NAND2xp5_ASAP7_75t_SL \i59/i331  (.A(\i59/n1 ),
    .B(\i59/n69 ),
    .Y(\i59/n10 ));
 NAND2xp33_ASAP7_75t_SL \i59/i332  (.A(\i59/n41 ),
    .B(\i59/n76 ),
    .Y(\i59/n202 ));
 NAND2xp5_ASAP7_75t_SL \i59/i333  (.A(\i59/n53 ),
    .B(\i59/n65 ),
    .Y(\i59/n9 ));
 NAND2xp5_ASAP7_75t_SL \i59/i334  (.A(\i59/n77 ),
    .B(\i59/n1 ),
    .Y(\i59/n8 ));
 NOR2xp33_ASAP7_75t_SL \i59/i335  (.A(\i59/n76 ),
    .B(\i59/n74 ),
    .Y(\i59/n149 ));
 NAND2xp5_ASAP7_75t_SL \i59/i336  (.A(\i59/n87 ),
    .B(\i59/n53 ),
    .Y(\i59/n200 ));
 NAND2xp5_ASAP7_75t_L \i59/i337  (.A(\i59/n81 ),
    .B(\i59/n87 ),
    .Y(\i59/n198 ));
 NAND2xp5_ASAP7_75t_SL \i59/i338  (.A(\i59/n69 ),
    .B(\i59/n63 ),
    .Y(\i59/n196 ));
 NOR2x1_ASAP7_75t_SL \i59/i339  (.A(\i59/n73 ),
    .B(\i59/n50 ),
    .Y(\i59/n193 ));
 INVxp67_ASAP7_75t_SL \i59/i34  (.A(\i59/n460 ),
    .Y(\i59/n461 ));
 AND2x2_ASAP7_75t_SL \i59/i340  (.A(\i59/n504 ),
    .B(\i59/n71 ),
    .Y(\i59/n192 ));
 NAND2xp5_ASAP7_75t_SL \i59/i341  (.A(\i59/n73 ),
    .B(\i59/n44 ),
    .Y(\i59/n191 ));
 NOR2xp33_ASAP7_75t_L \i59/i342  (.A(\i59/n42 ),
    .B(\i59/n62 ),
    .Y(\i59/n190 ));
 NAND2xp5_ASAP7_75t_SL \i59/i343  (.A(\i59/n77 ),
    .B(\i59/n80 ),
    .Y(\i59/n189 ));
 NAND2xp5_ASAP7_75t_SL \i59/i344  (.A(\i59/n44 ),
    .B(\i59/n63 ),
    .Y(\i59/n188 ));
 NAND2xp5_ASAP7_75t_SL \i59/i345  (.A(\i59/n47 ),
    .B(\i59/n85 ),
    .Y(\i59/n186 ));
 NAND2xp5_ASAP7_75t_SL \i59/i346  (.A(\i59/n62 ),
    .B(\i59/n38 ),
    .Y(\i59/n185 ));
 NAND2xp5_ASAP7_75t_SL \i59/i347  (.A(\i59/n62 ),
    .B(\i59/n81 ),
    .Y(\i59/n184 ));
 NOR2xp33_ASAP7_75t_SL \i59/i348  (.A(\i59/n509 ),
    .B(\i59/n506 ),
    .Y(\i59/n148 ));
 NOR2xp33_ASAP7_75t_L \i59/i349  (.A(\i59/n38 ),
    .B(\i59/n73 ),
    .Y(\i59/n182 ));
 INVxp67_ASAP7_75t_SL \i59/i35  (.A(\i59/n458 ),
    .Y(\i59/n459 ));
 NAND2xp5_ASAP7_75t_SL \i59/i350  (.A(\i59/n87 ),
    .B(\i59/n1 ),
    .Y(\i59/n180 ));
 NAND2xp33_ASAP7_75t_SL \i59/i351  (.A(\i59/n2 ),
    .B(\i59/n78 ),
    .Y(\i59/n178 ));
 NOR2xp33_ASAP7_75t_L \i59/i352  (.A(\i59/n83 ),
    .B(\i59/n79 ),
    .Y(\i59/n176 ));
 NOR2xp33_ASAP7_75t_SL \i59/i353  (.A(\i59/n83 ),
    .B(\i59/n73 ),
    .Y(\i59/n175 ));
 INVxp67_ASAP7_75t_SL \i59/i354  (.A(\i59/n535 ),
    .Y(\i59/n144 ));
 INVxp67_ASAP7_75t_SL \i59/i355  (.A(\i59/n138 ),
    .Y(\i59/n139 ));
 INVxp67_ASAP7_75t_SL \i59/i356  (.A(\i59/n132 ),
    .Y(\i59/n133 ));
 INVxp67_ASAP7_75t_SL \i59/i357  (.A(\i59/n129 ),
    .Y(\i59/n130 ));
 INVxp67_ASAP7_75t_SL \i59/i358  (.A(\i59/n5 ),
    .Y(\i59/n126 ));
 NOR2xp33_ASAP7_75t_SL \i59/i359  (.A(\i59/n42 ),
    .B(\i59/n56 ),
    .Y(\i59/n125 ));
 NAND3xp33_ASAP7_75t_SL \i59/i36  (.A(\i59/n413 ),
    .B(\i59/n368 ),
    .C(\i59/n374 ),
    .Y(\i59/n456 ));
 NOR2xp33_ASAP7_75t_SL \i59/i360  (.A(\i59/n82 ),
    .B(\i59/n486 ),
    .Y(\i59/n124 ));
 NAND2xp33_ASAP7_75t_SL \i59/i361  (.A(\i59/n54 ),
    .B(\i59/n78 ),
    .Y(\i59/n123 ));
 NAND2xp5_ASAP7_75t_SL \i59/i362  (.A(\i59/n42 ),
    .B(\i59/n81 ),
    .Y(\i59/n122 ));
 NAND2xp5_ASAP7_75t_SL \i59/i363  (.A(\i59/n83 ),
    .B(\i59/n40 ),
    .Y(\i59/n121 ));
 NOR2xp33_ASAP7_75t_SL \i59/i364  (.A(\i59/n83 ),
    .B(\i59/n50 ),
    .Y(\i59/n120 ));
 NAND2xp5_ASAP7_75t_SL \i59/i365  (.A(\i59/n47 ),
    .B(\i59/n38 ),
    .Y(\i59/n119 ));
 NAND2xp33_ASAP7_75t_L \i59/i366  (.A(\i59/n58 ),
    .B(\i59/n55 ),
    .Y(\i59/n118 ));
 NAND2xp33_ASAP7_75t_SL \i59/i367  (.A(\i59/n59 ),
    .B(\i59/n54 ),
    .Y(\i59/n117 ));
 NOR2xp33_ASAP7_75t_SL \i59/i368  (.A(\i59/n47 ),
    .B(\i59/n44 ),
    .Y(\i59/n116 ));
 NOR2xp33_ASAP7_75t_SL \i59/i369  (.A(\i59/n1 ),
    .B(\i59/n38 ),
    .Y(\i59/n115 ));
 NAND2xp5_ASAP7_75t_L \i59/i37  (.A(\i59/n552 ),
    .B(\i59/n393 ),
    .Y(\i59/n455 ));
 NAND2xp5_ASAP7_75t_SL \i59/i370  (.A(\i59/n75 ),
    .B(\i59/n47 ),
    .Y(\i59/n114 ));
 NOR2xp33_ASAP7_75t_L \i59/i371  (.A(\i59/n47 ),
    .B(\i59/n67 ),
    .Y(\i59/n113 ));
 NAND2xp5_ASAP7_75t_SL \i59/i372  (.A(\i59/n47 ),
    .B(\i59/n50 ),
    .Y(\i59/n112 ));
 NAND2xp5_ASAP7_75t_SL \i59/i373  (.A(\i59/n1 ),
    .B(\i59/n56 ),
    .Y(\i59/n111 ));
 NAND2xp5_ASAP7_75t_SL \i59/i374  (.A(\i59/n47 ),
    .B(\i59/n79 ),
    .Y(\i59/n110 ));
 NAND2xp33_ASAP7_75t_SL \i59/i375  (.A(\i59/n41 ),
    .B(\i59/n68 ),
    .Y(\i59/n109 ));
 NAND2xp33_ASAP7_75t_SL \i59/i376  (.A(\i59/n74 ),
    .B(\i59/n70 ),
    .Y(\i59/n108 ));
 NOR2xp33_ASAP7_75t_SL \i59/i377  (.A(\i59/n44 ),
    .B(\i59/n69 ),
    .Y(\i59/n107 ));
 NAND2xp33_ASAP7_75t_L \i59/i378  (.A(\i59/n43 ),
    .B(\i59/n52 ),
    .Y(\i59/n106 ));
 NAND2xp5_ASAP7_75t_SL \i59/i379  (.A(\i59/n44 ),
    .B(\i59/n61 ),
    .Y(\i59/n147 ));
 NOR2xp33_ASAP7_75t_SL \i59/i38  (.A(\i59/n421 ),
    .B(\i59/n351 ),
    .Y(\i59/n454 ));
 NAND2xp33_ASAP7_75t_SL \i59/i380  (.A(\i59/n486 ),
    .B(\i59/n43 ),
    .Y(\i59/n105 ));
 NAND2xp5_ASAP7_75t_SL \i59/i381  (.A(\i59/n50 ),
    .B(\i59/n71 ),
    .Y(\i59/n104 ));
 NAND2xp5_ASAP7_75t_SL \i59/i382  (.A(\i59/n44 ),
    .B(\i59/n48 ),
    .Y(\i59/n146 ));
 NOR2xp33_ASAP7_75t_SL \i59/i383  (.A(\i59/n509 ),
    .B(\i59/n68 ),
    .Y(\i59/n103 ));
 NOR2xp33_ASAP7_75t_SL \i59/i384  (.A(\i59/n56 ),
    .B(\i59/n40 ),
    .Y(\i59/n102 ));
 NAND2xp33_ASAP7_75t_SL \i59/i385  (.A(\i59/n486 ),
    .B(\i59/n66 ),
    .Y(\i59/n101 ));
 NAND2xp5_ASAP7_75t_SL \i59/i386  (.A(\i59/n53 ),
    .B(\i59/n45 ),
    .Y(\i59/n100 ));
 NOR2xp33_ASAP7_75t_SL \i59/i387  (.A(\i59/n53 ),
    .B(\i59/n38 ),
    .Y(\i59/n99 ));
 NAND2xp5_ASAP7_75t_L \i59/i388  (.A(\i59/n54 ),
    .B(\i59/n74 ),
    .Y(\i59/n98 ));
 NAND2xp5_ASAP7_75t_SL \i59/i389  (.A(\i59/n79 ),
    .B(\i59/n67 ),
    .Y(\i59/n97 ));
 NAND2xp33_ASAP7_75t_SL \i59/i39  (.A(\i59/n415 ),
    .B(\i59/n398 ),
    .Y(\i59/n453 ));
 NAND2xp5_ASAP7_75t_SL \i59/i390  (.A(\i59/n50 ),
    .B(\i59/n69 ),
    .Y(\i59/n145 ));
 NOR2xp33_ASAP7_75t_SL \i59/i391  (.A(\i59/n54 ),
    .B(\i59/n68 ),
    .Y(\i59/n96 ));
 NAND2xp5_ASAP7_75t_SL \i59/i392  (.A(\i59/n48 ),
    .B(\i59/n57 ),
    .Y(\i59/n95 ));
 NOR2xp33_ASAP7_75t_SL \i59/i393  (.A(\i59/n78 ),
    .B(\i59/n39 ),
    .Y(\i59/n94 ));
 NOR2xp33_ASAP7_75t_SL \i59/i394  (.A(\i59/n525 ),
    .B(\i59/n66 ),
    .Y(\i59/n93 ));
 NAND2xp5_ASAP7_75t_SL \i59/i395  (.A(\i59/n51 ),
    .B(\i59/n79 ),
    .Y(\i59/n143 ));
 NAND2xp5_ASAP7_75t_SL \i59/i396  (.A(\i59/n61 ),
    .B(\i59/n71 ),
    .Y(\i59/n7 ));
 NAND2x1p5_ASAP7_75t_SL \i59/i397  (.A(\i59/n74 ),
    .B(\i59/n78 ),
    .Y(\i59/n6 ));
 NOR2xp33_ASAP7_75t_L \i59/i398  (.A(\i59/n1 ),
    .B(\i59/n75 ),
    .Y(\i59/n142 ));
 NAND2xp5_ASAP7_75t_SL \i59/i399  (.A(\i59/n75 ),
    .B(\i59/n40 ),
    .Y(\i59/n141 ));
 AND2x4_ASAP7_75t_SL \i59/i4  (.A(\i59/n482 ),
    .B(\i59/n474 ),
    .Y(n2[3]));
 NAND3xp33_ASAP7_75t_SL \i59/i40  (.A(\i59/n426 ),
    .B(\i59/n267 ),
    .C(\i59/n540 ),
    .Y(\i59/n452 ));
 NAND2xp5_ASAP7_75t_SL \i59/i400  (.A(\i59/n53 ),
    .B(\i59/n40 ),
    .Y(\i59/n140 ));
 NOR2xp33_ASAP7_75t_SL \i59/i401  (.A(\i59/n52 ),
    .B(\i59/n60 ),
    .Y(\i59/n92 ));
 NAND2xp5_ASAP7_75t_SL \i59/i402  (.A(\i59/n51 ),
    .B(\i59/n83 ),
    .Y(\i59/n91 ));
 NAND2xp5_ASAP7_75t_SL \i59/i403  (.A(\i59/n38 ),
    .B(\i59/n57 ),
    .Y(\i59/n90 ));
 NAND2xp5_ASAP7_75t_SL \i59/i404  (.A(\i59/n48 ),
    .B(\i59/n45 ),
    .Y(\i59/n138 ));
 NAND2xp5_ASAP7_75t_SL \i59/i405  (.A(\i59/n48 ),
    .B(\i59/n67 ),
    .Y(\i59/n137 ));
 NAND2xp5_ASAP7_75t_SL \i59/i406  (.A(\i59/n61 ),
    .B(\i59/n45 ),
    .Y(\i59/n136 ));
 NOR2xp33_ASAP7_75t_SL \i59/i407  (.A(\i59/n486 ),
    .B(\i59/n49 ),
    .Y(\i59/n89 ));
 NAND2xp5_ASAP7_75t_SL \i59/i408  (.A(\i59/n38 ),
    .B(\i59/n56 ),
    .Y(\i59/n135 ));
 NAND2xp5_ASAP7_75t_SL \i59/i409  (.A(\i59/n50 ),
    .B(\i59/n56 ),
    .Y(\i59/n134 ));
 NAND2xp33_ASAP7_75t_SL \i59/i41  (.A(\i59/n408 ),
    .B(\i59/n412 ),
    .Y(\i59/n451 ));
 AND2x2_ASAP7_75t_SL \i59/i410  (.A(\i59/n53 ),
    .B(\i59/n42 ),
    .Y(\i59/n132 ));
 NAND4xp25_ASAP7_75t_SL \i59/i411  (.A(\i59/n32 ),
    .B(\i59/n34 ),
    .C(\i59/n23 ),
    .D(\i59/n24 ),
    .Y(\i59/n131 ));
 NAND2xp5_ASAP7_75t_SL \i59/i412  (.A(\i59/n44 ),
    .B(\i59/n38 ),
    .Y(\i59/n129 ));
 NAND2xp5_ASAP7_75t_SL \i59/i413  (.A(\i59/n47 ),
    .B(\i59/n61 ),
    .Y(\i59/n88 ));
 AND2x2_ASAP7_75t_SL \i59/i414  (.A(\i59/n50 ),
    .B(\i59/n42 ),
    .Y(\i59/n128 ));
 AND2x2_ASAP7_75t_SL \i59/i415  (.A(\i59/n48 ),
    .B(\i59/n56 ),
    .Y(\i59/n127 ));
 NAND2xp5_ASAP7_75t_SL \i59/i416  (.A(\i59/n81 ),
    .B(\i59/n56 ),
    .Y(\i59/n5 ));
 INVx2_ASAP7_75t_SL \i59/i417  (.A(\i59/n87 ),
    .Y(\i59/n86 ));
 INVx2_ASAP7_75t_SL \i59/i418  (.A(\i59/n85 ),
    .Y(\i59/n84 ));
 INVx4_ASAP7_75t_SL \i59/i419  (.A(\i59/n83 ),
    .Y(\i59/n82 ));
 NOR2xp33_ASAP7_75t_SL \i59/i42  (.A(\i59/n410 ),
    .B(\i59/n409 ),
    .Y(\i59/n450 ));
 INVx3_ASAP7_75t_SL \i59/i420  (.A(\i59/n79 ),
    .Y(\i59/n78 ));
 INVx2_ASAP7_75t_SL \i59/i421  (.A(\i59/n77 ),
    .Y(\i59/n76 ));
 INVx3_ASAP7_75t_SL \i59/i422  (.A(\i59/n75 ),
    .Y(\i59/n74 ));
 INVx2_ASAP7_75t_SL \i59/i423  (.A(\i59/n73 ),
    .Y(\i59/n72 ));
 INVx2_ASAP7_75t_SL \i59/i424  (.A(\i59/n71 ),
    .Y(\i59/n70 ));
 INVx2_ASAP7_75t_SL \i59/i425  (.A(\i59/n69 ),
    .Y(\i59/n68 ));
 INVx2_ASAP7_75t_SL \i59/i426  (.A(\i59/n67 ),
    .Y(\i59/n66 ));
 INVx3_ASAP7_75t_SL \i59/i427  (.A(\i59/n65 ),
    .Y(\i59/n64 ));
 AND2x4_ASAP7_75t_SL \i59/i428  (.A(\i59/n28 ),
    .B(\i59/n30 ),
    .Y(\i59/n87 ));
 AND2x4_ASAP7_75t_SL \i59/i429  (.A(\i59/n522 ),
    .B(\i59/n23 ),
    .Y(\i59/n85 ));
 NAND4xp25_ASAP7_75t_L \i59/i43  (.A(\i59/n388 ),
    .B(\i59/n327 ),
    .C(\i59/n249 ),
    .D(\i59/n290 ),
    .Y(\i59/n449 ));
 AND2x4_ASAP7_75t_SL \i59/i430  (.A(\i59/n35 ),
    .B(\i59/n521 ),
    .Y(\i59/n83 ));
 AND2x4_ASAP7_75t_SL \i59/i431  (.A(\i59/n36 ),
    .B(\i59/n24 ),
    .Y(\i59/n81 ));
 AND2x4_ASAP7_75t_SL \i59/i432  (.A(\i59/n25 ),
    .B(\i59/n23 ),
    .Y(\i59/n80 ));
 AND2x4_ASAP7_75t_SL \i59/i433  (.A(\i59/n554 ),
    .B(\i59/n24 ),
    .Y(\i59/n79 ));
 AND2x4_ASAP7_75t_SL \i59/i434  (.A(\i59/n536 ),
    .B(\i59/n33 ),
    .Y(\i59/n77 ));
 NAND2x1_ASAP7_75t_SL \i59/i435  (.A(\i59/n536 ),
    .B(\i59/n537 ),
    .Y(\i59/n4 ));
 AND2x4_ASAP7_75t_SL \i59/i436  (.A(\i59/n521 ),
    .B(\i59/n25 ),
    .Y(\i59/n75 ));
 AND2x4_ASAP7_75t_SL \i59/i437  (.A(\i59/n521 ),
    .B(\i59/n24 ),
    .Y(\i59/n73 ));
 AND2x4_ASAP7_75t_SL \i59/i438  (.A(\i59/n536 ),
    .B(\i59/n26 ),
    .Y(\i59/n71 ));
 AND2x4_ASAP7_75t_SL \i59/i439  (.A(\i59/n32 ),
    .B(\i59/n537 ),
    .Y(\i59/n69 ));
 NOR2xp33_ASAP7_75t_SL \i59/i44  (.A(\i59/n425 ),
    .B(\i59/n402 ),
    .Y(\i59/n448 ));
 AND2x4_ASAP7_75t_SL \i59/i440  (.A(\i59/n536 ),
    .B(\i59/n34 ),
    .Y(\i59/n67 ));
 AND2x4_ASAP7_75t_SL \i59/i441  (.A(\i59/n32 ),
    .B(\i59/n34 ),
    .Y(\i59/n65 ));
 INVx2_ASAP7_75t_SL \i59/i442  (.A(\i59/n61 ),
    .Y(\i59/n60 ));
 INVx2_ASAP7_75t_SL \i59/i443  (.A(\i59/n56 ),
    .Y(\i59/n55 ));
 INVx2_ASAP7_75t_SL \i59/i444  (.A(\i59/n52 ),
    .Y(\i59/n51 ));
 INVx2_ASAP7_75t_SL \i59/i445  (.A(\i59/n50 ),
    .Y(\i59/n49 ));
 INVx3_ASAP7_75t_SL \i59/i446  (.A(\i59/n47 ),
    .Y(\i59/n46 ));
 INVx4_ASAP7_75t_SL \i59/i447  (.A(\i59/n44 ),
    .Y(\i59/n43 ));
 INVx2_ASAP7_75t_SL \i59/i448  (.A(\i59/n42 ),
    .Y(\i59/n41 ));
 INVx3_ASAP7_75t_SL \i59/i449  (.A(\i59/n40 ),
    .Y(\i59/n39 ));
 NAND3xp33_ASAP7_75t_SL \i59/i45  (.A(\i59/n371 ),
    .B(\i59/n362 ),
    .C(\i59/n540 ),
    .Y(\i59/n447 ));
 INVx3_ASAP7_75t_SL \i59/i450  (.A(\i59/n38 ),
    .Y(\i59/n37 ));
 AND2x4_ASAP7_75t_SL \i59/i451  (.A(\i59/n25 ),
    .B(\i59/n36 ),
    .Y(\i59/n63 ));
 AND2x4_ASAP7_75t_SL \i59/i452  (.A(\i59/n21 ),
    .B(\i59/n33 ),
    .Y(\i59/n62 ));
 AND2x4_ASAP7_75t_SL \i59/i453  (.A(\i59/n24 ),
    .B(\i59/n23 ),
    .Y(\i59/n61 ));
 NAND2x1p5_ASAP7_75t_SL \i59/i454  (.A(\i59/n554 ),
    .B(\i59/n25 ),
    .Y(\i59/n59 ));
 AND2x4_ASAP7_75t_SL \i59/i455  (.A(\i59/n32 ),
    .B(\i59/n26 ),
    .Y(\i59/n57 ));
 AND2x4_ASAP7_75t_SL \i59/i456  (.A(\i59/n27 ),
    .B(\i59/n537 ),
    .Y(\i59/n56 ));
 NAND2xp5_ASAP7_75t_SL \i59/i457  (.A(\i59/n36 ),
    .B(\i59/n522 ),
    .Y(\i59/n54 ));
 AND4x1_ASAP7_75t_SL \i59/i458  (.A(n3[6]),
    .B(\i59/n0 ),
    .C(\i59/n3 ),
    .D(n3[4]),
    .Y(\i59/n53 ));
 OR2x6_ASAP7_75t_SL \i59/i459  (.A(\i59/n29 ),
    .B(\i59/n22 ),
    .Y(\i59/n52 ));
 NAND3xp33_ASAP7_75t_R \i59/i46  (.A(\i59/n388 ),
    .B(\i59/n372 ),
    .C(\i59/n359 ),
    .Y(\i59/n446 ));
 AND2x4_ASAP7_75t_SL \i59/i460  (.A(\i59/n36 ),
    .B(\i59/n35 ),
    .Y(\i59/n50 ));
 AND2x4_ASAP7_75t_SL \i59/i461  (.A(\i59/n522 ),
    .B(\i59/n554 ),
    .Y(\i59/n48 ));
 AND2x4_ASAP7_75t_SL \i59/i462  (.A(\i59/n31 ),
    .B(\i59/n28 ),
    .Y(\i59/n47 ));
 AND2x4_ASAP7_75t_SL \i59/i463  (.A(\i59/n20 ),
    .B(\i59/n26 ),
    .Y(\i59/n45 ));
 AND2x4_ASAP7_75t_SL \i59/i464  (.A(\i59/n33 ),
    .B(\i59/n27 ),
    .Y(\i59/n44 ));
 AND2x4_ASAP7_75t_SL \i59/i465  (.A(\i59/n33 ),
    .B(\i59/n32 ),
    .Y(\i59/n42 ));
 AND2x4_ASAP7_75t_SL \i59/i466  (.A(\i59/n34 ),
    .B(\i59/n27 ),
    .Y(\i59/n40 ));
 AND2x4_ASAP7_75t_SL \i59/i467  (.A(\i59/n35 ),
    .B(\i59/n554 ),
    .Y(\i59/n38 ));
 AND2x2_ASAP7_75t_SL \i59/i468  (.A(n3[1]),
    .B(n3[0]),
    .Y(\i59/n31 ));
 AND2x2_ASAP7_75t_SL \i59/i469  (.A(n3[6]),
    .B(\i59/n3 ),
    .Y(\i59/n36 ));
 NOR3xp33_ASAP7_75t_SL \i59/i47  (.A(\i59/n340 ),
    .B(\i59/n530 ),
    .C(\i59/n377 ),
    .Y(\i59/n460 ));
 AND2x2_ASAP7_75t_SL \i59/i470  (.A(n3[5]),
    .B(\i59/n17 ),
    .Y(\i59/n35 ));
 AND2x2_ASAP7_75t_SL \i59/i471  (.A(\i59/n19 ),
    .B(\i59/n16 ),
    .Y(\i59/n34 ));
 AND2x2_ASAP7_75t_SL \i59/i472  (.A(n3[3]),
    .B(n3[1]),
    .Y(\i59/n33 ));
 AND2x4_ASAP7_75t_L \i59/i473  (.A(\i59/n18 ),
    .B(\i59/n15 ),
    .Y(\i59/n32 ));
 INVx1_ASAP7_75t_SL \i59/i474  (.A(\i59/n29 ),
    .Y(\i59/n30 ));
 INVx3_ASAP7_75t_SL \i59/i475  (.A(\i59/n494 ),
    .Y(\i59/n23 ));
 NAND2xp5_ASAP7_75t_SL \i59/i476  (.A(n3[3]),
    .B(\i59/n18 ),
    .Y(\i59/n22 ));
 NOR2xp33_ASAP7_75t_SL \i59/i477  (.A(\i59/n15 ),
    .B(n3[2]),
    .Y(\i59/n21 ));
 NOR2xp33_ASAP7_75t_SL \i59/i478  (.A(\i59/n18 ),
    .B(n3[0]),
    .Y(\i59/n20 ));
 OR2x2_ASAP7_75t_SL \i59/i479  (.A(\i59/n15 ),
    .B(n3[1]),
    .Y(\i59/n29 ));
 NAND2xp5_ASAP7_75t_SL \i59/i48  (.A(\i59/n357 ),
    .B(\i59/n426 ),
    .Y(\i59/n458 ));
 AND2x2_ASAP7_75t_SL \i59/i480  (.A(\i59/n19 ),
    .B(\i59/n18 ),
    .Y(\i59/n28 ));
 AND2x2_ASAP7_75t_SL \i59/i481  (.A(n3[2]),
    .B(\i59/n15 ),
    .Y(\i59/n27 ));
 AND2x2_ASAP7_75t_SL \i59/i482  (.A(n3[3]),
    .B(\i59/n16 ),
    .Y(\i59/n26 ));
 AND2x2_ASAP7_75t_SL \i59/i483  (.A(\i59/n0 ),
    .B(\i59/n17 ),
    .Y(\i59/n25 ));
 AND2x2_ASAP7_75t_SL \i59/i484  (.A(n3[5]),
    .B(n3[4]),
    .Y(\i59/n24 ));
 INVx3_ASAP7_75t_SL \i59/i485  (.A(n3[7]),
    .Y(\i59/n3 ));
 INVx2_ASAP7_75t_SL \i59/i486  (.A(n3[3]),
    .Y(\i59/n19 ));
 INVx4_ASAP7_75t_SL \i59/i487  (.A(n3[2]),
    .Y(\i59/n18 ));
 INVx2_ASAP7_75t_SL \i59/i488  (.A(n3[4]),
    .Y(\i59/n17 ));
 INVx2_ASAP7_75t_SL \i59/i489  (.A(n3[1]),
    .Y(\i59/n16 ));
 NAND2xp5_ASAP7_75t_SL \i59/i49  (.A(\i59/n371 ),
    .B(\i59/n400 ),
    .Y(\i59/n457 ));
 INVx3_ASAP7_75t_SL \i59/i490  (.A(n3[0]),
    .Y(\i59/n15 ));
 OAI211xp5_ASAP7_75t_SL \i59/i491  (.A1(\i59/n496 ),
    .A2(\i59/n156 ),
    .B(\i59/n10 ),
    .C(\i59/n184 ),
    .Y(\i59/n485 ));
 INVx6_ASAP7_75t_SL \i59/i492  (.A(\i59/n57 ),
    .Y(\i59/n58 ));
 INVx3_ASAP7_75t_SL \i59/i493  (.A(\i59/n45 ),
    .Y(\i59/n486 ));
 INVx3_ASAP7_75t_SL \i59/i494  (.A(\i59/n81 ),
    .Y(\i59/n487 ));
 NOR4xp25_ASAP7_75t_SL \i59/i495  (.A(\i59/n380 ),
    .B(\i59/n340 ),
    .C(\i59/n228 ),
    .D(\i59/n488 ),
    .Y(\i59/n489 ));
 OAI211xp5_ASAP7_75t_SL \i59/i496  (.A1(\i59/n66 ),
    .A2(\i59/n496 ),
    .B(\i59/n191 ),
    .C(\i59/n532 ),
    .Y(\i59/n490 ));
 OAI22x1_ASAP7_75t_SL \i59/i497  (.A1(\i59/n2 ),
    .A2(\i59/n58 ),
    .B1(\i59/n486 ),
    .B2(\i59/n487 ),
    .Y(\i59/n488 ));
 OAI21xp5_ASAP7_75t_SL \i59/i498  (.A1(\i59/n52 ),
    .A2(\i59/n525 ),
    .B(\i59/n491 ),
    .Y(\i59/n492 ));
 NOR2x1_ASAP7_75t_SL \i59/i499  (.A(\i59/n505 ),
    .B(\i59/n488 ),
    .Y(\i59/n491 ));
 AND3x4_ASAP7_75t_SL \i59/i5  (.A(\i59/n551 ),
    .B(\i59/n476 ),
    .C(\i59/n473 ),
    .Y(n2[4]));
 INVx1_ASAP7_75t_SL \i59/i50  (.A(\i59/n519 ),
    .Y(\i59/n445 ));
 NAND5xp2_ASAP7_75t_SL \i59/i500  (.A(\i59/n366 ),
    .B(\i59/n336 ),
    .C(\i59/n309 ),
    .D(\i59/n307 ),
    .E(\i59/n491 ),
    .Y(\i59/n493 ));
 OR2x2_ASAP7_75t_SL \i59/i501  (.A(n3[7]),
    .B(n3[6]),
    .Y(\i59/n494 ));
 NAND2xp33_ASAP7_75t_SL \i59/i502  (.A(\i59/n509 ),
    .B(\i59/n496 ),
    .Y(\i59/n497 ));
 OR2x6_ASAP7_75t_SL \i59/i503  (.A(\i59/n495 ),
    .B(\i59/n494 ),
    .Y(\i59/n496 ));
 INVx2_ASAP7_75t_SL \i59/i504  (.A(\i59/n35 ),
    .Y(\i59/n495 ));
 NOR2xp67_ASAP7_75t_L \i59/i505  (.A(\i59/n496 ),
    .B(\i59/n4 ),
    .Y(\i59/n498 ));
 OAI22xp5_ASAP7_75t_SL \i59/i506  (.A1(\i59/n52 ),
    .A2(\i59/n496 ),
    .B1(\i59/n86 ),
    .B2(\i59/n72 ),
    .Y(\i59/n499 ));
 OAI22xp5_ASAP7_75t_SL \i59/i507  (.A1(\i59/n509 ),
    .A2(\i59/n39 ),
    .B1(\i59/n46 ),
    .B2(\i59/n496 ),
    .Y(\i59/n500 ));
 OAI22xp5_ASAP7_75t_SL \i59/i508  (.A1(\i59/n496 ),
    .A2(\i59/n64 ),
    .B1(\i59/n72 ),
    .B2(\i59/n39 ),
    .Y(\i59/n501 ));
 OAI22xp5_ASAP7_75t_SL \i59/i509  (.A1(\i59/n496 ),
    .A2(\i59/n169 ),
    .B1(\i59/n82 ),
    .B2(\i59/n64 ),
    .Y(\i59/n502 ));
 INVxp67_ASAP7_75t_SL \i59/i51  (.A(\i59/n443 ),
    .Y(\i59/n444 ));
 OAI222xp33_ASAP7_75t_SL \i59/i510  (.A1(\i59/n72 ),
    .A2(\i59/n76 ),
    .B1(\i59/n39 ),
    .B2(\i59/n496 ),
    .C1(\i59/n37 ),
    .C2(\i59/n86 ),
    .Y(\i59/n503 ));
 INVx3_ASAP7_75t_SL \i59/i511  (.A(\i59/n496 ),
    .Y(\i59/n504 ));
 OAI22xp5_ASAP7_75t_SL \i59/i512  (.A1(\i59/n43 ),
    .A2(\i59/n496 ),
    .B1(\i59/n82 ),
    .B2(\i59/n46 ),
    .Y(\i59/n505 ));
 INVx2_ASAP7_75t_SL \i59/i513  (.A(\i59/n62 ),
    .Y(\i59/n506 ));
 NAND2x1_ASAP7_75t_SL \i59/i514  (.A(\i59/n39 ),
    .B(\i59/n506 ),
    .Y(\i59/n507 ));
 NAND2xp5_ASAP7_75t_SL \i59/i515  (.A(\i59/n83 ),
    .B(\i59/n507 ),
    .Y(\i59/n508 ));
 INVx3_ASAP7_75t_SL \i59/i516  (.A(\i59/n48 ),
    .Y(\i59/n509 ));
 INVx2_ASAP7_75t_SL \i59/i517  (.A(\i59/n63 ),
    .Y(\i59/n510 ));
 NAND2xp5_ASAP7_75t_SL \i59/i518  (.A(\i59/n87 ),
    .B(\i59/n511 ),
    .Y(\i59/n512 ));
 NAND2x1_ASAP7_75t_SL \i59/i519  (.A(\i59/n509 ),
    .B(\i59/n510 ),
    .Y(\i59/n511 ));
 NAND3xp33_ASAP7_75t_L \i59/i52  (.A(\i59/n383 ),
    .B(\i59/n348 ),
    .C(\i59/n394 ),
    .Y(\i59/n442 ));
 AOI221xp5_ASAP7_75t_SL \i59/i520  (.A1(\i59/n511 ),
    .A2(\i59/n77 ),
    .B1(\i59/n63 ),
    .B2(\i59/n65 ),
    .C(\i59/n93 ),
    .Y(\i59/n513 ));
 OAI22xp5_ASAP7_75t_SL \i59/i521  (.A1(\i59/n86 ),
    .A2(\i59/n84 ),
    .B1(\i59/n41 ),
    .B2(\i59/n60 ),
    .Y(\i59/n514 ));
 AND2x2_ASAP7_75t_SL \i59/i522  (.A(\i59/n42 ),
    .B(\i59/n85 ),
    .Y(\i59/n515 ));
 NAND3xp33_ASAP7_75t_SL \i59/i523  (.A(\i59/n517 ),
    .B(\i59/n355 ),
    .C(\i59/n332 ),
    .Y(\i59/n518 ));
 NOR3xp33_ASAP7_75t_SL \i59/i524  (.A(\i59/n514 ),
    .B(\i59/n516 ),
    .C(\i59/n515 ),
    .Y(\i59/n517 ));
 OAI22xp5_ASAP7_75t_SL \i59/i525  (.A1(\i59/n37 ),
    .A2(\i59/n64 ),
    .B1(\i59/n506 ),
    .B2(\i59/n60 ),
    .Y(\i59/n516 ));
 NAND4xp25_ASAP7_75t_SL \i59/i526  (.A(\i59/n394 ),
    .B(\i59/n517 ),
    .C(\i59/n397 ),
    .D(\i59/n321 ),
    .Y(\i59/n519 ));
 NAND2xp5_ASAP7_75t_SL \i59/i527  (.A(\i59/n517 ),
    .B(\i59/n397 ),
    .Y(\i59/n520 ));
 AND2x2_ASAP7_75t_SL \i59/i528  (.A(n3[7]),
    .B(n3[6]),
    .Y(\i59/n521 ));
 AND2x4_ASAP7_75t_SL \i59/i529  (.A(n3[4]),
    .B(\i59/n0 ),
    .Y(\i59/n522 ));
 NAND3xp33_ASAP7_75t_L \i59/i53  (.A(\i59/n391 ),
    .B(\i59/n188 ),
    .C(\i59/n14 ),
    .Y(\i59/n441 ));
 OAI31xp33_ASAP7_75t_SL \i59/i530  (.A1(\i59/n507 ),
    .A2(\i59/n71 ),
    .A3(\i59/n57 ),
    .B(\i59/n523 ),
    .Y(\i59/n524 ));
 AND2x4_ASAP7_75t_SL \i59/i531  (.A(\i59/n521 ),
    .B(\i59/n522 ),
    .Y(\i59/n523 ));
 INVx3_ASAP7_75t_SL \i59/i532  (.A(\i59/n523 ),
    .Y(\i59/n525 ));
 AOI222xp33_ASAP7_75t_SL \i59/i533  (.A1(\i59/n56 ),
    .A2(\i59/n98 ),
    .B1(\i59/n69 ),
    .B2(\i59/n523 ),
    .C1(\i59/n71 ),
    .C2(\i59/n38 ),
    .Y(\i59/n526 ));
 AOI222xp33_ASAP7_75t_SL \i59/i534  (.A1(\i59/n69 ),
    .A2(\i59/n75 ),
    .B1(\i59/n57 ),
    .B2(\i59/n523 ),
    .C1(\i59/n45 ),
    .C2(\i59/n79 ),
    .Y(\i59/n527 ));
 AOI22xp5_ASAP7_75t_SL \i59/i535  (.A1(\i59/n80 ),
    .A2(\i59/n67 ),
    .B1(\i59/n523 ),
    .B2(\i59/n45 ),
    .Y(\i59/n528 ));
 AOI22xp5_ASAP7_75t_SL \i59/i536  (.A1(\i59/n51 ),
    .A2(\i59/n83 ),
    .B1(\i59/n523 ),
    .B2(\i59/n77 ),
    .Y(\i59/n529 ));
 AO22x1_ASAP7_75t_SL \i59/i537  (.A1(\i59/n61 ),
    .A2(\i59/n67 ),
    .B1(\i59/n523 ),
    .B2(\i59/n45 ),
    .Y(\i59/n530 ));
 NAND2xp5_ASAP7_75t_SL \i59/i538  (.A(\i59/n523 ),
    .B(\i59/n65 ),
    .Y(\i59/n531 ));
 NAND2xp5_ASAP7_75t_SL \i59/i539  (.A(\i59/n87 ),
    .B(\i59/n523 ),
    .Y(\i59/n532 ));
 A2O1A1Ixp33_ASAP7_75t_SL \i59/i54  (.A1(\i59/n59 ),
    .A2(\i59/n49 ),
    .B(\i59/n541 ),
    .C(\i59/n401 ),
    .Y(\i59/n440 ));
 NOR2xp33_ASAP7_75t_SL \i59/i540  (.A(\i59/n523 ),
    .B(\i59/n1 ),
    .Y(\i59/n533 ));
 NAND2xp5_ASAP7_75t_SL \i59/i541  (.A(\i59/n47 ),
    .B(\i59/n523 ),
    .Y(\i59/n534 ));
 NAND2xp5_ASAP7_75t_SL \i59/i542  (.A(\i59/n523 ),
    .B(\i59/n42 ),
    .Y(\i59/n535 ));
 AND2x2_ASAP7_75t_SL \i59/i543  (.A(n3[2]),
    .B(n3[0]),
    .Y(\i59/n536 ));
 AND2x2_ASAP7_75t_SL \i59/i544  (.A(n3[1]),
    .B(\i59/n19 ),
    .Y(\i59/n537 ));
 NAND2xp5_ASAP7_75t_SL \i59/i545  (.A(\i59/n538 ),
    .B(\i59/n523 ),
    .Y(\i59/n539 ));
 AND2x2_ASAP7_75t_SL \i59/i546  (.A(\i59/n536 ),
    .B(\i59/n537 ),
    .Y(\i59/n538 ));
 AOI22xp5_ASAP7_75t_SL \i59/i547  (.A1(\i59/n538 ),
    .A2(\i59/n511 ),
    .B1(\i59/n50 ),
    .B2(\i59/n77 ),
    .Y(\i59/n540 ));
 O2A1O1Ixp33_ASAP7_75t_SL \i59/i548  (.A1(\i59/n538 ),
    .A2(\i59/n507 ),
    .B(\i59/n1 ),
    .C(\i59/n71 ),
    .Y(\i59/n541 ));
 AOI221x1_ASAP7_75t_SL \i59/i549  (.A1(\i59/n1 ),
    .A2(\i59/n57 ),
    .B1(\i59/n538 ),
    .B2(\i59/n168 ),
    .C(\i59/n159 ),
    .Y(\i59/n542 ));
 NAND2xp33_ASAP7_75t_SL \i59/i55  (.A(\i59/n407 ),
    .B(\i59/n489 ),
    .Y(\i59/n439 ));
 NAND2xp5_ASAP7_75t_SL \i59/i550  (.A(\i59/n79 ),
    .B(\i59/n538 ),
    .Y(\i59/n543 ));
 NOR2xp33_ASAP7_75t_SL \i59/i551  (.A(\i59/n538 ),
    .B(\i59/n69 ),
    .Y(\i59/n544 ));
 AOI22xp5_ASAP7_75t_SL \i59/i552  (.A1(\i59/n538 ),
    .A2(\i59/n61 ),
    .B1(\i59/n75 ),
    .B2(\i59/n77 ),
    .Y(\i59/n545 ));
 NAND2xp5_ASAP7_75t_SL \i59/i553  (.A(\i59/n75 ),
    .B(\i59/n538 ),
    .Y(\i59/n546 ));
 NAND2xp5_ASAP7_75t_SL \i59/i554  (.A(\i59/n538 ),
    .B(\i59/n53 ),
    .Y(\i59/n547 ));
 AND2x2_ASAP7_75t_SL \i59/i555  (.A(\i59/n85 ),
    .B(\i59/n538 ),
    .Y(\i59/n548 ));
 AOI222xp33_ASAP7_75t_SL \i59/i556  (.A1(\i59/n57 ),
    .A2(\i59/n53 ),
    .B1(\i59/n538 ),
    .B2(\i59/n73 ),
    .C1(\i59/n62 ),
    .C2(\i59/n79 ),
    .Y(\i59/n349 ));
 NOR2xp33_ASAP7_75t_SL \i59/i557  (.A(\i59/n538 ),
    .B(\i59/n71 ),
    .Y(\i59/n549 ));
 OAI21xp5_ASAP7_75t_SL \i59/i558  (.A1(\i59/n538 ),
    .A2(\i59/n67 ),
    .B(\i59/n1 ),
    .Y(\i59/n550 ));
 AND4x1_ASAP7_75t_SL \i59/i559  (.A(\i59/n423 ),
    .B(\i59/n188 ),
    .C(\i59/n14 ),
    .D(\i59/n416 ),
    .Y(\i59/n551 ));
 NOR2xp33_ASAP7_75t_SL \i59/i56  (.A(\i59/n386 ),
    .B(\i59/n403 ),
    .Y(\i59/n438 ));
 NOR4xp25_ASAP7_75t_SL \i59/i560  (.A(\i59/n555 ),
    .B(\i59/n306 ),
    .C(\i59/n127 ),
    .D(\i59/n233 ),
    .Y(\i59/n552 ));
 AND4x1_ASAP7_75t_SL \i59/i561  (.A(\i59/n198 ),
    .B(\i59/n543 ),
    .C(\i59/n145 ),
    .D(\i59/n11 ),
    .Y(\i59/n553 ));
 NOR2x1p5_ASAP7_75t_SL \i59/i562  (.A(\i59/n3 ),
    .B(n3[6]),
    .Y(\i59/n554 ));
 NAND4xp25_ASAP7_75t_SL \i59/i563  (.A(\i59/n10 ),
    .B(\i59/n146 ),
    .C(\i59/n203 ),
    .D(\i59/n346 ),
    .Y(\i59/n555 ));
 NAND5xp2_ASAP7_75t_SL \i59/i57  (.A(\i59/n343 ),
    .B(\i59/n301 ),
    .C(\i59/n293 ),
    .D(\i59/n312 ),
    .E(\i59/n322 ),
    .Y(\i59/n437 ));
 NOR3xp33_ASAP7_75t_SL \i59/i58  (.A(\i59/n358 ),
    .B(\i59/n268 ),
    .C(\i59/n329 ),
    .Y(\i59/n436 ));
 NAND2xp33_ASAP7_75t_SL \i59/i59  (.A(\i59/n385 ),
    .B(\i59/n407 ),
    .Y(\i59/n435 ));
 AND5x2_ASAP7_75t_SL \i59/i6  (.A(\i59/n464 ),
    .B(\i59/n443 ),
    .C(\i59/n433 ),
    .D(\i59/n465 ),
    .E(\i59/n463 ),
    .Y(n2[1]));
 NAND4xp25_ASAP7_75t_SL \i59/i60  (.A(\i59/n395 ),
    .B(\i59/n372 ),
    .C(\i59/n298 ),
    .D(\i59/n317 ),
    .Y(\i59/n434 ));
 NOR3xp33_ASAP7_75t_SL \i59/i61  (.A(\i59/n406 ),
    .B(\i59/n369 ),
    .C(\i59/n390 ),
    .Y(\i59/n433 ));
 NAND5xp2_ASAP7_75t_SL \i59/i62  (.A(\i59/n376 ),
    .B(\i59/n344 ),
    .C(\i59/n339 ),
    .D(\i59/n220 ),
    .E(\i59/n305 ),
    .Y(\i59/n432 ));
 NOR4xp25_ASAP7_75t_SL \i59/i63  (.A(\i59/n363 ),
    .B(\i59/n364 ),
    .C(\i59/n222 ),
    .D(\i59/n192 ),
    .Y(\i59/n431 ));
 NAND2xp33_ASAP7_75t_SL \i59/i64  (.A(\i59/n411 ),
    .B(\i59/n389 ),
    .Y(\i59/n430 ));
 NOR3x1_ASAP7_75t_SL \i59/i65  (.A(\i59/n492 ),
    .B(\i59/n342 ),
    .C(\i59/n381 ),
    .Y(\i59/n443 ));
 INVxp67_ASAP7_75t_SL \i59/i66  (.A(\i59/n428 ),
    .Y(\i59/n429 ));
 INVx1_ASAP7_75t_SL \i59/i67  (.A(\i59/n424 ),
    .Y(\i59/n425 ));
 INVxp67_ASAP7_75t_SL \i59/i68  (.A(\i59/n422 ),
    .Y(\i59/n423 ));
 INVxp67_ASAP7_75t_SL \i59/i69  (.A(\i59/n420 ),
    .Y(\i59/n421 ));
 NOR2xp33_ASAP7_75t_SL \i59/i7  (.A(\i59/n455 ),
    .B(\i59/n483 ),
    .Y(\i59/n484 ));
 NOR3xp33_ASAP7_75t_SL \i59/i70  (.A(\i59/n384 ),
    .B(\i59/n13 ),
    .C(\i59/n235 ),
    .Y(\i59/n419 ));
 NAND3xp33_ASAP7_75t_SL \i59/i71  (.A(\i59/n266 ),
    .B(\i59/n524 ),
    .C(\i59/n286 ),
    .Y(\i59/n418 ));
 NAND2xp5_ASAP7_75t_SL \i59/i72  (.A(\i59/n373 ),
    .B(\i59/n387 ),
    .Y(\i59/n417 ));
 NOR2xp33_ASAP7_75t_SL \i59/i73  (.A(\i59/n396 ),
    .B(\i59/n365 ),
    .Y(\i59/n416 ));
 NOR2xp33_ASAP7_75t_SL \i59/i74  (.A(\i59/n356 ),
    .B(\i59/n297 ),
    .Y(\i59/n415 ));
 NOR5xp2_ASAP7_75t_SL \i59/i75  (.A(\i59/n288 ),
    .B(\i59/n530 ),
    .C(\i59/n222 ),
    .D(\i59/n262 ),
    .E(\i59/n259 ),
    .Y(\i59/n414 ));
 NOR2xp33_ASAP7_75t_SL \i59/i76  (.A(\i59/n341 ),
    .B(\i59/n367 ),
    .Y(\i59/n413 ));
 AOI211xp5_ASAP7_75t_SL \i59/i77  (.A1(\i59/n328 ),
    .A2(\i59/n108 ),
    .B(\i59/n279 ),
    .C(\i59/n236 ),
    .Y(\i59/n412 ));
 NAND2xp5_ASAP7_75t_SL \i59/i78  (.A(\i59/n292 ),
    .B(\i59/n388 ),
    .Y(\i59/n428 ));
 NAND3xp33_ASAP7_75t_SL \i59/i79  (.A(\i59/n370 ),
    .B(\i59/n349 ),
    .C(\i59/n320 ),
    .Y(\i59/n427 ));
 AND4x2_ASAP7_75t_SL \i59/i8  (.A(\i59/n473 ),
    .B(\i59/n481 ),
    .C(\i59/n480 ),
    .D(\i59/n431 ),
    .Y(n2[5]));
 NOR2x1_ASAP7_75t_SL \i59/i80  (.A(\i59/n378 ),
    .B(\i59/n300 ),
    .Y(\i59/n426 ));
 AND3x1_ASAP7_75t_SL \i59/i81  (.A(\i59/n508 ),
    .B(\i59/n302 ),
    .C(\i59/n280 ),
    .Y(\i59/n424 ));
 NAND3xp33_ASAP7_75t_SL \i59/i82  (.A(\i59/n298 ),
    .B(\i59/n540 ),
    .C(\i59/n553 ),
    .Y(\i59/n422 ));
 NOR3x1_ASAP7_75t_SL \i59/i83  (.A(\i59/n299 ),
    .B(\i59/n324 ),
    .C(\i59/n231 ),
    .Y(\i59/n420 ));
 INVxp33_ASAP7_75t_SL \i59/i84  (.A(\i59/n408 ),
    .Y(\i59/n409 ));
 OAI211xp5_ASAP7_75t_SL \i59/i85  (.A1(\i59/n486 ),
    .A2(\i59/n182 ),
    .B(\i59/n316 ),
    .C(\i59/n251 ),
    .Y(\i59/n405 ));
 AOI211xp5_ASAP7_75t_SL \i59/i86  (.A1(\i59/n183 ),
    .A2(\i59/n47 ),
    .B(\i59/n277 ),
    .C(\i59/n490 ),
    .Y(\i59/n404 ));
 NAND4xp25_ASAP7_75t_SL \i59/i87  (.A(\i59/n289 ),
    .B(\i59/n325 ),
    .C(\i59/n291 ),
    .D(\i59/n512 ),
    .Y(\i59/n403 ));
 NAND4xp25_ASAP7_75t_SL \i59/i88  (.A(\i59/n349 ),
    .B(\i59/n250 ),
    .C(\i59/n311 ),
    .D(\i59/n207 ),
    .Y(\i59/n402 ));
 NOR3xp33_ASAP7_75t_SL \i59/i89  (.A(\i59/n315 ),
    .B(\i59/n269 ),
    .C(\i59/n272 ),
    .Y(\i59/n401 ));
 AND3x4_ASAP7_75t_SL \i59/i9  (.A(\i59/n475 ),
    .B(\i59/n479 ),
    .C(\i59/n445 ),
    .Y(n2[0]));
 NOR3xp33_ASAP7_75t_SL \i59/i90  (.A(\i59/n502 ),
    .B(\i59/n253 ),
    .C(\i59/n278 ),
    .Y(\i59/n411 ));
 NOR2xp67_ASAP7_75t_SL \i59/i91  (.A(\i59/n390 ),
    .B(\i59/n354 ),
    .Y(\i59/n400 ));
 NOR2xp33_ASAP7_75t_SL \i59/i92  (.A(\i59/n379 ),
    .B(\i59/n361 ),
    .Y(\i59/n399 ));
 NAND5xp2_ASAP7_75t_SL \i59/i93  (.A(\i59/n295 ),
    .B(\i59/n314 ),
    .C(\i59/n219 ),
    .D(\i59/n227 ),
    .E(\i59/n220 ),
    .Y(\i59/n410 ));
 NOR3xp33_ASAP7_75t_SL \i59/i94  (.A(\i59/n350 ),
    .B(\i59/n103 ),
    .C(\i59/n226 ),
    .Y(\i59/n408 ));
 NOR2xp33_ASAP7_75t_L \i59/i95  (.A(\i59/n352 ),
    .B(\i59/n335 ),
    .Y(\i59/n407 ));
 NOR2xp33_ASAP7_75t_SL \i59/i96  (.A(\i59/n342 ),
    .B(\i59/n492 ),
    .Y(\i59/n398 ));
 NAND2xp5_ASAP7_75t_SL \i59/i97  (.A(\i59/n360 ),
    .B(\i59/n393 ),
    .Y(\i59/n406 ));
 INVxp33_ASAP7_75t_SL \i59/i98  (.A(\i59/n395 ),
    .Y(\i59/n396 ));
 INVxp67_ASAP7_75t_SL \i59/i99  (.A(\i59/n391 ),
    .Y(\i59/n392 ));
 OAI22xp5_ASAP7_75t_SL i590 (.A1(n124),
    .A2(n490),
    .B1(n474),
    .B2(n491),
    .Y(n882));
 AOI22xp5_ASAP7_75t_SL i591 (.A1(n125),
    .A2(n545),
    .B1(n544),
    .B2(n475),
    .Y(n881));
 OAI22xp5_ASAP7_75t_SL i592 (.A1(n504),
    .A2(n476),
    .B1(n1163),
    .B2(n505),
    .Y(n880));
 OAI22xp5_ASAP7_75t_SL i593 (.A1(n1163),
    .A2(n814),
    .B1(n476),
    .B2(n815),
    .Y(n879));
 INVxp67_ASAP7_75t_SL i594 (.A(n877),
    .Y(n878));
 INVx1_ASAP7_75t_SL i595 (.A(n875),
    .Y(n876));
 INVx1_ASAP7_75t_SL i596 (.A(n221),
    .Y(n874));
 INVx1_ASAP7_75t_SL i597 (.A(n872),
    .Y(n873));
 INVx1_ASAP7_75t_SL i598 (.A(n870),
    .Y(n871));
 INVx1_ASAP7_75t_SL i599 (.A(n868),
    .Y(n869));
 INVx2_ASAP7_75t_SL i6 (.A(n28[7]),
    .Y(n89));
 OR3x1_ASAP7_75t_SL i60 (.A(n1[2]),
    .B(n1[1]),
    .C(n1[3]),
    .Y(n1150));
 INVx1_ASAP7_75t_SL i600 (.A(n866),
    .Y(n867));
 INVx1_ASAP7_75t_SL i601 (.A(n864),
    .Y(n865));
 INVx1_ASAP7_75t_SL i602 (.A(n862),
    .Y(n863));
 INVx1_ASAP7_75t_SL i603 (.A(n860),
    .Y(n861));
 INVx1_ASAP7_75t_SL i604 (.A(n858),
    .Y(n859));
 INVx1_ASAP7_75t_SL i605 (.A(n855),
    .Y(n856));
 INVx1_ASAP7_75t_SL i606 (.A(n219),
    .Y(n854));
 INVx1_ASAP7_75t_SL i607 (.A(n852),
    .Y(n853));
 INVx1_ASAP7_75t_SL i608 (.A(n850),
    .Y(n851));
 INVx1_ASAP7_75t_SL i609 (.A(n848),
    .Y(n849));
 XOR2x1_ASAP7_75t_SL i61 (.A(n12[2]),
    .Y(n1151),
    .B(n2[2]));
 INVx1_ASAP7_75t_SL i610 (.A(n846),
    .Y(n847));
 INVx1_ASAP7_75t_SL i611 (.A(n844),
    .Y(n845));
 INVx1_ASAP7_75t_SL i612 (.A(n842),
    .Y(n843));
 INVx1_ASAP7_75t_SL i613 (.A(n839),
    .Y(n840));
 INVx1_ASAP7_75t_SL i614 (.A(n837),
    .Y(n838));
 INVx1_ASAP7_75t_SL i615 (.A(n224),
    .Y(n836));
 INVx1_ASAP7_75t_SL i616 (.A(n834),
    .Y(n835));
 INVx1_ASAP7_75t_SL i617 (.A(n832),
    .Y(n833));
 INVx1_ASAP7_75t_SL i618 (.A(n830),
    .Y(n831));
 INVx1_ASAP7_75t_SL i619 (.A(n828),
    .Y(n829));
 XOR2x1_ASAP7_75t_SL i62 (.A(n18[7]),
    .Y(n1153),
    .B(n16[7]));
 INVx1_ASAP7_75t_SL i620 (.A(n826),
    .Y(n827));
 INVx1_ASAP7_75t_SL i621 (.A(n824),
    .Y(n825));
 INVx1_ASAP7_75t_SL i622 (.A(n1174),
    .Y(n822));
 INVx1_ASAP7_75t_SL i623 (.A(n820),
    .Y(n821));
 INVx1_ASAP7_75t_SL i624 (.A(n816),
    .Y(n817));
 INVx2_ASAP7_75t_SL i625 (.A(n815),
    .Y(n814));
 INVx1_ASAP7_75t_SL i626 (.A(n812),
    .Y(n813));
 INVx2_ASAP7_75t_SL i627 (.A(n810),
    .Y(n809));
 INVx2_ASAP7_75t_SL i628 (.A(n808),
    .Y(n807));
 INVx2_ASAP7_75t_L i629 (.A(n806),
    .Y(n805));
 XOR2x1_ASAP7_75t_SL i63 (.A(n6[1]),
    .Y(n1152),
    .B(n16[1]));
 INVx2_ASAP7_75t_SL i630 (.A(n803),
    .Y(n802));
 INVx2_ASAP7_75t_L i631 (.A(n801),
    .Y(n800));
 INVx2_ASAP7_75t_SL i632 (.A(n799),
    .Y(n798));
 INVx1_ASAP7_75t_SL i633 (.A(n796),
    .Y(n797));
 INVx1_ASAP7_75t_SL i634 (.A(n1167),
    .Y(n795));
 INVx2_ASAP7_75t_SL i635 (.A(n794),
    .Y(n793));
 INVx2_ASAP7_75t_SL i636 (.A(n1175),
    .Y(n792));
 INVx2_ASAP7_75t_SL i637 (.A(n791),
    .Y(n790));
 INVx2_ASAP7_75t_SL i638 (.A(n1176),
    .Y(n789));
 INVx2_ASAP7_75t_SL i639 (.A(n788),
    .Y(n787));
 XOR2x1_ASAP7_75t_SL i64 (.A(n24[7]),
    .Y(n1155),
    .B(n14[7]));
 INVx2_ASAP7_75t_SL i640 (.A(n786),
    .Y(n785));
 INVx2_ASAP7_75t_SL i641 (.A(n784),
    .Y(n783));
 INVx2_ASAP7_75t_SL i642 (.A(n782),
    .Y(n781));
 INVx2_ASAP7_75t_SL i643 (.A(n779),
    .Y(n780));
 INVx2_ASAP7_75t_SL i644 (.A(n223),
    .Y(n778));
 INVx2_ASAP7_75t_SL i645 (.A(n1232),
    .Y(n777));
 INVx1_ASAP7_75t_SL i646 (.A(n773),
    .Y(n774));
 INVx1_ASAP7_75t_SL i647 (.A(n771),
    .Y(n772));
 INVx2_ASAP7_75t_SL i648 (.A(n1177),
    .Y(n769));
 INVx2_ASAP7_75t_SL i649 (.A(n768),
    .Y(n767));
 XOR2x1_ASAP7_75t_SL i65 (.A(n14[1]),
    .Y(n1154),
    .B(n4[1]));
 INVx2_ASAP7_75t_SL i650 (.A(n765),
    .Y(n764));
 INVx2_ASAP7_75t_SL i651 (.A(n763),
    .Y(n762));
 INVx2_ASAP7_75t_SL i652 (.A(n761),
    .Y(n760));
 INVx2_ASAP7_75t_SL i653 (.A(n759),
    .Y(n758));
 INVx2_ASAP7_75t_SL i654 (.A(n757),
    .Y(n756));
 AOI22xp5_ASAP7_75t_SL i655 (.A1(n38),
    .A2(n0[68]),
    .B1(net223),
    .B2(net129),
    .Y(n755));
 AOI22xp5_ASAP7_75t_SL i656 (.A1(n38),
    .A2(n0[98]),
    .B1(net256),
    .B2(net129),
    .Y(n754));
 AOI22xp5_ASAP7_75t_SL i657 (.A1(n38),
    .A2(n0[1]),
    .B1(net170),
    .B2(net129),
    .Y(n753));
 AOI22xp5_ASAP7_75t_SL i658 (.A1(n38),
    .A2(n0[121]),
    .B1(net155),
    .B2(net129),
    .Y(n752));
 AOI22xp5_ASAP7_75t_SL i659 (.A1(n38),
    .A2(n0[120]),
    .B1(net154),
    .B2(net129),
    .Y(n751));
 DFFHQNx1_ASAP7_75t_SL i66 (.CLK(clk),
    .D(n1027),
    .QN(n1[0]));
 AOI22xp5_ASAP7_75t_SL i660 (.A1(n38),
    .A2(n0[86]),
    .B1(net243),
    .B2(net129),
    .Y(n750));
 AOI22xp5_ASAP7_75t_SL i661 (.A1(n38),
    .A2(n0[23]),
    .B1(net174),
    .B2(net129),
    .Y(n749));
 AOI22xp5_ASAP7_75t_SL i662 (.A1(n38),
    .A2(n0[49]),
    .B1(net202),
    .B2(net129),
    .Y(n748));
 AOI22xp5_ASAP7_75t_SL i663 (.A1(n38),
    .A2(n0[109]),
    .B1(net141),
    .B2(net129),
    .Y(n747));
 AOI22xp5_ASAP7_75t_SL i664 (.A1(n38),
    .A2(n0[43]),
    .B1(net196),
    .B2(net129),
    .Y(n746));
 AOI22xp5_ASAP7_75t_SL i665 (.A1(n38),
    .A2(n0[115]),
    .B1(net148),
    .B2(net129),
    .Y(n745));
 AOI22xp5_ASAP7_75t_SL i666 (.A1(n38),
    .A2(n0[96]),
    .B1(net254),
    .B2(net129),
    .Y(n744));
 AOI22xp5_ASAP7_75t_SL i667 (.A1(n38),
    .A2(n0[19]),
    .B1(net169),
    .B2(net129),
    .Y(n743));
 AOI22xp5_ASAP7_75t_SL i668 (.A1(n38),
    .A2(n0[53]),
    .B1(net207),
    .B2(net129),
    .Y(n742));
 AOI22xp5_ASAP7_75t_SL i669 (.A1(n38),
    .A2(n0[114]),
    .B1(net147),
    .B2(net129),
    .Y(n741));
 DFFHQNx1_ASAP7_75t_SL i67 (.CLK(clk),
    .D(n1029),
    .QN(n1[1]));
 AOI22xp5_ASAP7_75t_SL i670 (.A1(n38),
    .A2(n0[80]),
    .B1(net237),
    .B2(net129),
    .Y(n740));
 AOI22xp5_ASAP7_75t_SL i671 (.A1(n38),
    .A2(n0[113]),
    .B1(net146),
    .B2(net129),
    .Y(n739));
 AOI22xp5_ASAP7_75t_SL i672 (.A1(n38),
    .A2(n0[79]),
    .B1(net235),
    .B2(net129),
    .Y(n738));
 AOI22xp5_ASAP7_75t_SL i673 (.A1(n38),
    .A2(n0[11]),
    .B1(net153),
    .B2(net129),
    .Y(n737));
 AOI22xp5_ASAP7_75t_SL i674 (.A1(n38),
    .A2(n0[110]),
    .B1(net143),
    .B2(net129),
    .Y(n736));
 AOI22xp5_ASAP7_75t_SL i675 (.A1(n38),
    .A2(n0[52]),
    .B1(net206),
    .B2(net129),
    .Y(n735));
 AOI22xp5_ASAP7_75t_SL i676 (.A1(n38),
    .A2(n0[126]),
    .B1(net160),
    .B2(net129),
    .Y(n734));
 AOI22xp5_ASAP7_75t_SL i677 (.A1(n38),
    .A2(n0[95]),
    .B1(net253),
    .B2(net129),
    .Y(n733));
 AOI22xp5_ASAP7_75t_SL i678 (.A1(n38),
    .A2(n0[51]),
    .B1(net205),
    .B2(net129),
    .Y(n732));
 AOI22xp5_ASAP7_75t_SL i679 (.A1(n38),
    .A2(n0[75]),
    .B1(net231),
    .B2(net129),
    .Y(n731));
 DFFHQNx1_ASAP7_75t_SL i68 (.CLK(clk),
    .D(n1028),
    .QN(n1[2]));
 AOI22xp5_ASAP7_75t_SL i680 (.A1(n38),
    .A2(n0[74]),
    .B1(net230),
    .B2(net129),
    .Y(n730));
 AOI22xp5_ASAP7_75t_SL i681 (.A1(n38),
    .A2(n0[125]),
    .B1(net159),
    .B2(net129),
    .Y(n729));
 AOI22xp5_ASAP7_75t_SL i682 (.A1(n38),
    .A2(n0[103]),
    .B1(net135),
    .B2(net129),
    .Y(n728));
 AOI22xp5_ASAP7_75t_SL i683 (.A1(n38),
    .A2(n0[0]),
    .B1(net131),
    .B2(net129),
    .Y(n727));
 AOI22xp5_ASAP7_75t_SL i684 (.A1(n38),
    .A2(n0[2]),
    .B1(net181),
    .B2(net129),
    .Y(n726));
 AOI22xp5_ASAP7_75t_SL i685 (.A1(n38),
    .A2(n0[3]),
    .B1(net192),
    .B2(net129),
    .Y(n725));
 AOI22xp5_ASAP7_75t_SL i686 (.A1(n38),
    .A2(n0[4]),
    .B1(net203),
    .B2(net129),
    .Y(n724));
 AOI22xp5_ASAP7_75t_SL i687 (.A1(n38),
    .A2(n0[5]),
    .B1(net214),
    .B2(net129),
    .Y(n723));
 AOI22xp5_ASAP7_75t_SL i688 (.A1(n38),
    .A2(n0[6]),
    .B1(net225),
    .B2(net129),
    .Y(n722));
 AOI22xp5_ASAP7_75t_SL i689 (.A1(n38),
    .A2(n0[7]),
    .B1(net236),
    .B2(net129),
    .Y(n721));
 DFFHQNx1_ASAP7_75t_SL i69 (.CLK(clk),
    .D(n1030),
    .QN(n1[3]));
 AOI22xp5_ASAP7_75t_SL i690 (.A1(n38),
    .A2(n0[8]),
    .B1(net247),
    .B2(net129),
    .Y(n720));
 AOI22xp5_ASAP7_75t_SL i691 (.A1(n38),
    .A2(n0[9]),
    .B1(net258),
    .B2(net129),
    .Y(n719));
 AOI22xp5_ASAP7_75t_SL i692 (.A1(n38),
    .A2(n0[10]),
    .B1(net142),
    .B2(net129),
    .Y(n718));
 AOI22xp5_ASAP7_75t_SL i693 (.A1(n38),
    .A2(n0[12]),
    .B1(net162),
    .B2(net129),
    .Y(n717));
 AOI22xp5_ASAP7_75t_SL i694 (.A1(n38),
    .A2(n0[13]),
    .B1(net163),
    .B2(net129),
    .Y(n716));
 AOI22xp5_ASAP7_75t_SL i695 (.A1(n38),
    .A2(n0[14]),
    .B1(net164),
    .B2(net129),
    .Y(n715));
 AOI22xp5_ASAP7_75t_SL i696 (.A1(n38),
    .A2(n0[15]),
    .B1(net165),
    .B2(net129),
    .Y(n714));
 AOI22xp5_ASAP7_75t_SL i697 (.A1(n38),
    .A2(n0[16]),
    .B1(net166),
    .B2(net129),
    .Y(n713));
 AOI22xp5_ASAP7_75t_SL i698 (.A1(n38),
    .A2(n0[17]),
    .B1(net167),
    .B2(net129),
    .Y(n712));
 AOI22xp5_ASAP7_75t_SL i699 (.A1(n38),
    .A2(n0[18]),
    .B1(net168),
    .B2(net129),
    .Y(n711));
 INVx2_ASAP7_75t_SL i7 (.A(n26[7]),
    .Y(n90));
 SDFHx4_ASAP7_75t_SL i70 (.CLK(clk),
    .D(n352),
    .QN(n33[0]),
    .SE(n1229),
    .SI(n1103));
 AOI22xp5_ASAP7_75t_SL i700 (.A1(n38),
    .A2(n0[20]),
    .B1(net171),
    .B2(net129),
    .Y(n710));
 AOI22xp5_ASAP7_75t_SL i701 (.A1(n38),
    .A2(n0[21]),
    .B1(net172),
    .B2(net129),
    .Y(n709));
 AOI22xp5_ASAP7_75t_SL i702 (.A1(n38),
    .A2(n0[22]),
    .B1(net173),
    .B2(net129),
    .Y(n708));
 AOI22xp5_ASAP7_75t_SL i703 (.A1(n38),
    .A2(n0[24]),
    .B1(net175),
    .B2(net129),
    .Y(n707));
 AOI22xp5_ASAP7_75t_SL i704 (.A1(n38),
    .A2(n0[25]),
    .B1(net176),
    .B2(net129),
    .Y(n706));
 AOI22xp5_ASAP7_75t_SL i705 (.A1(n38),
    .A2(n0[26]),
    .B1(net177),
    .B2(net129),
    .Y(n705));
 AOI22xp5_ASAP7_75t_SL i706 (.A1(n38),
    .A2(n0[27]),
    .B1(net178),
    .B2(net129),
    .Y(n704));
 AOI22xp5_ASAP7_75t_SL i707 (.A1(n38),
    .A2(n0[28]),
    .B1(net179),
    .B2(net129),
    .Y(n703));
 AOI22xp5_ASAP7_75t_SL i708 (.A1(n38),
    .A2(n0[29]),
    .B1(net180),
    .B2(net129),
    .Y(n702));
 AOI22xp5_ASAP7_75t_SL i709 (.A1(n38),
    .A2(n0[30]),
    .B1(net182),
    .B2(net129),
    .Y(n701));
 SDFHx4_ASAP7_75t_SL i71 (.CLK(clk),
    .D(n370),
    .QN(n33[1]),
    .SE(n1229),
    .SI(n1096));
 AOI22xp5_ASAP7_75t_SL i710 (.A1(n38),
    .A2(n0[31]),
    .B1(net183),
    .B2(net129),
    .Y(n700));
 AOI22xp5_ASAP7_75t_SL i711 (.A1(n38),
    .A2(n0[32]),
    .B1(net184),
    .B2(net129),
    .Y(n699));
 AOI22xp5_ASAP7_75t_SL i712 (.A1(n38),
    .A2(n0[33]),
    .B1(net185),
    .B2(net129),
    .Y(n698));
 AOI22xp5_ASAP7_75t_SL i713 (.A1(n38),
    .A2(n0[34]),
    .B1(net186),
    .B2(net129),
    .Y(n697));
 AOI22xp5_ASAP7_75t_SL i714 (.A1(n38),
    .A2(n0[35]),
    .B1(net187),
    .B2(net129),
    .Y(n696));
 AOI22xp5_ASAP7_75t_SL i715 (.A1(n38),
    .A2(n0[36]),
    .B1(net188),
    .B2(net129),
    .Y(n695));
 AOI22xp5_ASAP7_75t_SL i716 (.A1(n38),
    .A2(n0[37]),
    .B1(net189),
    .B2(net129),
    .Y(n694));
 AOI22xp5_ASAP7_75t_SL i717 (.A1(n38),
    .A2(n0[38]),
    .B1(net190),
    .B2(net129),
    .Y(n693));
 AOI22xp5_ASAP7_75t_SL i718 (.A1(n38),
    .A2(n0[39]),
    .B1(net191),
    .B2(net129),
    .Y(n692));
 AOI22xp5_ASAP7_75t_SL i719 (.A1(n38),
    .A2(n0[40]),
    .B1(net193),
    .B2(net129),
    .Y(n691));
 SDFHx4_ASAP7_75t_SL i72 (.CLK(clk),
    .D(n378),
    .QN(n33[2]),
    .SE(n1229),
    .SI(n1143));
 AOI22xp5_ASAP7_75t_SL i720 (.A1(n38),
    .A2(n0[41]),
    .B1(net194),
    .B2(net129),
    .Y(n690));
 AOI22xp5_ASAP7_75t_SL i721 (.A1(n38),
    .A2(n0[42]),
    .B1(net195),
    .B2(net129),
    .Y(n689));
 AOI22xp5_ASAP7_75t_SL i722 (.A1(n38),
    .A2(n0[44]),
    .B1(net197),
    .B2(net129),
    .Y(n688));
 AOI22xp5_ASAP7_75t_SL i723 (.A1(n38),
    .A2(n0[45]),
    .B1(net198),
    .B2(net129),
    .Y(n687));
 AOI22xp5_ASAP7_75t_SL i724 (.A1(n38),
    .A2(n0[46]),
    .B1(net199),
    .B2(net129),
    .Y(n686));
 AOI22xp5_ASAP7_75t_SL i725 (.A1(n38),
    .A2(n0[47]),
    .B1(net200),
    .B2(net129),
    .Y(n685));
 AOI22xp5_ASAP7_75t_SL i726 (.A1(n38),
    .A2(n0[48]),
    .B1(net201),
    .B2(net129),
    .Y(n684));
 AOI22xp5_ASAP7_75t_SL i727 (.A1(n38),
    .A2(n0[50]),
    .B1(net204),
    .B2(net129),
    .Y(n683));
 AOI22xp5_ASAP7_75t_SL i728 (.A1(n38),
    .A2(n0[54]),
    .B1(net208),
    .B2(net129),
    .Y(n682));
 AOI22xp5_ASAP7_75t_SL i729 (.A1(n38),
    .A2(n0[55]),
    .B1(net209),
    .B2(net129),
    .Y(n681));
 SDFHx4_ASAP7_75t_SL i73 (.CLK(clk),
    .D(n386),
    .QN(n33[3]),
    .SE(n1229),
    .SI(n1092));
 AOI22xp5_ASAP7_75t_SL i730 (.A1(n38),
    .A2(n0[56]),
    .B1(net210),
    .B2(net129),
    .Y(n680));
 AOI22xp5_ASAP7_75t_SL i731 (.A1(n38),
    .A2(n0[57]),
    .B1(net211),
    .B2(net129),
    .Y(n679));
 AOI22xp5_ASAP7_75t_SL i732 (.A1(n38),
    .A2(n0[58]),
    .B1(net212),
    .B2(net129),
    .Y(n678));
 AOI22xp5_ASAP7_75t_SL i733 (.A1(n38),
    .A2(n0[59]),
    .B1(net213),
    .B2(net129),
    .Y(n677));
 AOI22xp5_ASAP7_75t_SL i734 (.A1(n38),
    .A2(n0[60]),
    .B1(net215),
    .B2(net129),
    .Y(n676));
 AOI22xp5_ASAP7_75t_SL i735 (.A1(n38),
    .A2(n0[61]),
    .B1(net216),
    .B2(net129),
    .Y(n675));
 AOI22xp5_ASAP7_75t_SL i736 (.A1(n38),
    .A2(n0[62]),
    .B1(net217),
    .B2(net129),
    .Y(n674));
 AOI22xp5_ASAP7_75t_SL i737 (.A1(n38),
    .A2(n0[63]),
    .B1(net218),
    .B2(net129),
    .Y(n673));
 AOI22xp5_ASAP7_75t_SL i738 (.A1(n38),
    .A2(n0[64]),
    .B1(net219),
    .B2(net129),
    .Y(n672));
 AOI22xp5_ASAP7_75t_SL i739 (.A1(n38),
    .A2(n0[65]),
    .B1(net220),
    .B2(net129),
    .Y(n671));
 SDFHx4_ASAP7_75t_SL i74 (.CLK(clk),
    .D(n395),
    .QN(n33[4]),
    .SE(n1229),
    .SI(n1088));
 AOI22xp5_ASAP7_75t_SL i740 (.A1(n38),
    .A2(n0[66]),
    .B1(net221),
    .B2(net129),
    .Y(n670));
 AOI22xp5_ASAP7_75t_SL i741 (.A1(n38),
    .A2(n0[67]),
    .B1(net222),
    .B2(net129),
    .Y(n669));
 AOI22xp5_ASAP7_75t_SL i742 (.A1(n38),
    .A2(n0[69]),
    .B1(net224),
    .B2(net129),
    .Y(n668));
 AOI22xp5_ASAP7_75t_SL i743 (.A1(n38),
    .A2(n0[70]),
    .B1(net226),
    .B2(net129),
    .Y(n667));
 AOI22xp5_ASAP7_75t_SL i744 (.A1(n38),
    .A2(n0[71]),
    .B1(net227),
    .B2(net129),
    .Y(n666));
 AOI22xp5_ASAP7_75t_SL i745 (.A1(n38),
    .A2(n0[72]),
    .B1(net228),
    .B2(net129),
    .Y(n665));
 AOI22xp5_ASAP7_75t_SL i746 (.A1(n38),
    .A2(n0[73]),
    .B1(net229),
    .B2(net129),
    .Y(n664));
 AOI22xp5_ASAP7_75t_SL i747 (.A1(n38),
    .A2(n0[76]),
    .B1(net232),
    .B2(net129),
    .Y(n663));
 AOI22xp5_ASAP7_75t_SL i748 (.A1(n38),
    .A2(n0[77]),
    .B1(net233),
    .B2(net129),
    .Y(n662));
 AOI22xp5_ASAP7_75t_SL i749 (.A1(n38),
    .A2(n0[78]),
    .B1(net234),
    .B2(net129),
    .Y(n661));
 SDFHx4_ASAP7_75t_SL i75 (.CLK(clk),
    .D(n406),
    .QN(n33[5]),
    .SE(n1229),
    .SI(n1081));
 AOI22xp5_ASAP7_75t_SL i750 (.A1(n38),
    .A2(n0[81]),
    .B1(net238),
    .B2(net129),
    .Y(n660));
 AOI22xp5_ASAP7_75t_SL i751 (.A1(n38),
    .A2(n0[82]),
    .B1(net239),
    .B2(net129),
    .Y(n659));
 AOI22xp5_ASAP7_75t_SL i752 (.A1(n38),
    .A2(n0[83]),
    .B1(net240),
    .B2(net129),
    .Y(n658));
 AOI22xp5_ASAP7_75t_SL i753 (.A1(n38),
    .A2(n0[84]),
    .B1(net241),
    .B2(net129),
    .Y(n657));
 AOI22xp5_ASAP7_75t_SL i754 (.A1(n38),
    .A2(n0[85]),
    .B1(net242),
    .B2(net129),
    .Y(n656));
 AOI22xp5_ASAP7_75t_SL i755 (.A1(n38),
    .A2(n0[87]),
    .B1(net244),
    .B2(net129),
    .Y(n655));
 AOI22xp5_ASAP7_75t_SL i756 (.A1(n38),
    .A2(n0[88]),
    .B1(net245),
    .B2(net129),
    .Y(n654));
 AOI22xp5_ASAP7_75t_SL i757 (.A1(n38),
    .A2(n0[89]),
    .B1(net246),
    .B2(net129),
    .Y(n653));
 AOI22xp5_ASAP7_75t_SL i758 (.A1(n38),
    .A2(n0[91]),
    .B1(net249),
    .B2(net129),
    .Y(n652));
 AOI22xp5_ASAP7_75t_SL i759 (.A1(n38),
    .A2(n0[92]),
    .B1(net250),
    .B2(net129),
    .Y(n651));
 SDFHx4_ASAP7_75t_SL i76 (.CLK(clk),
    .D(n415),
    .QN(n33[6]),
    .SE(n1229),
    .SI(n1076));
 AOI22xp5_ASAP7_75t_SL i760 (.A1(n38),
    .A2(n0[93]),
    .B1(net251),
    .B2(net129),
    .Y(n650));
 AOI22xp5_ASAP7_75t_SL i761 (.A1(n38),
    .A2(n0[94]),
    .B1(net252),
    .B2(net129),
    .Y(n649));
 AOI22xp5_ASAP7_75t_SL i762 (.A1(n38),
    .A2(n0[97]),
    .B1(net255),
    .B2(net129),
    .Y(n648));
 AOI22xp5_ASAP7_75t_SL i763 (.A1(n38),
    .A2(n0[101]),
    .B1(net133),
    .B2(net129),
    .Y(n647));
 AOI22xp5_ASAP7_75t_SL i764 (.A1(n38),
    .A2(n0[102]),
    .B1(net134),
    .B2(net129),
    .Y(n646));
 AOI22xp5_ASAP7_75t_SL i765 (.A1(n38),
    .A2(n0[104]),
    .B1(net136),
    .B2(net129),
    .Y(n645));
 AOI22xp5_ASAP7_75t_SL i766 (.A1(n38),
    .A2(n0[105]),
    .B1(net137),
    .B2(net129),
    .Y(n644));
 AOI22xp5_ASAP7_75t_SL i767 (.A1(n38),
    .A2(n0[106]),
    .B1(net138),
    .B2(net129),
    .Y(n643));
 AOI22xp5_ASAP7_75t_SL i768 (.A1(n38),
    .A2(n0[107]),
    .B1(net139),
    .B2(net129),
    .Y(n642));
 AOI22xp5_ASAP7_75t_SL i769 (.A1(n38),
    .A2(n0[108]),
    .B1(net140),
    .B2(net129),
    .Y(n641));
 SDFHx4_ASAP7_75t_SL i77 (.CLK(clk),
    .D(n422),
    .QN(n33[7]),
    .SE(n1229),
    .SI(n1068));
 AOI22xp5_ASAP7_75t_SL i770 (.A1(n38),
    .A2(n0[111]),
    .B1(net144),
    .B2(net129),
    .Y(n640));
 AOI22xp5_ASAP7_75t_SL i771 (.A1(n38),
    .A2(n0[112]),
    .B1(net145),
    .B2(net129),
    .Y(n639));
 AOI22xp5_ASAP7_75t_SL i772 (.A1(n38),
    .A2(n0[116]),
    .B1(net149),
    .B2(net129),
    .Y(n638));
 AOI22xp5_ASAP7_75t_SL i773 (.A1(n38),
    .A2(n0[117]),
    .B1(net150),
    .B2(net129),
    .Y(n637));
 AOI22xp5_ASAP7_75t_SL i774 (.A1(n38),
    .A2(n0[118]),
    .B1(net151),
    .B2(net129),
    .Y(n636));
 AOI22xp5_ASAP7_75t_SL i775 (.A1(n38),
    .A2(n0[119]),
    .B1(net152),
    .B2(net129),
    .Y(n635));
 AOI22xp5_ASAP7_75t_SL i776 (.A1(n38),
    .A2(n0[122]),
    .B1(net156),
    .B2(net129),
    .Y(n634));
 AOI22xp5_ASAP7_75t_SL i777 (.A1(n38),
    .A2(n0[123]),
    .B1(net157),
    .B2(net129),
    .Y(n633));
 AOI22xp5_ASAP7_75t_SL i778 (.A1(n38),
    .A2(n0[124]),
    .B1(net158),
    .B2(net129),
    .Y(n632));
 AOI22xp5_ASAP7_75t_SL i779 (.A1(n38),
    .A2(n0[127]),
    .B1(net161),
    .B2(net129),
    .Y(n631));
 SDFHx4_ASAP7_75t_SL i78 (.CLK(clk),
    .D(n451),
    .QN(n31[0]),
    .SE(n1229),
    .SI(n1066));
 AOI22xp5_ASAP7_75t_SL i780 (.A1(n38),
    .A2(n0[99]),
    .B1(net257),
    .B2(net129),
    .Y(n630));
 AOI22xp5_ASAP7_75t_SL i781 (.A1(n38),
    .A2(n0[100]),
    .B1(net132),
    .B2(net129),
    .Y(n629));
 AOI22xp5_ASAP7_75t_SL i782 (.A1(n38),
    .A2(n0[90]),
    .B1(net248),
    .B2(net129),
    .Y(n628));
 NOR2xp33_ASAP7_75t_SL i783 (.A(n1[2]),
    .B(n293),
    .Y(n877));
 AOI22xp5_ASAP7_75t_SL i784 (.A1(n35[16]),
    .A2(n146),
    .B1(n291),
    .B2(n28[0]),
    .Y(n875));
 OAI22xp33_ASAP7_75t_SL i785 (.A1(n239),
    .A2(n10[3]),
    .B1(n36[3]),
    .B2(n1158),
    .Y(n627));
 OAI22xp5_ASAP7_75t_SL i786 (.A1(n262),
    .A2(n6[4]),
    .B1(n35[28]),
    .B2(n115),
    .Y(n626));
 AOI22xp5_ASAP7_75t_SL i787 (.A1(n22[5]),
    .A2(n1221),
    .B1(n22[4]),
    .B2(n94),
    .Y(n625));
 OAI22xp5_ASAP7_75t_SL i788 (.A1(n245),
    .A2(n8[0]),
    .B1(n36[8]),
    .B2(n149),
    .Y(n872));
 OAI22xp5_ASAP7_75t_SL i789 (.A1(n43),
    .A2(n22[2]),
    .B1(n37[26]),
    .B2(n229),
    .Y(n870));
 SDFHx4_ASAP7_75t_SL i79 (.CLK(clk),
    .D(n424),
    .QN(n31[1]),
    .SE(n1229),
    .SI(n1059));
 OAI22xp5_ASAP7_75t_SL i790 (.A1(n150),
    .A2(n10[2]),
    .B1(n8[1]),
    .B2(n145),
    .Y(n868));
 OAI22xp5_ASAP7_75t_SL i791 (.A1(n139),
    .A2(n10[6]),
    .B1(n8[5]),
    .B2(n171),
    .Y(n624));
 XOR2xp5_ASAP7_75t_SL i792 (.A(n30[1]),
    .B(n36[2]),
    .Y(n623));
 OAI22xp5_ASAP7_75t_SL i793 (.A1(n282),
    .A2(n8[1]),
    .B1(n36[9]),
    .B2(n150),
    .Y(n866));
 OAI22xp5_ASAP7_75t_SL i794 (.A1(n249),
    .A2(n8[2]),
    .B1(n36[10]),
    .B2(n113),
    .Y(n864));
 AOI22xp5_ASAP7_75t_SL i795 (.A1(n37[29]),
    .A2(n197),
    .B1(n41),
    .B2(n32[4]),
    .Y(n622));
 OAI22xp5_ASAP7_75t_SL i796 (.A1(n16[6]),
    .A2(n1161),
    .B1(n185),
    .B2(n16[7]),
    .Y(n862));
 AOI22xp5_ASAP7_75t_SL i797 (.A1(n18[5]),
    .A2(n178),
    .B1(n144),
    .B2(n18[4]),
    .Y(n621));
 OAI22xp5_ASAP7_75t_SL i798 (.A1(n257),
    .A2(n8[3]),
    .B1(n36[11]),
    .B2(n112),
    .Y(n860));
 AOI22xp5_ASAP7_75t_SL i799 (.A1(n35[29]),
    .A2(n154),
    .B1(n290),
    .B2(n28[4]),
    .Y(n620));
 INVxp67_ASAP7_75t_SL i8 (.A(n26[6]),
    .Y(n91));
 SDFHx4_ASAP7_75t_SL i80 (.CLK(clk),
    .D(n367),
    .QN(n31[2]),
    .SE(n1229),
    .SI(n1054));
 OAI22xp5_ASAP7_75t_SL i800 (.A1(n266),
    .A2(n10[5]),
    .B1(n36[5]),
    .B2(n199),
    .Y(n619));
 OAI22xp5_ASAP7_75t_SL i801 (.A1(n283),
    .A2(n20[4]),
    .B1(n36[12]),
    .B2(n162),
    .Y(n858));
 AOI22xp33_ASAP7_75t_SL i802 (.A1(n8[0]),
    .A2(n88),
    .B1(n149),
    .B2(n30[0]),
    .Y(n618));
 AOI22xp5_ASAP7_75t_SL i803 (.A1(n36[1]),
    .A2(n109),
    .B1(n237),
    .B2(n10[1]),
    .Y(n617));
 OAI22xp5_ASAP7_75t_R i804 (.A1(n274),
    .A2(n10[4]),
    .B1(n36[13]),
    .B2(n196),
    .Y(n616));
 OAI22xp5_ASAP7_75t_SL i805 (.A1(n12[2]),
    .A2(n229),
    .B1(n22[2]),
    .B2(n153),
    .Y(n615));
 AOI22xp5_ASAP7_75t_SL i806 (.A1(n8[5]),
    .A2(n111),
    .B1(n139),
    .B2(n8[4]),
    .Y(n857));
 OAI22xp5_ASAP7_75t_SL i807 (.A1(n256),
    .A2(n18[6]),
    .B1(n35[30]),
    .B2(n193),
    .Y(n614));
 OAI22xp5_ASAP7_75t_SL i808 (.A1(n232),
    .A2(n8[6]),
    .B1(n36[14]),
    .B2(n134),
    .Y(n613));
 XOR2xp5_ASAP7_75t_SL i809 (.A(n26[7]),
    .B(n34[7]),
    .Y(n612));
 SDFHx4_ASAP7_75t_SL i81 (.CLK(clk),
    .D(n445),
    .QN(n31[3]),
    .SE(n1229),
    .SI(n1050));
 XOR2xp5_ASAP7_75t_SL i810 (.A(n24[1]),
    .B(n34[18]),
    .Y(n611));
 AOI22xp5_ASAP7_75t_SL i811 (.A1(n180),
    .A2(n36[0]),
    .B1(n10[0]),
    .B2(n278),
    .Y(n855));
 OAI22xp5_ASAP7_75t_SL i812 (.A1(n238),
    .A2(n32[7]),
    .B1(n37[7]),
    .B2(n84),
    .Y(n610));
 OAI22xp5_ASAP7_75t_SL i813 (.A1(n246),
    .A2(n6[0]),
    .B1(n35[8]),
    .B2(n169),
    .Y(n852));
 OAI22xp33_ASAP7_75t_SL i814 (.A1(n122),
    .A2(n32[6]),
    .B1(n85),
    .B2(n2[6]),
    .Y(n609));
 AOI22xp5_ASAP7_75t_SL i815 (.A1(n37[17]),
    .A2(n147),
    .B1(n258),
    .B2(n32[1]),
    .Y(n608));
 AOI22xp33_ASAP7_75t_SL i816 (.A1(n137),
    .A2(n22[0]),
    .B1(n12[0]),
    .B2(n1225),
    .Y(n607));
 OAI22xp5_ASAP7_75t_SL i817 (.A1(n265),
    .A2(n22[0]),
    .B1(n37[24]),
    .B2(n1225),
    .Y(n850));
 OAI22xp5_ASAP7_75t_SL i818 (.A1(n260),
    .A2(n6[2]),
    .B1(n35[10]),
    .B2(n148),
    .Y(n848));
 OAI22xp5_ASAP7_75t_SL i819 (.A1(n247),
    .A2(n6[3]),
    .B1(n35[11]),
    .B2(n116),
    .Y(n846));
 SDFHx4_ASAP7_75t_SL i82 (.CLK(clk),
    .D(n460),
    .QN(n31[4]),
    .SE(n1229),
    .SI(n1049));
 OAI22xp5_ASAP7_75t_SL i820 (.A1(n77),
    .A2(n26[5]),
    .B1(n34[6]),
    .B2(n140),
    .Y(n606));
 OAI22xp5_ASAP7_75t_SL i821 (.A1(n56),
    .A2(n24[6]),
    .B1(n34[30]),
    .B2(n92),
    .Y(n605));
 OAI22xp5_ASAP7_75t_SL i822 (.A1(n50),
    .A2(n32[5]),
    .B1(n37[6]),
    .B2(n157),
    .Y(n604));
 OAI22xp5_ASAP7_75t_SL i823 (.A1(n236),
    .A2(n18[4]),
    .B1(n35[12]),
    .B2(n178),
    .Y(n844));
 OAI22xp5_ASAP7_75t_SL i824 (.A1(n16[3]),
    .A2(n98),
    .B1(n16[4]),
    .B2(n99),
    .Y(n603));
 AOI22xp33_ASAP7_75t_SL i825 (.A1(n24[2]),
    .A2(n141),
    .B1(n14[2]),
    .B2(n160),
    .Y(n602));
 AOI22xp5_ASAP7_75t_SL i826 (.A1(n230),
    .A2(n34[25]),
    .B1(n61),
    .B2(n24[1]),
    .Y(n842));
 AOI22xp5_ASAP7_75t_SL i827 (.A1(n6[5]),
    .A2(n115),
    .B1(n170),
    .B2(n6[4]),
    .Y(n841));
 OAI22xp33_ASAP7_75t_SL i828 (.A1(n181),
    .A2(n12[6]),
    .B1(n104),
    .B2(n2[5]),
    .Y(n601));
 OAI22xp5_ASAP7_75t_SL i829 (.A1(n51),
    .A2(n12[5]),
    .B1(n37[5]),
    .B2(n105),
    .Y(n600));
 SDFHx4_ASAP7_75t_SL i83 (.CLK(clk),
    .D(n450),
    .QN(n31[5]),
    .SE(n1229),
    .SI(n1046));
 OAI22xp5_ASAP7_75t_SL i830 (.A1(n268),
    .A2(n32[0]),
    .B1(n37[16]),
    .B2(n1165),
    .Y(n839));
 OAI22xp5_ASAP7_75t_SL i831 (.A1(n271),
    .A2(n6[6]),
    .B1(n35[14]),
    .B2(n167),
    .Y(n599));
 AOI22xp5_ASAP7_75t_SL i832 (.A1(n37[4]),
    .A2(n197),
    .B1(n234),
    .B2(n32[4]),
    .Y(n598));
 OAI22xp5_ASAP7_75t_SL i833 (.A1(n60),
    .A2(n24[2]),
    .B1(n34[26]),
    .B2(n160),
    .Y(n837));
 OAI22xp5_ASAP7_75t_SL i834 (.A1(n42),
    .A2(n2[4]),
    .B1(n37[28]),
    .B2(n184),
    .Y(n597));
 OAI22xp5_ASAP7_75t_SL i835 (.A1(n123),
    .A2(n32[3]),
    .B1(n2[3]),
    .B2(n1162),
    .Y(n596));
 OAI22xp5_ASAP7_75t_SL i836 (.A1(n76),
    .A2(n4[0]),
    .B1(n34[8]),
    .B2(n138),
    .Y(n834));
 OAI22xp5_ASAP7_75t_SL i837 (.A1(n231),
    .A2(n12[3]),
    .B1(n37[3]),
    .B2(n107),
    .Y(n595));
 OAI22xp5_ASAP7_75t_R i838 (.A1(n255),
    .A2(n18[6]),
    .B1(n35[23]),
    .B2(n193),
    .Y(n594));
 AOI22xp5_ASAP7_75t_SL i839 (.A1(n143),
    .A2(n36[22]),
    .B1(n276),
    .B2(n20[5]),
    .Y(n593));
 SDFHx4_ASAP7_75t_SL i84 (.CLK(clk),
    .D(n468),
    .QN(n31[6]),
    .SE(n1229),
    .SI(n1045));
 OAI22xp5_ASAP7_75t_SL i840 (.A1(n192),
    .A2(n12[2]),
    .B1(n2[1]),
    .B2(n153),
    .Y(n832));
 XOR2xp5_ASAP7_75t_SL i841 (.A(n32[1]),
    .B(n37[2]),
    .Y(n592));
 AOI22xp5_ASAP7_75t_SL i842 (.A1(n1222),
    .A2(n34[27]),
    .B1(n24[3]),
    .B2(n59),
    .Y(n830));
 OAI22xp5_ASAP7_75t_SL i843 (.A1(n74),
    .A2(n4[2]),
    .B1(n34[10]),
    .B2(n183),
    .Y(n828));
 OAI22xp5_ASAP7_75t_SL i844 (.A1(n52),
    .A2(n20[6]),
    .B1(n36[30]),
    .B2(n96),
    .Y(n591));
 OAI22xp5_ASAP7_75t_SL i845 (.A1(n78),
    .A2(n14[5]),
    .B1(n34[5]),
    .B2(n190),
    .Y(n590));
 OAI22xp5_ASAP7_75t_SL i846 (.A1(n194),
    .A2(n32[0]),
    .B1(n2[0]),
    .B2(n1165),
    .Y(n589));
 OAI22xp5_ASAP7_75t_SL i847 (.A1(n73),
    .A2(n4[3]),
    .B1(n34[11]),
    .B2(n120),
    .Y(n826));
 AOI22xp33_ASAP7_75t_SL i848 (.A1(n4[3]),
    .A2(n1227),
    .B1(n120),
    .B2(n26[3]),
    .Y(n588));
 OAI22xp5_ASAP7_75t_SL i849 (.A1(n58),
    .A2(n4[4]),
    .B1(n34[28]),
    .B2(n119),
    .Y(n587));
 SDFHx4_ASAP7_75t_SL i85 (.CLK(clk),
    .D(n389),
    .QN(n31[7]),
    .SE(n1229),
    .SI(n1044));
 OAI22xp5_ASAP7_75t_SL i850 (.A1(n72),
    .A2(n24[4]),
    .B1(n34[12]),
    .B2(n158),
    .Y(n824));
 AOI22xp5_ASAP7_75t_SL i851 (.A1(n4[5]),
    .A2(n119),
    .B1(n155),
    .B2(n4[4]),
    .Y(n823));
 AOI22xp5_ASAP7_75t_SL i852 (.A1(n137),
    .A2(n37[0]),
    .B1(n12[0]),
    .B2(n284),
    .Y(n820));
 OAI22xp5_ASAP7_75t_SL i853 (.A1(n71),
    .A2(n4[6]),
    .B1(n34[14]),
    .B2(n118),
    .Y(n586));
 AOI22xp5_ASAP7_75t_SL i854 (.A1(n24[5]),
    .A2(n158),
    .B1(n195),
    .B2(n24[4]),
    .Y(n585));
 AOI22xp5_ASAP7_75t_SL i855 (.A1(n34[29]),
    .A2(n161),
    .B1(n57),
    .B2(n26[4]),
    .Y(n584));
 AND3x1_ASAP7_75t_SL i856 (.A(n1150),
    .B(n38),
    .C(net130),
    .Y(n819));
 AO22x1_ASAP7_75t_SL i857 (.A1(n4[5]),
    .A2(n190),
    .B1(n155),
    .B2(n14[5]),
    .Y(n818));
 AOI22x1_ASAP7_75t_SL i858 (.A1(n140),
    .A2(n24[5]),
    .B1(n195),
    .B2(n26[5]),
    .Y(n816));
 OAI22x1_ASAP7_75t_SL i859 (.A1(n111),
    .A2(n30[4]),
    .B1(n8[4]),
    .B2(n87),
    .Y(n815));
 SDFHx4_ASAP7_75t_SL i86 (.CLK(clk),
    .D(n456),
    .QN(n29[0]),
    .SE(n1229),
    .SI(n1115));
 AOI22x1_ASAP7_75t_SL i860 (.A1(n101),
    .A2(n24[4]),
    .B1(n158),
    .B2(n14[4]),
    .Y(n812));
 OAI22xp5_ASAP7_75t_SL i861 (.A1(n118),
    .A2(n14[6]),
    .B1(n4[6]),
    .B2(n100),
    .Y(n811));
 AOI22x1_ASAP7_75t_SL i862 (.A1(n131),
    .A2(n22[2]),
    .B1(n229),
    .B2(n32[2]),
    .Y(n810));
 OAI22x1_ASAP7_75t_SL i863 (.A1(n176),
    .A2(n32[1]),
    .B1(n147),
    .B2(n22[1]),
    .Y(n808));
 AOI22x1_ASAP7_75t_SL i864 (.A1(n163),
    .A2(n24[2]),
    .B1(n160),
    .B2(n26[2]),
    .Y(n806));
 OAI22xp5_ASAP7_75t_SL i865 (.A1(n26[6]),
    .A2(n92),
    .B1(n24[6]),
    .B2(n91),
    .Y(n804));
 OAI22x1_ASAP7_75t_SL i866 (.A1(n120),
    .A2(n14[3]),
    .B1(n102),
    .B2(n4[3]),
    .Y(n803));
 AOI22x1_ASAP7_75t_SL i867 (.A1(n198),
    .A2(n20[2]),
    .B1(n168),
    .B2(n30[2]),
    .Y(n801));
 XNOR2x1_ASAP7_75t_SL i868 (.B(n22[4]),
    .Y(n799),
    .A(n12[4]));
 AOI22x1_ASAP7_75t_SL i869 (.A1(n98),
    .A2(n18[4]),
    .B1(n178),
    .B2(n16[4]),
    .Y(n796));
 SDFHx4_ASAP7_75t_SL i87 (.CLK(clk),
    .D(n459),
    .QN(n29[1]),
    .SE(n1229),
    .SI(n1128));
 OAI22x1_ASAP7_75t_SL i870 (.A1(n183),
    .A2(n14[2]),
    .B1(n4[2]),
    .B2(n141),
    .Y(n794));
 OAI22x1_ASAP7_75t_SL i871 (.A1(n26[1]),
    .A2(n230),
    .B1(n24[1]),
    .B2(n174),
    .Y(n791));
 OAI22x1_ASAP7_75t_SL i872 (.A1(n30[1]),
    .A2(n142),
    .B1(n20[1]),
    .B2(n159),
    .Y(n788));
 OAI22x1_ASAP7_75t_SL i873 (.A1(n26[0]),
    .A2(n130),
    .B1(n24[0]),
    .B2(n136),
    .Y(n786));
 OAI22x1_ASAP7_75t_SL i874 (.A1(n14[0]),
    .A2(n138),
    .B1(n4[0]),
    .B2(n132),
    .Y(n784));
 OAI22x1_ASAP7_75t_SL i875 (.A1(n194),
    .A2(n12[0]),
    .B1(n2[0]),
    .B2(n137),
    .Y(n782));
 OAI22x1_ASAP7_75t_SL i876 (.A1(n123),
    .A2(n12[3]),
    .B1(n107),
    .B2(n2[3]),
    .Y(n779));
 OAI22xp5_ASAP7_75t_SL i877 (.A1(n28[6]),
    .A2(n193),
    .B1(n18[6]),
    .B2(n1220),
    .Y(n776));
 OAI22xp5_ASAP7_75t_SL i878 (.A1(n167),
    .A2(n16[6]),
    .B1(n6[6]),
    .B2(n185),
    .Y(n775));
 AOI22x1_ASAP7_75t_SL i879 (.A1(n188),
    .A2(n18[5]),
    .B1(n144),
    .B2(n28[5]),
    .Y(n773));
 SDFHx4_ASAP7_75t_SL i88 (.CLK(clk),
    .D(n464),
    .QN(n29[2]),
    .SE(n1229),
    .SI(n225));
 AOI22xp5_ASAP7_75t_SL i880 (.A1(n105),
    .A2(n2[5]),
    .B1(n12[5]),
    .B2(n181),
    .Y(n771));
 OAI22xp5_ASAP7_75t_SL i881 (.A1(n30[6]),
    .A2(n96),
    .B1(n135),
    .B2(n20[6]),
    .Y(n770));
 OAI22x1_ASAP7_75t_SL i882 (.A1(n115),
    .A2(n28[4]),
    .B1(n154),
    .B2(n6[4]),
    .Y(n768));
 AO22x1_ASAP7_75t_SL i883 (.A1(n6[5]),
    .A2(n200),
    .B1(n170),
    .B2(n16[5]),
    .Y(n766));
 OAI22x1_ASAP7_75t_SL i884 (.A1(n114),
    .A2(n16[7]),
    .B1(n6[7]),
    .B2(n1161),
    .Y(n765));
 OAI22x1_ASAP7_75t_SL i885 (.A1(n110),
    .A2(n10[7]),
    .B1(n108),
    .B2(n8[7]),
    .Y(n763));
 OA22x2_ASAP7_75t_SL i886 (.A1(n32[7]),
    .A2(n93),
    .B1(n22[7]),
    .B2(n84),
    .Y(n761));
 OA22x2_ASAP7_75t_SL i887 (.A1(n1156),
    .A2(n26[7]),
    .B1(n90),
    .B2(n24[7]),
    .Y(n759));
 OAI22x1_ASAP7_75t_SL i888 (.A1(n117),
    .A2(n14[7]),
    .B1(n4[7]),
    .B2(n1157),
    .Y(n757));
 INVx1_ASAP7_75t_SL i889 (.A(n582),
    .Y(n583));
 SDFHx4_ASAP7_75t_SL i89 (.CLK(clk),
    .D(n469),
    .QN(n29[3]),
    .SE(n1229),
    .SI(n1038));
 INVx1_ASAP7_75t_SL i890 (.A(n1231),
    .Y(n581));
 INVx1_ASAP7_75t_SL i891 (.A(n579),
    .Y(n580));
 INVx1_ASAP7_75t_SL i892 (.A(n1230),
    .Y(n577));
 INVx1_ASAP7_75t_SL i893 (.A(n575),
    .Y(n576));
 INVx1_ASAP7_75t_SL i894 (.A(n573),
    .Y(n574));
 INVx1_ASAP7_75t_SL i895 (.A(n571),
    .Y(n572));
 INVx1_ASAP7_75t_SL i896 (.A(n569),
    .Y(n570));
 INVx1_ASAP7_75t_SL i897 (.A(n567),
    .Y(n568));
 INVx1_ASAP7_75t_SL i898 (.A(n565),
    .Y(n566));
 INVx1_ASAP7_75t_SL i899 (.A(n563),
    .Y(n564));
 INVx2_ASAP7_75t_SL i9 (.A(n24[6]),
    .Y(n92));
 SDFHx4_ASAP7_75t_SL i90 (.CLK(clk),
    .D(n363),
    .QN(n29[4]),
    .SE(n1229),
    .SI(n1113));
 INVx1_ASAP7_75t_SL i900 (.A(n561),
    .Y(n562));
 INVx1_ASAP7_75t_SL i901 (.A(n559),
    .Y(n560));
 INVx1_ASAP7_75t_SL i902 (.A(n557),
    .Y(n558));
 INVx1_ASAP7_75t_SL i903 (.A(n555),
    .Y(n556));
 INVx1_ASAP7_75t_SL i904 (.A(n553),
    .Y(n554));
 INVx1_ASAP7_75t_SL i905 (.A(n551),
    .Y(n552));
 INVx1_ASAP7_75t_SL i906 (.A(n218),
    .Y(n550));
 INVx1_ASAP7_75t_SL i907 (.A(n548),
    .Y(n549));
 INVx1_ASAP7_75t_SL i908 (.A(n546),
    .Y(n547));
 INVx1_ASAP7_75t_SL i909 (.A(n544),
    .Y(n545));
 SDFHx4_ASAP7_75t_SL i91 (.CLK(clk),
    .D(n360),
    .QN(n29[5]),
    .SE(n1229),
    .SI(n1110));
 INVx1_ASAP7_75t_SL i910 (.A(n1180),
    .Y(n543));
 INVx1_ASAP7_75t_SL i911 (.A(n541),
    .Y(n542));
 INVx1_ASAP7_75t_SL i912 (.A(n539),
    .Y(n540));
 INVx1_ASAP7_75t_SL i913 (.A(n537),
    .Y(n538));
 INVx1_ASAP7_75t_SL i914 (.A(n535),
    .Y(n536));
 INVx1_ASAP7_75t_SL i915 (.A(n1181),
    .Y(n534));
 INVx1_ASAP7_75t_SL i916 (.A(n217),
    .Y(n533));
 INVx1_ASAP7_75t_SL i917 (.A(n531),
    .Y(n532));
 INVx1_ASAP7_75t_SL i918 (.A(n529),
    .Y(n530));
 INVx1_ASAP7_75t_SL i919 (.A(n527),
    .Y(n528));
 SDFHx4_ASAP7_75t_SL i92 (.CLK(clk),
    .D(n356),
    .QN(n29[6]),
    .SE(n1229),
    .SI(n1107));
 INVx1_ASAP7_75t_SL i920 (.A(n525),
    .Y(n526));
 INVx1_ASAP7_75t_SL i921 (.A(n523),
    .Y(n524));
 INVx1_ASAP7_75t_SL i922 (.A(n521),
    .Y(n522));
 INVx1_ASAP7_75t_SL i923 (.A(n519),
    .Y(n520));
 INVx1_ASAP7_75t_SL i924 (.A(n517),
    .Y(n518));
 INVxp67_ASAP7_75t_SL i925 (.A(n515),
    .Y(n516));
 INVx1_ASAP7_75t_SL i926 (.A(n513),
    .Y(n514));
 INVx2_ASAP7_75t_L i927 (.A(n511),
    .Y(n510));
 INVx2_ASAP7_75t_SL i928 (.A(n509),
    .Y(n508));
 INVx2_ASAP7_75t_SL i929 (.A(n507),
    .Y(n506));
 SDFHx4_ASAP7_75t_SL i93 (.CLK(clk),
    .D(n351),
    .QN(n29[7]),
    .SE(n1229),
    .SI(n1125));
 INVx2_ASAP7_75t_SL i930 (.A(n504),
    .Y(n505));
 INVx1_ASAP7_75t_SL i931 (.A(n1210),
    .Y(n502));
 INVx2_ASAP7_75t_SL i932 (.A(n500),
    .Y(n499));
 INVx2_ASAP7_75t_SL i933 (.A(n498),
    .Y(n497));
 INVx1_ASAP7_75t_SL i934 (.A(n495),
    .Y(n496));
 INVx2_ASAP7_75t_SL i935 (.A(n493),
    .Y(n492));
 INVx2_ASAP7_75t_SL i936 (.A(n491),
    .Y(n490));
 INVx2_ASAP7_75t_SL i937 (.A(n489),
    .Y(n488));
 INVx2_ASAP7_75t_SL i938 (.A(n487),
    .Y(n486));
 INVx1_ASAP7_75t_SL i939 (.A(n484),
    .Y(n485));
 SDFHx4_ASAP7_75t_SL i94 (.CLK(clk),
    .D(n473),
    .QN(n27[0]),
    .SE(n1229),
    .SI(n1117));
 INVx2_ASAP7_75t_SL i940 (.A(n483),
    .Y(n482));
 INVx2_ASAP7_75t_SL i941 (.A(n481),
    .Y(n480));
 INVx2_ASAP7_75t_SL i942 (.A(n1211),
    .Y(n479));
 INVx2_ASAP7_75t_SL i943 (.A(n478),
    .Y(n477));
 XNOR2xp5_ASAP7_75t_SL i944 (.A(n0[24]),
    .B(n34[24]),
    .Y(n473));
 XNOR2xp5_ASAP7_75t_SL i945 (.A(n0[110]),
    .B(n37[14]),
    .Y(n472));
 XNOR2xp5_ASAP7_75t_SL i946 (.A(n0[118]),
    .B(n37[22]),
    .Y(n471));
 XNOR2xp5_ASAP7_75t_SL i947 (.A(n0[109]),
    .B(n37[13]),
    .Y(n470));
 XNOR2xp5_ASAP7_75t_SL i948 (.A(n0[59]),
    .B(n35[27]),
    .Y(n469));
 XNOR2xp5_ASAP7_75t_SL i949 (.A(n0[94]),
    .B(n36[30]),
    .Y(n468));
 SDFHx4_ASAP7_75t_SL i95 (.CLK(clk),
    .D(n369),
    .QN(n27[1]),
    .SE(n1229),
    .SI(n1146));
 XNOR2xp5_ASAP7_75t_SL i950 (.A(n0[108]),
    .B(n37[12]),
    .Y(n467));
 XNOR2xp5_ASAP7_75t_SL i951 (.A(n0[107]),
    .B(n37[11]),
    .Y(n466));
 XNOR2xp5_ASAP7_75t_SL i952 (.A(n0[81]),
    .B(n36[17]),
    .Y(n465));
 XNOR2xp5_ASAP7_75t_SL i953 (.A(n0[58]),
    .B(n35[26]),
    .Y(n464));
 XNOR2xp5_ASAP7_75t_SL i954 (.A(n0[106]),
    .B(n37[10]),
    .Y(n463));
 XNOR2xp5_ASAP7_75t_SL i955 (.A(n0[105]),
    .B(n37[9]),
    .Y(n462));
 XNOR2xp5_ASAP7_75t_SL i956 (.A(n0[104]),
    .B(n37[8]),
    .Y(n461));
 XNOR2xp5_ASAP7_75t_SL i957 (.A(n0[92]),
    .B(n36[28]),
    .Y(n460));
 XNOR2xp5_ASAP7_75t_SL i958 (.A(n0[57]),
    .B(n35[25]),
    .Y(n459));
 XNOR2xp5_ASAP7_75t_SL i959 (.A(n34[23]),
    .B(n0[23]),
    .Y(n458));
 SDFHx4_ASAP7_75t_SL i96 (.CLK(clk),
    .D(n373),
    .QN(n27[2]),
    .SE(n1229),
    .SI(n1119));
 XNOR2xp5_ASAP7_75t_SL i960 (.A(n34[22]),
    .B(n0[22]),
    .Y(n457));
 XNOR2xp5_ASAP7_75t_SL i961 (.A(n0[56]),
    .B(n35[24]),
    .Y(n456));
 XNOR2xp5_ASAP7_75t_SL i962 (.A(n34[21]),
    .B(n0[21]),
    .Y(n455));
 XNOR2xp5_ASAP7_75t_SL i963 (.A(n34[20]),
    .B(n0[20]),
    .Y(n454));
 XNOR2xp5_ASAP7_75t_SL i964 (.A(n34[16]),
    .B(n0[16]),
    .Y(n453));
 XNOR2xp5_ASAP7_75t_SL i965 (.A(n0[34]),
    .B(n35[2]),
    .Y(n452));
 XNOR2xp5_ASAP7_75t_SL i966 (.A(n0[88]),
    .B(n36[24]),
    .Y(n451));
 XNOR2xp5_ASAP7_75t_SL i967 (.A(n0[93]),
    .B(n36[29]),
    .Y(n450));
 XNOR2xp5_ASAP7_75t_SL i968 (.A(n0[53]),
    .B(n35[21]),
    .Y(n449));
 XNOR2xp5_ASAP7_75t_SL i969 (.A(n0[52]),
    .B(n35[20]),
    .Y(n448));
 SDFHx4_ASAP7_75t_SL i97 (.CLK(clk),
    .D(n377),
    .QN(n27[3]),
    .SE(n1229),
    .SI(n1098));
 XNOR2xp5_ASAP7_75t_SL i970 (.A(n0[50]),
    .B(n35[18]),
    .Y(n447));
 XNOR2xp5_ASAP7_75t_SL i971 (.A(n0[48]),
    .B(n35[16]),
    .Y(n446));
 XNOR2xp5_ASAP7_75t_SL i972 (.A(n0[91]),
    .B(n36[27]),
    .Y(n445));
 XNOR2xp5_ASAP7_75t_SL i973 (.A(n0[87]),
    .B(n36[23]),
    .Y(n444));
 XNOR2xp5_ASAP7_75t_SL i974 (.A(n0[54]),
    .B(n35[22]),
    .Y(n443));
 XNOR2xp5_ASAP7_75t_SL i975 (.A(n34[7]),
    .B(n0[7]),
    .Y(n442));
 XNOR2xp5_ASAP7_75t_SL i976 (.A(n34[6]),
    .B(n0[6]),
    .Y(n441));
 XNOR2xp5_ASAP7_75t_SL i977 (.A(n34[5]),
    .B(n0[5]),
    .Y(n440));
 XNOR2xp5_ASAP7_75t_SL i978 (.A(n34[18]),
    .B(n0[18]),
    .Y(n439));
 XNOR2xp5_ASAP7_75t_SL i979 (.A(n0[84]),
    .B(n36[20]),
    .Y(n438));
 SDFHx4_ASAP7_75t_SL i98 (.CLK(clk),
    .D(n383),
    .QN(n27[4]),
    .SE(n1229),
    .SI(n1094));
 XNOR2xp5_ASAP7_75t_SL i980 (.A(n34[2]),
    .B(n0[2]),
    .Y(n437));
 XNOR2xp5_ASAP7_75t_SL i981 (.A(n0[83]),
    .B(n36[19]),
    .Y(n436));
 XNOR2xp5_ASAP7_75t_SL i982 (.A(n0[0]),
    .B(n34[0]),
    .Y(n435));
 XNOR2xp5_ASAP7_75t_SL i983 (.A(n0[33]),
    .B(n35[1]),
    .Y(n434));
 XNOR2xp5_ASAP7_75t_SL i984 (.A(n34[1]),
    .B(n0[1]),
    .Y(n433));
 XNOR2xp5_ASAP7_75t_SL i985 (.A(n0[39]),
    .B(n35[7]),
    .Y(n432));
 XNOR2xp5_ASAP7_75t_SL i986 (.A(n0[82]),
    .B(n36[18]),
    .Y(n431));
 XNOR2xp5_ASAP7_75t_SL i987 (.A(n0[51]),
    .B(n35[19]),
    .Y(n430));
 XNOR2xp5_ASAP7_75t_SL i988 (.A(n0[38]),
    .B(n35[6]),
    .Y(n429));
 XNOR2xp5_ASAP7_75t_SL i989 (.A(n0[37]),
    .B(n35[5]),
    .Y(n428));
 SDFHx4_ASAP7_75t_SL i99 (.CLK(clk),
    .D(n387),
    .QN(n27[5]),
    .SE(n1229),
    .SI(n1091));
 XNOR2xp5_ASAP7_75t_SL i990 (.A(n0[36]),
    .B(n35[4]),
    .Y(n427));
 XNOR2xp5_ASAP7_75t_SL i991 (.A(n0[80]),
    .B(n36[16]),
    .Y(n426));
 XNOR2xp5_ASAP7_75t_SL i992 (.A(n0[35]),
    .B(n35[3]),
    .Y(n425));
 XNOR2xp5_ASAP7_75t_SL i993 (.A(n0[89]),
    .B(n36[25]),
    .Y(n424));
 XNOR2xp5_ASAP7_75t_SL i994 (.A(n0[119]),
    .B(n37[23]),
    .Y(n423));
 XNOR2xp5_ASAP7_75t_SL i995 (.A(n0[127]),
    .B(n37[31]),
    .Y(n422));
 XNOR2xp5_ASAP7_75t_SL i996 (.A(n0[32]),
    .B(n35[0]),
    .Y(n421));
 XNOR2xp5_ASAP7_75t_SL i997 (.A(n0[71]),
    .B(n36[7]),
    .Y(n420));
 XNOR2xp5_ASAP7_75t_SL i998 (.A(n0[70]),
    .B(n36[6]),
    .Y(n419));
 XNOR2xp5_ASAP7_75t_SL i999 (.A(n0[69]),
    .B(n36[5]),
    .Y(n418));
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_208_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_207_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_206_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_205_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_204_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_203_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_202_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_201_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_200_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_199_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_198_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_197_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_196_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_195_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_194_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_193_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_192_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_191_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_190_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_189_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_188_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_187_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_186_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_185_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_184_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_183_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_182_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_181_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_180_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_179_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_178_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_177_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_176_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_175_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_174_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_173_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_172_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_171_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_170_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_169_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_168_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_167_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_166_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_165_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_164_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_163_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_162_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_161_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_160_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_159_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_158_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_157_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_156_Right_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_155_Right_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_154_Right_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_153_Right_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_152_Right_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_151_Right_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_150_Right_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_149_Right_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_148_Right_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_147_Right_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_146_Right_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_145_Right_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_144_Right_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_143_Right_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_142_Right_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_141_Right_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_140_Right_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_139_Right_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_138_Right_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_137_Right_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_136_Right_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_135_Right_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_134_Right_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_133_Right_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_132_Right_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_131_Right_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_130_Right_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_129_Right_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_128_Right_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_127_Right_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_126_Right_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_125_Right_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_124_Right_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_123_Right_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_122_Right_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_121_Right_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_120_Right_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_119_Right_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_118_Right_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_117_Right_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_116_Right_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_115_Right_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_114_Right_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_113_Right_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_112_Right_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_111_Right_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_110_Right_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_109_Right_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_108_Right_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_107_Right_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_106_Right_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_105_Right_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_104_Right_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_103_Right_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_102_Right_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_101_Right_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_100_Right_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_99_Right_109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_98_Right_110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_97_Right_111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_96_Right_112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_95_Right_113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_94_Right_114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_93_Right_115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_92_Right_116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_91_Right_117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_90_Right_118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_89_Right_119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_88_Right_120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_87_Right_121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_86_Right_122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_85_Right_123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_84_Right_124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_83_Right_125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_82_Right_126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_81_Right_127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_80_Right_128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_79_Right_129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_78_Right_130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_77_Right_131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_76_Right_132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_75_Right_133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_74_Right_134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_73_Right_135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_72_Right_136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_71_Right_137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_70_Right_138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_69_Right_139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_68_Right_140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_67_Right_141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_66_Right_142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_65_Right_143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_64_Right_144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_63_Right_145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_62_Right_146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_61_Right_147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_60_Right_148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_59_Right_149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_58_Right_150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_57_Right_151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_56_Right_152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_55_Right_153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_54_Right_154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_53_Right_155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_52_Right_156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_51_Right_157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_50_Right_158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_49_Right_159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_48_Right_160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_47_Right_161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_46_Right_162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_45_Right_163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_44_Right_164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_43_Right_165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_42_Right_166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_41_Right_167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_40_Right_168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_39_Right_169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_38_Right_170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_37_Right_171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_36_Right_172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_35_Right_173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_34_Right_174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_33_Right_175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_32_Right_176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_31_Right_177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_30_Right_178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_29_Right_179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_28_Right_180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_27_Right_181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_26_Right_182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_25_Right_183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_24_Right_184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_23_Right_185 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_22_Right_186 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_21_Right_187 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_20_Right_188 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_19_Right_189 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_18_Right_190 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_17_Right_191 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_16_Right_192 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_15_Right_193 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_14_Right_194 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_13_Right_195 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_12_Right_196 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_11_Right_197 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_10_Right_198 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_9_Right_199 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_8_Right_200 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_7_Right_201 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_6_Right_202 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_5_Right_203 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_4_Right_204 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_3_Right_205 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_2_Right_206 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_1_Right_207 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_0_Right_208 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_208_Left_209 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_207_Left_210 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_206_Left_211 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_205_Left_212 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_204_Left_213 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_203_Left_214 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_202_Left_215 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_201_Left_216 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_200_Left_217 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_199_Left_218 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_198_Left_219 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_197_Left_220 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_196_Left_221 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_195_Left_222 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_194_Left_223 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_193_Left_224 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_192_Left_225 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_191_Left_226 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_190_Left_227 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_189_Left_228 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_188_Left_229 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_187_Left_230 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_186_Left_231 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_185_Left_232 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_184_Left_233 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_183_Left_234 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_182_Left_235 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_181_Left_236 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_180_Left_237 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_179_Left_238 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_178_Left_239 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_177_Left_240 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_176_Left_241 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_175_Left_242 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_174_Left_243 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_173_Left_244 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_172_Left_245 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_171_Left_246 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_170_Left_247 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_169_Left_248 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_168_Left_249 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_167_Left_250 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_166_Left_251 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_165_Left_252 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_164_Left_253 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_163_Left_254 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_162_Left_255 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_161_Left_256 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_160_Left_257 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_159_Left_258 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_158_Left_259 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_157_Left_260 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_156_Left_261 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_155_Left_262 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_154_Left_263 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_153_Left_264 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_152_Left_265 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_151_Left_266 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_150_Left_267 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_149_Left_268 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_148_Left_269 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_147_Left_270 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_146_Left_271 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_145_Left_272 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_144_Left_273 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_143_Left_274 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_142_Left_275 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_141_Left_276 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_140_Left_277 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_139_Left_278 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_138_Left_279 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_137_Left_280 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_136_Left_281 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_135_Left_282 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_134_Left_283 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_133_Left_284 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_132_Left_285 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_131_Left_286 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_130_Left_287 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_129_Left_288 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_128_Left_289 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_127_Left_290 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_126_Left_291 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_125_Left_292 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_124_Left_293 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_123_Left_294 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_122_Left_295 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_121_Left_296 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_120_Left_297 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_119_Left_298 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_118_Left_299 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_117_Left_300 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_116_Left_301 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_115_Left_302 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_114_Left_303 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_113_Left_304 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_112_Left_305 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_111_Left_306 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_110_Left_307 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_109_Left_308 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_108_Left_309 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_107_Left_310 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_106_Left_311 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_105_Left_312 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_104_Left_313 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_103_Left_314 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_102_Left_315 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_101_Left_316 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_100_Left_317 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_99_Left_318 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_98_Left_319 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_97_Left_320 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_96_Left_321 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_95_Left_322 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_94_Left_323 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_93_Left_324 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_92_Left_325 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_91_Left_326 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_90_Left_327 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_89_Left_328 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_88_Left_329 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_87_Left_330 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_86_Left_331 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_85_Left_332 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_84_Left_333 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_83_Left_334 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_82_Left_335 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_81_Left_336 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_80_Left_337 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_79_Left_338 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_78_Left_339 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_77_Left_340 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_76_Left_341 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_75_Left_342 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_74_Left_343 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_73_Left_344 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_72_Left_345 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_71_Left_346 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_70_Left_347 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_69_Left_348 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_68_Left_349 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_67_Left_350 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_66_Left_351 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_65_Left_352 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_64_Left_353 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_63_Left_354 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_62_Left_355 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_61_Left_356 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_60_Left_357 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_59_Left_358 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_58_Left_359 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_57_Left_360 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_56_Left_361 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_55_Left_362 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_54_Left_363 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_53_Left_364 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_52_Left_365 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_51_Left_366 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_50_Left_367 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_49_Left_368 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_48_Left_369 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_47_Left_370 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_46_Left_371 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_45_Left_372 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_44_Left_373 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_43_Left_374 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_42_Left_375 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_41_Left_376 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_40_Left_377 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_39_Left_378 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_38_Left_379 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_37_Left_380 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_36_Left_381 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_35_Left_382 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_34_Left_383 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_33_Left_384 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_32_Left_385 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_31_Left_386 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_30_Left_387 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_29_Left_388 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_28_Left_389 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_27_Left_390 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_26_Left_391 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_25_Left_392 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_24_Left_393 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_23_Left_394 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_22_Left_395 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_21_Left_396 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_20_Left_397 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_19_Left_398 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_18_Left_399 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_17_Left_400 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_16_Left_401 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_15_Left_402 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_14_Left_403 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_13_Left_404 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_12_Left_405 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_11_Left_406 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_10_Left_407 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_9_Left_408 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_8_Left_409 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_7_Left_410 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_6_Left_411 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_5_Left_412 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_4_Left_413 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_3_Left_414 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_2_Left_415 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_1_Left_416 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_CORE_ROW_0_Left_417 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_208_418 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_208_419 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_207_420 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_206_421 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_205_422 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_204_423 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_203_424 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_202_425 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_201_426 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_200_427 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_199_428 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_198_429 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_197_430 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_196_431 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_195_432 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_194_433 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_193_434 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_192_435 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_191_436 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_190_437 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_189_438 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_188_439 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_187_440 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_186_441 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_185_442 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_184_443 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_183_444 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_182_445 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_181_446 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_180_447 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_179_448 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_178_449 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_177_450 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_176_451 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_175_452 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_174_453 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_173_454 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_172_455 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_171_456 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_170_457 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_169_458 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_168_459 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_167_460 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_166_461 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_165_462 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_164_463 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_163_464 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_162_465 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_161_466 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_160_467 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_159_468 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_158_469 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_157_470 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_156_471 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_155_472 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_154_473 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_153_474 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_152_475 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_151_476 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_150_477 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_149_478 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_148_479 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_147_480 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_146_481 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_145_482 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_144_483 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_143_484 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_142_485 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_141_486 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_140_487 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_139_488 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_138_489 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_137_490 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_136_491 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_135_492 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_134_493 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_133_494 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_132_495 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_131_496 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_130_497 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_129_498 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_128_499 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_127_500 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_126_501 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_125_502 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_124_503 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_123_504 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_122_505 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_121_506 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_120_507 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_119_508 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_118_509 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_117_510 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_116_511 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_115_512 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_114_513 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_113_514 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_112_515 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_111_516 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_110_517 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_109_518 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_108_519 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_107_520 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_106_521 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_105_522 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_104_523 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_103_524 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_102_525 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_101_526 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_100_527 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_99_528 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_98_529 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_97_530 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_96_531 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_95_532 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_94_533 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_93_534 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_92_535 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_91_536 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_90_537 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_89_538 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_88_539 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_87_540 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_86_541 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_85_542 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_84_543 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_83_544 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_82_545 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_81_546 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_80_547 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_79_548 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_78_549 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_77_550 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_76_551 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_75_552 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_74_553 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_73_554 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_72_555 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_71_556 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_70_557 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_69_558 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_68_559 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_67_560 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_66_561 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_65_562 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_64_563 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_63_564 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_62_565 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_61_566 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_60_567 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_59_568 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_58_569 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_57_570 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_56_571 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_55_572 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_54_573 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_53_574 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_52_575 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_51_576 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_50_577 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_49_578 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_48_579 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_47_580 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_46_581 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_45_582 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_44_583 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_43_584 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_42_585 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_41_586 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_40_587 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_39_588 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_38_589 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_37_590 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_36_591 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_35_592 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_34_593 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_33_594 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_32_595 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_31_596 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_30_597 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_29_598 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_28_599 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_27_600 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_26_601 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_25_602 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_24_603 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_23_604 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_22_605 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_21_606 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_20_607 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_19_608 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_18_609 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_17_610 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_16_611 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_15_612 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_14_613 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_13_614 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_12_615 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_11_616 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_10_617 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_9_618 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_8_619 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_7_620 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_6_621 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_5_622 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_4_623 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_3_624 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_2_625 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_1_626 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_0_627 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_CORE_ROW_0_628 ();
 BUFx2_ASAP7_75t_L input1 (.A(key[0]),
    .Y(net1));
 BUFx2_ASAP7_75t_L input2 (.A(key[100]),
    .Y(net2));
 BUFx2_ASAP7_75t_L input3 (.A(key[101]),
    .Y(net3));
 BUFx2_ASAP7_75t_L input4 (.A(key[102]),
    .Y(net4));
 BUFx2_ASAP7_75t_L input5 (.A(key[103]),
    .Y(net5));
 BUFx2_ASAP7_75t_L input6 (.A(key[104]),
    .Y(net6));
 BUFx2_ASAP7_75t_L input7 (.A(key[105]),
    .Y(net7));
 BUFx2_ASAP7_75t_L input8 (.A(key[106]),
    .Y(net8));
 BUFx2_ASAP7_75t_L input9 (.A(key[107]),
    .Y(net9));
 BUFx2_ASAP7_75t_L input10 (.A(key[108]),
    .Y(net10));
 BUFx2_ASAP7_75t_L input11 (.A(key[109]),
    .Y(net11));
 BUFx2_ASAP7_75t_L input12 (.A(key[10]),
    .Y(net12));
 BUFx2_ASAP7_75t_L input13 (.A(key[110]),
    .Y(net13));
 BUFx2_ASAP7_75t_L input14 (.A(key[111]),
    .Y(net14));
 BUFx2_ASAP7_75t_L input15 (.A(key[112]),
    .Y(net15));
 BUFx2_ASAP7_75t_L input16 (.A(key[113]),
    .Y(net16));
 BUFx2_ASAP7_75t_L input17 (.A(key[114]),
    .Y(net17));
 BUFx2_ASAP7_75t_L input18 (.A(key[115]),
    .Y(net18));
 BUFx2_ASAP7_75t_L input19 (.A(key[116]),
    .Y(net19));
 BUFx2_ASAP7_75t_L input20 (.A(key[117]),
    .Y(net20));
 BUFx2_ASAP7_75t_L input21 (.A(key[118]),
    .Y(net21));
 BUFx2_ASAP7_75t_L input22 (.A(key[119]),
    .Y(net22));
 BUFx2_ASAP7_75t_L input23 (.A(key[11]),
    .Y(net23));
 BUFx2_ASAP7_75t_L input24 (.A(key[120]),
    .Y(net24));
 BUFx2_ASAP7_75t_L input25 (.A(key[121]),
    .Y(net25));
 BUFx2_ASAP7_75t_L input26 (.A(key[122]),
    .Y(net26));
 BUFx2_ASAP7_75t_L input27 (.A(key[123]),
    .Y(net27));
 BUFx2_ASAP7_75t_L input28 (.A(key[124]),
    .Y(net28));
 BUFx2_ASAP7_75t_L input29 (.A(key[125]),
    .Y(net29));
 BUFx2_ASAP7_75t_L input30 (.A(key[126]),
    .Y(net30));
 BUFx2_ASAP7_75t_L input31 (.A(key[127]),
    .Y(net31));
 BUFx2_ASAP7_75t_L input32 (.A(key[12]),
    .Y(net32));
 BUFx2_ASAP7_75t_L input33 (.A(key[13]),
    .Y(net33));
 BUFx2_ASAP7_75t_L input34 (.A(key[14]),
    .Y(net34));
 BUFx2_ASAP7_75t_L input35 (.A(key[15]),
    .Y(net35));
 BUFx2_ASAP7_75t_L input36 (.A(key[16]),
    .Y(net36));
 BUFx2_ASAP7_75t_L input37 (.A(key[17]),
    .Y(net37));
 BUFx2_ASAP7_75t_L input38 (.A(key[18]),
    .Y(net38));
 BUFx2_ASAP7_75t_L input39 (.A(key[19]),
    .Y(net39));
 BUFx2_ASAP7_75t_L input40 (.A(key[1]),
    .Y(net40));
 BUFx2_ASAP7_75t_L input41 (.A(key[20]),
    .Y(net41));
 BUFx2_ASAP7_75t_L input42 (.A(key[21]),
    .Y(net42));
 BUFx2_ASAP7_75t_L input43 (.A(key[22]),
    .Y(net43));
 BUFx2_ASAP7_75t_L input44 (.A(key[23]),
    .Y(net44));
 BUFx2_ASAP7_75t_L input45 (.A(key[24]),
    .Y(net45));
 BUFx2_ASAP7_75t_L input46 (.A(key[25]),
    .Y(net46));
 BUFx2_ASAP7_75t_L input47 (.A(key[26]),
    .Y(net47));
 BUFx2_ASAP7_75t_L input48 (.A(key[27]),
    .Y(net48));
 BUFx2_ASAP7_75t_L input49 (.A(key[28]),
    .Y(net49));
 BUFx2_ASAP7_75t_L input50 (.A(key[29]),
    .Y(net50));
 BUFx2_ASAP7_75t_L input51 (.A(key[2]),
    .Y(net51));
 BUFx2_ASAP7_75t_L input52 (.A(key[30]),
    .Y(net52));
 BUFx2_ASAP7_75t_L input53 (.A(key[31]),
    .Y(net53));
 BUFx2_ASAP7_75t_L input54 (.A(key[32]),
    .Y(net54));
 BUFx2_ASAP7_75t_L input55 (.A(key[33]),
    .Y(net55));
 BUFx2_ASAP7_75t_L input56 (.A(key[34]),
    .Y(net56));
 BUFx2_ASAP7_75t_L input57 (.A(key[35]),
    .Y(net57));
 BUFx2_ASAP7_75t_L input58 (.A(key[36]),
    .Y(net58));
 BUFx2_ASAP7_75t_L input59 (.A(key[37]),
    .Y(net59));
 BUFx2_ASAP7_75t_L input60 (.A(key[38]),
    .Y(net60));
 BUFx2_ASAP7_75t_L input61 (.A(key[39]),
    .Y(net61));
 BUFx2_ASAP7_75t_L input62 (.A(key[3]),
    .Y(net62));
 BUFx2_ASAP7_75t_L input63 (.A(key[40]),
    .Y(net63));
 BUFx2_ASAP7_75t_L input64 (.A(key[41]),
    .Y(net64));
 BUFx2_ASAP7_75t_L input65 (.A(key[42]),
    .Y(net65));
 BUFx2_ASAP7_75t_L input66 (.A(key[43]),
    .Y(net66));
 BUFx2_ASAP7_75t_L input67 (.A(key[44]),
    .Y(net67));
 BUFx2_ASAP7_75t_L input68 (.A(key[45]),
    .Y(net68));
 BUFx2_ASAP7_75t_L input69 (.A(key[46]),
    .Y(net69));
 BUFx2_ASAP7_75t_L input70 (.A(key[47]),
    .Y(net70));
 BUFx2_ASAP7_75t_L input71 (.A(key[48]),
    .Y(net71));
 BUFx2_ASAP7_75t_L input72 (.A(key[49]),
    .Y(net72));
 BUFx2_ASAP7_75t_L input73 (.A(key[4]),
    .Y(net73));
 BUFx2_ASAP7_75t_L input74 (.A(key[50]),
    .Y(net74));
 BUFx2_ASAP7_75t_L input75 (.A(key[51]),
    .Y(net75));
 BUFx2_ASAP7_75t_L input76 (.A(key[52]),
    .Y(net76));
 BUFx2_ASAP7_75t_L input77 (.A(key[53]),
    .Y(net77));
 BUFx2_ASAP7_75t_L input78 (.A(key[54]),
    .Y(net78));
 BUFx2_ASAP7_75t_L input79 (.A(key[55]),
    .Y(net79));
 BUFx2_ASAP7_75t_L input80 (.A(key[56]),
    .Y(net80));
 BUFx2_ASAP7_75t_L input81 (.A(key[57]),
    .Y(net81));
 BUFx2_ASAP7_75t_L input82 (.A(key[58]),
    .Y(net82));
 BUFx2_ASAP7_75t_L input83 (.A(key[59]),
    .Y(net83));
 BUFx2_ASAP7_75t_L input84 (.A(key[5]),
    .Y(net84));
 BUFx2_ASAP7_75t_L input85 (.A(key[60]),
    .Y(net85));
 BUFx2_ASAP7_75t_L input86 (.A(key[61]),
    .Y(net86));
 BUFx2_ASAP7_75t_L input87 (.A(key[62]),
    .Y(net87));
 BUFx2_ASAP7_75t_L input88 (.A(key[63]),
    .Y(net88));
 BUFx2_ASAP7_75t_L input89 (.A(key[64]),
    .Y(net89));
 BUFx2_ASAP7_75t_L input90 (.A(key[65]),
    .Y(net90));
 BUFx2_ASAP7_75t_L input91 (.A(key[66]),
    .Y(net91));
 BUFx2_ASAP7_75t_L input92 (.A(key[67]),
    .Y(net92));
 BUFx2_ASAP7_75t_L input93 (.A(key[68]),
    .Y(net93));
 BUFx2_ASAP7_75t_L input94 (.A(key[69]),
    .Y(net94));
 BUFx2_ASAP7_75t_L input95 (.A(key[6]),
    .Y(net95));
 BUFx2_ASAP7_75t_L input96 (.A(key[70]),
    .Y(net96));
 BUFx2_ASAP7_75t_L input97 (.A(key[71]),
    .Y(net97));
 BUFx2_ASAP7_75t_L input98 (.A(key[72]),
    .Y(net98));
 BUFx2_ASAP7_75t_L input99 (.A(key[73]),
    .Y(net99));
 BUFx2_ASAP7_75t_L input100 (.A(key[74]),
    .Y(net100));
 BUFx2_ASAP7_75t_L input101 (.A(key[75]),
    .Y(net101));
 BUFx2_ASAP7_75t_L input102 (.A(key[76]),
    .Y(net102));
 BUFx2_ASAP7_75t_L input103 (.A(key[77]),
    .Y(net103));
 BUFx2_ASAP7_75t_L input104 (.A(key[78]),
    .Y(net104));
 BUFx2_ASAP7_75t_L input105 (.A(key[79]),
    .Y(net105));
 BUFx2_ASAP7_75t_L input106 (.A(key[7]),
    .Y(net106));
 BUFx2_ASAP7_75t_L input107 (.A(key[80]),
    .Y(net107));
 BUFx2_ASAP7_75t_L input108 (.A(key[81]),
    .Y(net108));
 BUFx2_ASAP7_75t_L input109 (.A(key[82]),
    .Y(net109));
 BUFx2_ASAP7_75t_L input110 (.A(key[83]),
    .Y(net110));
 BUFx2_ASAP7_75t_L input111 (.A(key[84]),
    .Y(net111));
 BUFx2_ASAP7_75t_L input112 (.A(key[85]),
    .Y(net112));
 BUFx2_ASAP7_75t_L input113 (.A(key[86]),
    .Y(net113));
 BUFx2_ASAP7_75t_L input114 (.A(key[87]),
    .Y(net114));
 BUFx2_ASAP7_75t_L input115 (.A(key[88]),
    .Y(net115));
 BUFx2_ASAP7_75t_L input116 (.A(key[89]),
    .Y(net116));
 BUFx2_ASAP7_75t_L input117 (.A(key[8]),
    .Y(net117));
 BUFx2_ASAP7_75t_L input118 (.A(key[90]),
    .Y(net118));
 BUFx2_ASAP7_75t_L input119 (.A(key[91]),
    .Y(net119));
 BUFx2_ASAP7_75t_L input120 (.A(key[92]),
    .Y(net120));
 BUFx2_ASAP7_75t_L input121 (.A(key[93]),
    .Y(net121));
 BUFx2_ASAP7_75t_L input122 (.A(key[94]),
    .Y(net122));
 BUFx2_ASAP7_75t_L input123 (.A(key[95]),
    .Y(net123));
 BUFx2_ASAP7_75t_L input124 (.A(key[96]),
    .Y(net124));
 BUFx2_ASAP7_75t_L input125 (.A(key[97]),
    .Y(net125));
 BUFx2_ASAP7_75t_L input126 (.A(key[98]),
    .Y(net126));
 BUFx2_ASAP7_75t_L input127 (.A(key[99]),
    .Y(net127));
 BUFx2_ASAP7_75t_L input128 (.A(key[9]),
    .Y(net128));
 BUFx2_ASAP7_75t_L input129 (.A(ld),
    .Y(net129));
 BUFx2_ASAP7_75t_L input130 (.A(rst),
    .Y(net130));
 BUFx2_ASAP7_75t_L input131 (.A(text_in[0]),
    .Y(net131));
 BUFx2_ASAP7_75t_L input132 (.A(text_in[100]),
    .Y(net132));
 BUFx2_ASAP7_75t_L input133 (.A(text_in[101]),
    .Y(net133));
 BUFx2_ASAP7_75t_L input134 (.A(text_in[102]),
    .Y(net134));
 BUFx2_ASAP7_75t_L input135 (.A(text_in[103]),
    .Y(net135));
 BUFx2_ASAP7_75t_L input136 (.A(text_in[104]),
    .Y(net136));
 BUFx2_ASAP7_75t_L input137 (.A(text_in[105]),
    .Y(net137));
 BUFx2_ASAP7_75t_L input138 (.A(text_in[106]),
    .Y(net138));
 BUFx2_ASAP7_75t_L input139 (.A(text_in[107]),
    .Y(net139));
 BUFx2_ASAP7_75t_L input140 (.A(text_in[108]),
    .Y(net140));
 BUFx2_ASAP7_75t_L input141 (.A(text_in[109]),
    .Y(net141));
 BUFx2_ASAP7_75t_L input142 (.A(text_in[10]),
    .Y(net142));
 BUFx2_ASAP7_75t_L input143 (.A(text_in[110]),
    .Y(net143));
 BUFx2_ASAP7_75t_L input144 (.A(text_in[111]),
    .Y(net144));
 BUFx2_ASAP7_75t_L input145 (.A(text_in[112]),
    .Y(net145));
 BUFx2_ASAP7_75t_L input146 (.A(text_in[113]),
    .Y(net146));
 BUFx2_ASAP7_75t_L input147 (.A(text_in[114]),
    .Y(net147));
 BUFx2_ASAP7_75t_L input148 (.A(text_in[115]),
    .Y(net148));
 BUFx2_ASAP7_75t_L input149 (.A(text_in[116]),
    .Y(net149));
 BUFx2_ASAP7_75t_L input150 (.A(text_in[117]),
    .Y(net150));
 BUFx2_ASAP7_75t_L input151 (.A(text_in[118]),
    .Y(net151));
 BUFx2_ASAP7_75t_L input152 (.A(text_in[119]),
    .Y(net152));
 BUFx2_ASAP7_75t_L input153 (.A(text_in[11]),
    .Y(net153));
 BUFx2_ASAP7_75t_L input154 (.A(text_in[120]),
    .Y(net154));
 BUFx2_ASAP7_75t_L input155 (.A(text_in[121]),
    .Y(net155));
 BUFx2_ASAP7_75t_L input156 (.A(text_in[122]),
    .Y(net156));
 BUFx2_ASAP7_75t_L input157 (.A(text_in[123]),
    .Y(net157));
 BUFx2_ASAP7_75t_L input158 (.A(text_in[124]),
    .Y(net158));
 BUFx2_ASAP7_75t_L input159 (.A(text_in[125]),
    .Y(net159));
 BUFx2_ASAP7_75t_L input160 (.A(text_in[126]),
    .Y(net160));
 BUFx2_ASAP7_75t_L input161 (.A(text_in[127]),
    .Y(net161));
 BUFx2_ASAP7_75t_L input162 (.A(text_in[12]),
    .Y(net162));
 BUFx2_ASAP7_75t_L input163 (.A(text_in[13]),
    .Y(net163));
 BUFx2_ASAP7_75t_L input164 (.A(text_in[14]),
    .Y(net164));
 BUFx2_ASAP7_75t_L input165 (.A(text_in[15]),
    .Y(net165));
 BUFx2_ASAP7_75t_L input166 (.A(text_in[16]),
    .Y(net166));
 BUFx2_ASAP7_75t_L input167 (.A(text_in[17]),
    .Y(net167));
 BUFx2_ASAP7_75t_L input168 (.A(text_in[18]),
    .Y(net168));
 BUFx2_ASAP7_75t_L input169 (.A(text_in[19]),
    .Y(net169));
 BUFx2_ASAP7_75t_L input170 (.A(text_in[1]),
    .Y(net170));
 BUFx2_ASAP7_75t_L input171 (.A(text_in[20]),
    .Y(net171));
 BUFx2_ASAP7_75t_L input172 (.A(text_in[21]),
    .Y(net172));
 BUFx2_ASAP7_75t_L input173 (.A(text_in[22]),
    .Y(net173));
 BUFx2_ASAP7_75t_L input174 (.A(text_in[23]),
    .Y(net174));
 BUFx2_ASAP7_75t_L input175 (.A(text_in[24]),
    .Y(net175));
 BUFx2_ASAP7_75t_L input176 (.A(text_in[25]),
    .Y(net176));
 BUFx2_ASAP7_75t_L input177 (.A(text_in[26]),
    .Y(net177));
 BUFx2_ASAP7_75t_L input178 (.A(text_in[27]),
    .Y(net178));
 BUFx2_ASAP7_75t_L input179 (.A(text_in[28]),
    .Y(net179));
 BUFx2_ASAP7_75t_L input180 (.A(text_in[29]),
    .Y(net180));
 BUFx2_ASAP7_75t_L input181 (.A(text_in[2]),
    .Y(net181));
 BUFx2_ASAP7_75t_L input182 (.A(text_in[30]),
    .Y(net182));
 BUFx2_ASAP7_75t_L input183 (.A(text_in[31]),
    .Y(net183));
 BUFx2_ASAP7_75t_L input184 (.A(text_in[32]),
    .Y(net184));
 BUFx2_ASAP7_75t_L input185 (.A(text_in[33]),
    .Y(net185));
 BUFx2_ASAP7_75t_L input186 (.A(text_in[34]),
    .Y(net186));
 BUFx2_ASAP7_75t_L input187 (.A(text_in[35]),
    .Y(net187));
 BUFx2_ASAP7_75t_L input188 (.A(text_in[36]),
    .Y(net188));
 BUFx2_ASAP7_75t_L input189 (.A(text_in[37]),
    .Y(net189));
 BUFx2_ASAP7_75t_L input190 (.A(text_in[38]),
    .Y(net190));
 BUFx2_ASAP7_75t_L input191 (.A(text_in[39]),
    .Y(net191));
 BUFx2_ASAP7_75t_L input192 (.A(text_in[3]),
    .Y(net192));
 BUFx2_ASAP7_75t_L input193 (.A(text_in[40]),
    .Y(net193));
 BUFx2_ASAP7_75t_L input194 (.A(text_in[41]),
    .Y(net194));
 BUFx2_ASAP7_75t_L input195 (.A(text_in[42]),
    .Y(net195));
 BUFx2_ASAP7_75t_L input196 (.A(text_in[43]),
    .Y(net196));
 BUFx2_ASAP7_75t_L input197 (.A(text_in[44]),
    .Y(net197));
 BUFx2_ASAP7_75t_L input198 (.A(text_in[45]),
    .Y(net198));
 BUFx2_ASAP7_75t_L input199 (.A(text_in[46]),
    .Y(net199));
 BUFx2_ASAP7_75t_L input200 (.A(text_in[47]),
    .Y(net200));
 BUFx2_ASAP7_75t_L input201 (.A(text_in[48]),
    .Y(net201));
 BUFx2_ASAP7_75t_L input202 (.A(text_in[49]),
    .Y(net202));
 BUFx2_ASAP7_75t_L input203 (.A(text_in[4]),
    .Y(net203));
 BUFx2_ASAP7_75t_L input204 (.A(text_in[50]),
    .Y(net204));
 BUFx2_ASAP7_75t_L input205 (.A(text_in[51]),
    .Y(net205));
 BUFx2_ASAP7_75t_L input206 (.A(text_in[52]),
    .Y(net206));
 BUFx2_ASAP7_75t_L input207 (.A(text_in[53]),
    .Y(net207));
 BUFx2_ASAP7_75t_L input208 (.A(text_in[54]),
    .Y(net208));
 BUFx2_ASAP7_75t_L input209 (.A(text_in[55]),
    .Y(net209));
 BUFx2_ASAP7_75t_L input210 (.A(text_in[56]),
    .Y(net210));
 BUFx2_ASAP7_75t_L input211 (.A(text_in[57]),
    .Y(net211));
 BUFx2_ASAP7_75t_L input212 (.A(text_in[58]),
    .Y(net212));
 BUFx2_ASAP7_75t_L input213 (.A(text_in[59]),
    .Y(net213));
 BUFx2_ASAP7_75t_L input214 (.A(text_in[5]),
    .Y(net214));
 BUFx2_ASAP7_75t_L input215 (.A(text_in[60]),
    .Y(net215));
 BUFx2_ASAP7_75t_L input216 (.A(text_in[61]),
    .Y(net216));
 BUFx2_ASAP7_75t_L input217 (.A(text_in[62]),
    .Y(net217));
 BUFx2_ASAP7_75t_L input218 (.A(text_in[63]),
    .Y(net218));
 BUFx2_ASAP7_75t_L input219 (.A(text_in[64]),
    .Y(net219));
 BUFx2_ASAP7_75t_L input220 (.A(text_in[65]),
    .Y(net220));
 BUFx2_ASAP7_75t_L input221 (.A(text_in[66]),
    .Y(net221));
 BUFx2_ASAP7_75t_L input222 (.A(text_in[67]),
    .Y(net222));
 BUFx2_ASAP7_75t_L input223 (.A(text_in[68]),
    .Y(net223));
 BUFx2_ASAP7_75t_L input224 (.A(text_in[69]),
    .Y(net224));
 BUFx2_ASAP7_75t_L input225 (.A(text_in[6]),
    .Y(net225));
 BUFx2_ASAP7_75t_L input226 (.A(text_in[70]),
    .Y(net226));
 BUFx2_ASAP7_75t_L input227 (.A(text_in[71]),
    .Y(net227));
 BUFx2_ASAP7_75t_L input228 (.A(text_in[72]),
    .Y(net228));
 BUFx2_ASAP7_75t_L input229 (.A(text_in[73]),
    .Y(net229));
 BUFx2_ASAP7_75t_L input230 (.A(text_in[74]),
    .Y(net230));
 BUFx2_ASAP7_75t_L input231 (.A(text_in[75]),
    .Y(net231));
 BUFx2_ASAP7_75t_L input232 (.A(text_in[76]),
    .Y(net232));
 BUFx2_ASAP7_75t_L input233 (.A(text_in[77]),
    .Y(net233));
 BUFx2_ASAP7_75t_L input234 (.A(text_in[78]),
    .Y(net234));
 BUFx2_ASAP7_75t_L input235 (.A(text_in[79]),
    .Y(net235));
 BUFx2_ASAP7_75t_L input236 (.A(text_in[7]),
    .Y(net236));
 BUFx2_ASAP7_75t_L input237 (.A(text_in[80]),
    .Y(net237));
 BUFx2_ASAP7_75t_L input238 (.A(text_in[81]),
    .Y(net238));
 BUFx2_ASAP7_75t_L input239 (.A(text_in[82]),
    .Y(net239));
 BUFx2_ASAP7_75t_L input240 (.A(text_in[83]),
    .Y(net240));
 BUFx2_ASAP7_75t_L input241 (.A(text_in[84]),
    .Y(net241));
 BUFx2_ASAP7_75t_L input242 (.A(text_in[85]),
    .Y(net242));
 BUFx2_ASAP7_75t_L input243 (.A(text_in[86]),
    .Y(net243));
 BUFx2_ASAP7_75t_L input244 (.A(text_in[87]),
    .Y(net244));
 BUFx2_ASAP7_75t_L input245 (.A(text_in[88]),
    .Y(net245));
 BUFx2_ASAP7_75t_L input246 (.A(text_in[89]),
    .Y(net246));
 BUFx2_ASAP7_75t_L input247 (.A(text_in[8]),
    .Y(net247));
 BUFx2_ASAP7_75t_L input248 (.A(text_in[90]),
    .Y(net248));
 BUFx2_ASAP7_75t_L input249 (.A(text_in[91]),
    .Y(net249));
 BUFx2_ASAP7_75t_L input250 (.A(text_in[92]),
    .Y(net250));
 BUFx2_ASAP7_75t_L input251 (.A(text_in[93]),
    .Y(net251));
 BUFx2_ASAP7_75t_L input252 (.A(text_in[94]),
    .Y(net252));
 BUFx2_ASAP7_75t_L input253 (.A(text_in[95]),
    .Y(net253));
 BUFx2_ASAP7_75t_L input254 (.A(text_in[96]),
    .Y(net254));
 BUFx2_ASAP7_75t_L input255 (.A(text_in[97]),
    .Y(net255));
 BUFx2_ASAP7_75t_L input256 (.A(text_in[98]),
    .Y(net256));
 BUFx2_ASAP7_75t_L input257 (.A(text_in[99]),
    .Y(net257));
 BUFx2_ASAP7_75t_L input258 (.A(text_in[9]),
    .Y(net258));
 BUFx2_ASAP7_75t_L output259 (.A(net259),
    .Y(done));
 BUFx2_ASAP7_75t_L output260 (.A(net260),
    .Y(text_out[0]));
 BUFx2_ASAP7_75t_L output261 (.A(net261),
    .Y(text_out[100]));
 BUFx2_ASAP7_75t_L output262 (.A(net262),
    .Y(text_out[101]));
 BUFx2_ASAP7_75t_L output263 (.A(net263),
    .Y(text_out[102]));
 BUFx2_ASAP7_75t_L output264 (.A(net264),
    .Y(text_out[103]));
 BUFx2_ASAP7_75t_L output265 (.A(net265),
    .Y(text_out[104]));
 BUFx2_ASAP7_75t_L output266 (.A(net266),
    .Y(text_out[105]));
 BUFx2_ASAP7_75t_L output267 (.A(net267),
    .Y(text_out[106]));
 BUFx2_ASAP7_75t_L output268 (.A(net268),
    .Y(text_out[107]));
 BUFx2_ASAP7_75t_L output269 (.A(net269),
    .Y(text_out[108]));
 BUFx2_ASAP7_75t_L output270 (.A(net270),
    .Y(text_out[109]));
 BUFx2_ASAP7_75t_L output271 (.A(net271),
    .Y(text_out[10]));
 BUFx2_ASAP7_75t_L output272 (.A(net272),
    .Y(text_out[110]));
 BUFx2_ASAP7_75t_L output273 (.A(net273),
    .Y(text_out[111]));
 BUFx2_ASAP7_75t_L output274 (.A(net274),
    .Y(text_out[112]));
 BUFx2_ASAP7_75t_L output275 (.A(net275),
    .Y(text_out[113]));
 BUFx2_ASAP7_75t_L output276 (.A(net276),
    .Y(text_out[114]));
 BUFx2_ASAP7_75t_L output277 (.A(net277),
    .Y(text_out[115]));
 BUFx2_ASAP7_75t_L output278 (.A(net278),
    .Y(text_out[116]));
 BUFx2_ASAP7_75t_L output279 (.A(net279),
    .Y(text_out[117]));
 BUFx2_ASAP7_75t_L output280 (.A(net280),
    .Y(text_out[118]));
 BUFx2_ASAP7_75t_L output281 (.A(net281),
    .Y(text_out[119]));
 BUFx2_ASAP7_75t_L output282 (.A(net282),
    .Y(text_out[11]));
 BUFx2_ASAP7_75t_L output283 (.A(net283),
    .Y(text_out[120]));
 BUFx2_ASAP7_75t_L output284 (.A(net284),
    .Y(text_out[121]));
 BUFx2_ASAP7_75t_L output285 (.A(net285),
    .Y(text_out[122]));
 BUFx2_ASAP7_75t_L output286 (.A(net286),
    .Y(text_out[123]));
 BUFx2_ASAP7_75t_L output287 (.A(net287),
    .Y(text_out[124]));
 BUFx2_ASAP7_75t_L output288 (.A(net288),
    .Y(text_out[125]));
 BUFx2_ASAP7_75t_L output289 (.A(net289),
    .Y(text_out[126]));
 BUFx2_ASAP7_75t_L output290 (.A(net290),
    .Y(text_out[127]));
 BUFx2_ASAP7_75t_L output291 (.A(net291),
    .Y(text_out[12]));
 BUFx2_ASAP7_75t_L output292 (.A(net292),
    .Y(text_out[13]));
 BUFx2_ASAP7_75t_L output293 (.A(net293),
    .Y(text_out[14]));
 BUFx2_ASAP7_75t_L output294 (.A(net294),
    .Y(text_out[15]));
 BUFx2_ASAP7_75t_L output295 (.A(net295),
    .Y(text_out[16]));
 BUFx2_ASAP7_75t_L output296 (.A(net296),
    .Y(text_out[17]));
 BUFx2_ASAP7_75t_L output297 (.A(net297),
    .Y(text_out[18]));
 BUFx2_ASAP7_75t_L output298 (.A(net298),
    .Y(text_out[19]));
 BUFx2_ASAP7_75t_L output299 (.A(net299),
    .Y(text_out[1]));
 BUFx2_ASAP7_75t_L output300 (.A(net300),
    .Y(text_out[20]));
 BUFx2_ASAP7_75t_L output301 (.A(net301),
    .Y(text_out[21]));
 BUFx2_ASAP7_75t_L output302 (.A(net302),
    .Y(text_out[22]));
 BUFx2_ASAP7_75t_L output303 (.A(net303),
    .Y(text_out[23]));
 BUFx2_ASAP7_75t_L output304 (.A(net304),
    .Y(text_out[24]));
 BUFx2_ASAP7_75t_L output305 (.A(net305),
    .Y(text_out[25]));
 BUFx2_ASAP7_75t_L output306 (.A(net306),
    .Y(text_out[26]));
 BUFx2_ASAP7_75t_L output307 (.A(net307),
    .Y(text_out[27]));
 BUFx2_ASAP7_75t_L output308 (.A(net308),
    .Y(text_out[28]));
 BUFx2_ASAP7_75t_L output309 (.A(net309),
    .Y(text_out[29]));
 BUFx2_ASAP7_75t_L output310 (.A(net310),
    .Y(text_out[2]));
 BUFx2_ASAP7_75t_L output311 (.A(net311),
    .Y(text_out[30]));
 BUFx2_ASAP7_75t_L output312 (.A(net312),
    .Y(text_out[31]));
 BUFx2_ASAP7_75t_L output313 (.A(net313),
    .Y(text_out[32]));
 BUFx2_ASAP7_75t_L output314 (.A(net314),
    .Y(text_out[33]));
 BUFx2_ASAP7_75t_L output315 (.A(net315),
    .Y(text_out[34]));
 BUFx2_ASAP7_75t_L output316 (.A(net316),
    .Y(text_out[35]));
 BUFx2_ASAP7_75t_L output317 (.A(net317),
    .Y(text_out[36]));
 BUFx2_ASAP7_75t_L output318 (.A(net318),
    .Y(text_out[37]));
 BUFx2_ASAP7_75t_L output319 (.A(net319),
    .Y(text_out[38]));
 BUFx2_ASAP7_75t_L output320 (.A(net320),
    .Y(text_out[39]));
 BUFx2_ASAP7_75t_L output321 (.A(net321),
    .Y(text_out[3]));
 BUFx2_ASAP7_75t_L output322 (.A(net322),
    .Y(text_out[40]));
 BUFx2_ASAP7_75t_L output323 (.A(net323),
    .Y(text_out[41]));
 BUFx2_ASAP7_75t_L output324 (.A(net324),
    .Y(text_out[42]));
 BUFx2_ASAP7_75t_L output325 (.A(net325),
    .Y(text_out[43]));
 BUFx2_ASAP7_75t_L output326 (.A(net326),
    .Y(text_out[44]));
 BUFx2_ASAP7_75t_L output327 (.A(net327),
    .Y(text_out[45]));
 BUFx2_ASAP7_75t_L output328 (.A(net328),
    .Y(text_out[46]));
 BUFx2_ASAP7_75t_L output329 (.A(net329),
    .Y(text_out[47]));
 BUFx2_ASAP7_75t_L output330 (.A(net330),
    .Y(text_out[48]));
 BUFx2_ASAP7_75t_L output331 (.A(net331),
    .Y(text_out[49]));
 BUFx2_ASAP7_75t_L output332 (.A(net332),
    .Y(text_out[4]));
 BUFx2_ASAP7_75t_L output333 (.A(net333),
    .Y(text_out[50]));
 BUFx2_ASAP7_75t_L output334 (.A(net334),
    .Y(text_out[51]));
 BUFx2_ASAP7_75t_L output335 (.A(net335),
    .Y(text_out[52]));
 BUFx2_ASAP7_75t_L output336 (.A(net336),
    .Y(text_out[53]));
 BUFx2_ASAP7_75t_L output337 (.A(net337),
    .Y(text_out[54]));
 BUFx2_ASAP7_75t_L output338 (.A(net338),
    .Y(text_out[55]));
 BUFx2_ASAP7_75t_L output339 (.A(net339),
    .Y(text_out[56]));
 BUFx2_ASAP7_75t_L output340 (.A(net340),
    .Y(text_out[57]));
 BUFx2_ASAP7_75t_L output341 (.A(net341),
    .Y(text_out[58]));
 BUFx2_ASAP7_75t_L output342 (.A(net342),
    .Y(text_out[59]));
 BUFx2_ASAP7_75t_L output343 (.A(net343),
    .Y(text_out[5]));
 BUFx2_ASAP7_75t_L output344 (.A(net344),
    .Y(text_out[60]));
 BUFx2_ASAP7_75t_L output345 (.A(net345),
    .Y(text_out[61]));
 BUFx2_ASAP7_75t_L output346 (.A(net346),
    .Y(text_out[62]));
 BUFx2_ASAP7_75t_L output347 (.A(net347),
    .Y(text_out[63]));
 BUFx2_ASAP7_75t_L output348 (.A(net348),
    .Y(text_out[64]));
 BUFx2_ASAP7_75t_L output349 (.A(net349),
    .Y(text_out[65]));
 BUFx2_ASAP7_75t_L output350 (.A(net350),
    .Y(text_out[66]));
 BUFx2_ASAP7_75t_L output351 (.A(net351),
    .Y(text_out[67]));
 BUFx2_ASAP7_75t_L output352 (.A(net352),
    .Y(text_out[68]));
 BUFx2_ASAP7_75t_L output353 (.A(net353),
    .Y(text_out[69]));
 BUFx2_ASAP7_75t_L output354 (.A(net354),
    .Y(text_out[6]));
 BUFx2_ASAP7_75t_L output355 (.A(net355),
    .Y(text_out[70]));
 BUFx2_ASAP7_75t_L output356 (.A(net356),
    .Y(text_out[71]));
 BUFx2_ASAP7_75t_L output357 (.A(net357),
    .Y(text_out[72]));
 BUFx2_ASAP7_75t_L output358 (.A(net358),
    .Y(text_out[73]));
 BUFx2_ASAP7_75t_L output359 (.A(net359),
    .Y(text_out[74]));
 BUFx2_ASAP7_75t_L output360 (.A(net360),
    .Y(text_out[75]));
 BUFx2_ASAP7_75t_L output361 (.A(net361),
    .Y(text_out[76]));
 BUFx2_ASAP7_75t_L output362 (.A(net362),
    .Y(text_out[77]));
 BUFx2_ASAP7_75t_L output363 (.A(net363),
    .Y(text_out[78]));
 BUFx2_ASAP7_75t_L output364 (.A(net364),
    .Y(text_out[79]));
 BUFx2_ASAP7_75t_L output365 (.A(net365),
    .Y(text_out[7]));
 BUFx2_ASAP7_75t_L output366 (.A(net366),
    .Y(text_out[80]));
 BUFx2_ASAP7_75t_L output367 (.A(net367),
    .Y(text_out[81]));
 BUFx2_ASAP7_75t_L output368 (.A(net368),
    .Y(text_out[82]));
 BUFx2_ASAP7_75t_L output369 (.A(net369),
    .Y(text_out[83]));
 BUFx2_ASAP7_75t_L output370 (.A(net370),
    .Y(text_out[84]));
 BUFx2_ASAP7_75t_L output371 (.A(net371),
    .Y(text_out[85]));
 BUFx2_ASAP7_75t_L output372 (.A(net372),
    .Y(text_out[86]));
 BUFx2_ASAP7_75t_L output373 (.A(net373),
    .Y(text_out[87]));
 BUFx2_ASAP7_75t_L output374 (.A(net374),
    .Y(text_out[88]));
 BUFx2_ASAP7_75t_L output375 (.A(net375),
    .Y(text_out[89]));
 BUFx2_ASAP7_75t_L output376 (.A(net376),
    .Y(text_out[8]));
 BUFx2_ASAP7_75t_L output377 (.A(net377),
    .Y(text_out[90]));
 BUFx2_ASAP7_75t_L output378 (.A(net378),
    .Y(text_out[91]));
 BUFx2_ASAP7_75t_L output379 (.A(net379),
    .Y(text_out[92]));
 BUFx2_ASAP7_75t_L output380 (.A(net380),
    .Y(text_out[93]));
 BUFx2_ASAP7_75t_L output381 (.A(net381),
    .Y(text_out[94]));
 BUFx2_ASAP7_75t_L output382 (.A(net382),
    .Y(text_out[95]));
 BUFx2_ASAP7_75t_L output383 (.A(net383),
    .Y(text_out[96]));
 BUFx2_ASAP7_75t_L output384 (.A(net384),
    .Y(text_out[97]));
 BUFx2_ASAP7_75t_L output385 (.A(net385),
    .Y(text_out[98]));
 BUFx2_ASAP7_75t_L output386 (.A(net386),
    .Y(text_out[99]));
 BUFx2_ASAP7_75t_L output387 (.A(net387),
    .Y(text_out[9]));
endmodule

module aes_cipher_top (clk,
    done,
    ld,
    rst,
    key,
    text_in,
    text_out);
 input clk;
 output done;
 input ld;
 input rst;
 input [127:0] key;
 input [127:0] text_in;
 output [127:0] text_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00978_;
 wire _00979_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01022_;
 wire _01023_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01108_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01129_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01150_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01171_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01213_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01326_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01347_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01368_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01389_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01727_;
 wire _01729_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01772_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01787_;
 wire _01790_;
 wire _01791_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01803_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01813_;
 wire _01814_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01888_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02375_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02392_;
 wire _02396_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02428_;
 wire _02429_;
 wire _02431_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02443_;
 wire _02444_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02453_;
 wire _02454_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02470_;
 wire _02472_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02541_;
 wire _02542_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03070_;
 wire _03071_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03083_;
 wire _03084_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03106_;
 wire _03107_;
 wire _03112_;
 wire _03113_;
 wire _03117_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03152_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03165_;
 wire _03166_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03179_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03291_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03766_;
 wire _03767_;
 wire _03769_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03869_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03937_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04410_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04451_;
 wire _04452_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04467_;
 wire _04468_;
 wire _04472_;
 wire _04473_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04502_;
 wire _04503_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04510_;
 wire _04512_;
 wire _04513_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04551_;
 wire _04552_;
 wire _04555_;
 wire _04557_;
 wire _04558_;
 wire _04560_;
 wire _04561_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05086_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05106_;
 wire _05107_;
 wire _05109_;
 wire _05112_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05146_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05178_;
 wire _05179_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05231_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05315_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05329_;
 wire _05330_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05778_;
 wire _05779_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05823_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05836_;
 wire _05837_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05846_;
 wire _05847_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05870_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05930_;
 wire _05931_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06482_;
 wire _06483_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06515_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06523_;
 wire _06524_;
 wire _06527_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06533_;
 wire _06534_;
 wire _06537_;
 wire _06538_;
 wire _06540_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06547_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06563_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06587_;
 wire _06589_;
 wire _06590_;
 wire _06592_;
 wire _06594_;
 wire _06595_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07138_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07150_;
 wire _07152_;
 wire _07153_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07212_;
 wire _07214_;
 wire _07215_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07222_;
 wire _07223_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07233_;
 wire _07234_;
 wire _07236_;
 wire _07237_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07263_;
 wire _07264_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07737_;
 wire _07738_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07749_;
 wire _07750_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07761_;
 wire _07762_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07773_;
 wire _07774_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07785_;
 wire _07786_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07797_;
 wire _07798_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07809_;
 wire _07810_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07821_;
 wire _07822_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07833_;
 wire _07834_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07845_;
 wire _07846_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07857_;
 wire _07858_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07869_;
 wire _07870_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _08005_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08017_;
 wire _08018_;
 wire _08020_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08081_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08088_;
 wire _08089_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08107_;
 wire _08108_;
 wire _08110_;
 wire _08111_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08143_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08178_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08191_;
 wire _08193_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08200_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08664_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08733_;
 wire _08734_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08789_;
 wire _08790_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08994_;
 wire _08995_;
 wire _08997_;
 wire _09000_;
 wire _09001_;
 wire _09004_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09037_;
 wire _09039_;
 wire _09041_;
 wire _09042_;
 wire _09044_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09051_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09064_;
 wire _09065_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09084_;
 wire _09085_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09144_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09157_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09204_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09566_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09613_;
 wire _09614_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09660_;
 wire _09661_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09667_;
 wire _09668_;
 wire _09670_;
 wire _09671_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09735_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10123_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10131_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10277_;
 wire _10278_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10678_;
 wire _10679_;
 wire _10681_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10758_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10798_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10810_;
 wire _10812_;
 wire _10813_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10845_;
 wire _10846_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10866_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10895_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10915_;
 wire _10916_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10966_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11492_;
 wire _11493_;
 wire _11495_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11525_;
 wire _11526_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11576_;
 wire _11577_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11666_;
 wire _11668_;
 wire _11669_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12169_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12199_;
 wire _12200_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12219_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12236_;
 wire _12237_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12294_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12311_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12336_;
 wire _12337_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12356_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12881_;
 wire _12882_;
 wire _12884_;
 wire _12885_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12895_;
 wire _12897_;
 wire _12899_;
 wire _12900_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12950_;
 wire _12952_;
 wire _12953_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12961_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12972_;
 wire _12973_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13017_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13072_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13516_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13599_;
 wire _13600_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13660_;
 wire _13662_;
 wire _13663_;
 wire _13665_;
 wire _13666_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13696_;
 wire _13697_;
 wire _13699_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13707_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14232_;
 wire _14233_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14288_;
 wire _14289_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14341_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14349_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14406_;
 wire _14407_;
 wire _14409_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14416_;
 wire _14417_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14438_;
 wire _14440_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14452_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15019_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15025_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15034_;
 wire _15035_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15055_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15071_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15104_;
 wire _15105_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15133_;
 wire _15134_;
 wire _15136_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15169_;
 wire _15171_;
 wire _15173_;
 wire _15174_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire \u0.r0.rcnt[0] ;
 wire \u0.r0.rcnt[1] ;
 wire \u0.r0.rcnt_next[0] ;

 XOR2x2_ASAP7_75t_R _15811_ (.A(_00695_),
    .B(_00934_),
    .Y(_00265_));
 XOR2x2_ASAP7_75t_R _15814_ (.A(_00696_),
    .B(_00945_),
    .Y(_00266_));
 XOR2x2_ASAP7_75t_R _15817_ (.A(_00697_),
    .B(_00956_),
    .Y(_00267_));
 XOR2x2_ASAP7_75t_R _15818_ (.A(_00698_),
    .B(_00959_),
    .Y(_00268_));
 XOR2x2_ASAP7_75t_R _15819_ (.A(_00699_),
    .B(_00960_),
    .Y(_00269_));
 XOR2x2_ASAP7_75t_R _15820_ (.A(_00700_),
    .B(_00961_),
    .Y(_00270_));
 XOR2x2_ASAP7_75t_R _15821_ (.A(_00701_),
    .B(_00962_),
    .Y(_00271_));
 XOR2x2_ASAP7_75t_R _15823_ (.A(_00569_),
    .B(_00963_),
    .Y(_00272_));
 XOR2x2_ASAP7_75t_R _15826_ (.A(_00687_),
    .B(_00902_),
    .Y(_00217_));
 XOR2x2_ASAP7_75t_R _15829_ (.A(_00688_),
    .B(_00913_),
    .Y(_00218_));
 XOR2x2_ASAP7_75t_R _15832_ (.A(_00689_),
    .B(_00924_),
    .Y(_00219_));
 XOR2x2_ASAP7_75t_R _15833_ (.A(_00690_),
    .B(_00927_),
    .Y(_00220_));
 XOR2x2_ASAP7_75t_R _15834_ (.A(_00691_),
    .B(_00928_),
    .Y(_00221_));
 XOR2x2_ASAP7_75t_R _15835_ (.A(_00692_),
    .B(_00929_),
    .Y(_00222_));
 XOR2x2_ASAP7_75t_R _15836_ (.A(_00693_),
    .B(_00930_),
    .Y(_00223_));
 XOR2x2_ASAP7_75t_R _15837_ (.A(_00694_),
    .B(_00931_),
    .Y(_00224_));
 XOR2x2_ASAP7_75t_R _15840_ (.A(_00679_),
    .B(_00870_),
    .Y(_00249_));
 XOR2x2_ASAP7_75t_R _15843_ (.A(_00680_),
    .B(_00881_),
    .Y(_00250_));
 XOR2x2_ASAP7_75t_R _15846_ (.A(_00681_),
    .B(_00892_),
    .Y(_00251_));
 XOR2x2_ASAP7_75t_R _15847_ (.A(_00682_),
    .B(_00895_),
    .Y(_00252_));
 XOR2x2_ASAP7_75t_R _15848_ (.A(_00683_),
    .B(_00896_),
    .Y(_00253_));
 XOR2x2_ASAP7_75t_R _15849_ (.A(_00684_),
    .B(_00897_),
    .Y(_00254_));
 XOR2x2_ASAP7_75t_R _15850_ (.A(_00685_),
    .B(_00898_),
    .Y(_00255_));
 XOR2x2_ASAP7_75t_R _15852_ (.A(_00686_),
    .B(_00899_),
    .Y(_00256_));
 XOR2x2_ASAP7_75t_R _15855_ (.A(_00671_),
    .B(_00838_),
    .Y(_00161_));
 XOR2x2_ASAP7_75t_R _15858_ (.A(_00672_),
    .B(_00849_),
    .Y(_00162_));
 XOR2x2_ASAP7_75t_R _15861_ (.A(_00673_),
    .B(_00860_),
    .Y(_00163_));
 XOR2x2_ASAP7_75t_R _15863_ (.A(_00674_),
    .B(_00863_),
    .Y(_00164_));
 XOR2x2_ASAP7_75t_R _15864_ (.A(_00675_),
    .B(_00864_),
    .Y(_00165_));
 XOR2x2_ASAP7_75t_R _15866_ (.A(_00676_),
    .B(_00865_),
    .Y(_00166_));
 XOR2x2_ASAP7_75t_R _15867_ (.A(_00677_),
    .B(_00866_),
    .Y(_00167_));
 XOR2x2_ASAP7_75t_R _15868_ (.A(_00678_),
    .B(_00867_),
    .Y(_00168_));
 XOR2x2_ASAP7_75t_R _15870_ (.A(_00663_),
    .B(_00964_),
    .Y(_00193_));
 XOR2x2_ASAP7_75t_R _15872_ (.A(_00486_),
    .B(_00664_),
    .Y(_00194_));
 XOR2x2_ASAP7_75t_R _15875_ (.A(_00665_),
    .B(_00935_),
    .Y(_00195_));
 XOR2x2_ASAP7_75t_R _15876_ (.A(_00666_),
    .B(_00936_),
    .Y(_00196_));
 XOR2x2_ASAP7_75t_R _15877_ (.A(_00667_),
    .B(_00937_),
    .Y(_00197_));
 XOR2x2_ASAP7_75t_R _15878_ (.A(_00668_),
    .B(_00938_),
    .Y(_00198_));
 XOR2x2_ASAP7_75t_R _15879_ (.A(_00669_),
    .B(_00939_),
    .Y(_00199_));
 XOR2x2_ASAP7_75t_R _15881_ (.A(_00670_),
    .B(_00940_),
    .Y(_00200_));
 XOR2x2_ASAP7_75t_R _15883_ (.A(_00655_),
    .B(_00932_),
    .Y(_00225_));
 XOR2x2_ASAP7_75t_R _15885_ (.A(_00656_),
    .B(_00933_),
    .Y(_00226_));
 XOR2x2_ASAP7_75t_R _15888_ (.A(_00657_),
    .B(_00903_),
    .Y(_00227_));
 XOR2x2_ASAP7_75t_R _15889_ (.A(_00658_),
    .B(_00904_),
    .Y(_00228_));
 XOR2x2_ASAP7_75t_R _15890_ (.A(_00659_),
    .B(_00905_),
    .Y(_00229_));
 XOR2x2_ASAP7_75t_R _15891_ (.A(_00660_),
    .B(_00906_),
    .Y(_00230_));
 XOR2x2_ASAP7_75t_R _15892_ (.A(_00661_),
    .B(_00907_),
    .Y(_00231_));
 XOR2x2_ASAP7_75t_R _15894_ (.A(_00662_),
    .B(_00908_),
    .Y(_00232_));
 XOR2x2_ASAP7_75t_R _15896_ (.A(_00647_),
    .B(_00900_),
    .Y(_00257_));
 XOR2x2_ASAP7_75t_R _15899_ (.A(_00648_),
    .B(_00901_),
    .Y(_00258_));
 XOR2x2_ASAP7_75t_R _15902_ (.A(_00649_),
    .B(_00871_),
    .Y(_00259_));
 XOR2x2_ASAP7_75t_R _15903_ (.A(_00650_),
    .B(_00872_),
    .Y(_00260_));
 XOR2x2_ASAP7_75t_R _15904_ (.A(_00651_),
    .B(_00873_),
    .Y(_00261_));
 XOR2x2_ASAP7_75t_R _15905_ (.A(_00652_),
    .B(_00874_),
    .Y(_00262_));
 XOR2x2_ASAP7_75t_R _15906_ (.A(_00653_),
    .B(_00875_),
    .Y(_00263_));
 XOR2x2_ASAP7_75t_R _15908_ (.A(_00654_),
    .B(_00876_),
    .Y(_00264_));
 XOR2x2_ASAP7_75t_R _15910_ (.A(_00639_),
    .B(_00868_),
    .Y(_00169_));
 XOR2x2_ASAP7_75t_R _15912_ (.A(_00640_),
    .B(_00869_),
    .Y(_00170_));
 XOR2x2_ASAP7_75t_R _15915_ (.A(_00641_),
    .B(_00839_),
    .Y(_00171_));
 XOR2x2_ASAP7_75t_R _15916_ (.A(_00642_),
    .B(_00840_),
    .Y(_00172_));
 XOR2x2_ASAP7_75t_R _15917_ (.A(_00643_),
    .B(_00841_),
    .Y(_00173_));
 XOR2x2_ASAP7_75t_R _15918_ (.A(_00644_),
    .B(_00842_),
    .Y(_00174_));
 XOR2x2_ASAP7_75t_R _15919_ (.A(_00645_),
    .B(_00843_),
    .Y(_00175_));
 XOR2x2_ASAP7_75t_R _15921_ (.A(_00646_),
    .B(_00844_),
    .Y(_00176_));
 XOR2x2_ASAP7_75t_R _15922_ (.A(_00631_),
    .B(_00941_),
    .Y(_00201_));
 XOR2x2_ASAP7_75t_R _15923_ (.A(_00632_),
    .B(_00942_),
    .Y(_00202_));
 XOR2x2_ASAP7_75t_R _15926_ (.A(_00633_),
    .B(_00943_),
    .Y(_00203_));
 XOR2x2_ASAP7_75t_R _15927_ (.A(_00634_),
    .B(_00944_),
    .Y(_00204_));
 XOR2x2_ASAP7_75t_R _15928_ (.A(_00635_),
    .B(_00946_),
    .Y(_00205_));
 XOR2x2_ASAP7_75t_R _15929_ (.A(_00636_),
    .B(_00947_),
    .Y(_00206_));
 XOR2x2_ASAP7_75t_R _15930_ (.A(_00637_),
    .B(_00948_),
    .Y(_00207_));
 XOR2x2_ASAP7_75t_R _15932_ (.A(_00638_),
    .B(_00949_),
    .Y(_00208_));
 XOR2x2_ASAP7_75t_R _15934_ (.A(_00623_),
    .B(_00909_),
    .Y(_00233_));
 XOR2x2_ASAP7_75t_R _15936_ (.A(_00624_),
    .B(_00910_),
    .Y(_00234_));
 XOR2x2_ASAP7_75t_R _15939_ (.A(_00625_),
    .B(_00911_),
    .Y(_00235_));
 XOR2x2_ASAP7_75t_R _15941_ (.A(_00626_),
    .B(_00912_),
    .Y(_00236_));
 XOR2x2_ASAP7_75t_R _15943_ (.A(_00627_),
    .B(_00914_),
    .Y(_00237_));
 XOR2x2_ASAP7_75t_R _15944_ (.A(_00628_),
    .B(_00915_),
    .Y(_00238_));
 XOR2x2_ASAP7_75t_R _15945_ (.A(_00629_),
    .B(_00916_),
    .Y(_00239_));
 XOR2x2_ASAP7_75t_R _15947_ (.A(_00630_),
    .B(_00917_),
    .Y(_00240_));
 XOR2x2_ASAP7_75t_R _15949_ (.A(_00615_),
    .B(_00877_),
    .Y(_00273_));
 XOR2x2_ASAP7_75t_R _15950_ (.A(_00616_),
    .B(_00878_),
    .Y(_00274_));
 XOR2x2_ASAP7_75t_R _15953_ (.A(_00617_),
    .B(_00879_),
    .Y(_00275_));
 XOR2x2_ASAP7_75t_R _15955_ (.A(_00618_),
    .B(_00880_),
    .Y(_00276_));
 XOR2x2_ASAP7_75t_R _15956_ (.A(_00619_),
    .B(_00882_),
    .Y(_00277_));
 XOR2x2_ASAP7_75t_R _15957_ (.A(_00620_),
    .B(_00883_),
    .Y(_00278_));
 XOR2x2_ASAP7_75t_R _15958_ (.A(_00621_),
    .B(_00884_),
    .Y(_00279_));
 XOR2x2_ASAP7_75t_R _15960_ (.A(_00622_),
    .B(_00885_),
    .Y(_00280_));
 XOR2x2_ASAP7_75t_R _15962_ (.A(_00607_),
    .B(_00845_),
    .Y(_00177_));
 XOR2x2_ASAP7_75t_R _15964_ (.A(_00608_),
    .B(_00846_),
    .Y(_00178_));
 XOR2x2_ASAP7_75t_R _15967_ (.A(_00609_),
    .B(_00847_),
    .Y(_00179_));
 XOR2x2_ASAP7_75t_R _15969_ (.A(_00610_),
    .B(_00848_),
    .Y(_00180_));
 XOR2x2_ASAP7_75t_R _15970_ (.A(_00611_),
    .B(_00850_),
    .Y(_00181_));
 XOR2x2_ASAP7_75t_R _15972_ (.A(_00612_),
    .B(_00851_),
    .Y(_00182_));
 XOR2x2_ASAP7_75t_R _15973_ (.A(_00613_),
    .B(_00852_),
    .Y(_00183_));
 XOR2x2_ASAP7_75t_R _15975_ (.A(_00614_),
    .B(_00853_),
    .Y(_00184_));
 XOR2x2_ASAP7_75t_R _15977_ (.A(_00599_),
    .B(_00950_),
    .Y(_00209_));
 XOR2x2_ASAP7_75t_R _15979_ (.A(_00600_),
    .B(_00951_),
    .Y(_00210_));
 XOR2x2_ASAP7_75t_R _15982_ (.A(_00601_),
    .B(_00952_),
    .Y(_00211_));
 XOR2x2_ASAP7_75t_R _15983_ (.A(_00602_),
    .B(_00953_),
    .Y(_00212_));
 XOR2x2_ASAP7_75t_R _15985_ (.A(_00603_),
    .B(_00954_),
    .Y(_00213_));
 XOR2x2_ASAP7_75t_R _15986_ (.A(_00604_),
    .B(_00955_),
    .Y(_00214_));
 XOR2x2_ASAP7_75t_R _15987_ (.A(_00605_),
    .B(_00957_),
    .Y(_00215_));
 XOR2x2_ASAP7_75t_R _15989_ (.A(_00606_),
    .B(_00958_),
    .Y(_00216_));
 XOR2x2_ASAP7_75t_R _15992_ (.A(_00591_),
    .B(_00918_),
    .Y(_00241_));
 XOR2x2_ASAP7_75t_R _15995_ (.A(_00592_),
    .B(_00919_),
    .Y(_00242_));
 XOR2x2_ASAP7_75t_R _15997_ (.A(_00593_),
    .B(_00920_),
    .Y(_00243_));
 XOR2x2_ASAP7_75t_R _15998_ (.A(_00594_),
    .B(_00921_),
    .Y(_00244_));
 XOR2x2_ASAP7_75t_R _16000_ (.A(_00595_),
    .B(_00922_),
    .Y(_00245_));
 XOR2x2_ASAP7_75t_R _16001_ (.A(_00596_),
    .B(_00923_),
    .Y(_00246_));
 XOR2x2_ASAP7_75t_R _16002_ (.A(_00597_),
    .B(_00925_),
    .Y(_00247_));
 XOR2x2_ASAP7_75t_R _16004_ (.A(_00598_),
    .B(_00926_),
    .Y(_00248_));
 XOR2x2_ASAP7_75t_R _16007_ (.A(_00583_),
    .B(_00886_),
    .Y(_00281_));
 XOR2x2_ASAP7_75t_R _16009_ (.A(_00584_),
    .B(_00887_),
    .Y(_00282_));
 XOR2x2_ASAP7_75t_R _16011_ (.A(_00585_),
    .B(_00888_),
    .Y(_00283_));
 XOR2x2_ASAP7_75t_R _16012_ (.A(_00586_),
    .B(_00889_),
    .Y(_00284_));
 XOR2x2_ASAP7_75t_R _16013_ (.A(_00587_),
    .B(_00890_),
    .Y(_00285_));
 XOR2x2_ASAP7_75t_R _16014_ (.A(_00588_),
    .B(_00891_),
    .Y(_00286_));
 XOR2x2_ASAP7_75t_R _16015_ (.A(_00589_),
    .B(_00893_),
    .Y(_00287_));
 XOR2x2_ASAP7_75t_R _16017_ (.A(_00590_),
    .B(_00894_),
    .Y(_00288_));
 XOR2x2_ASAP7_75t_R _16019_ (.A(_00575_),
    .B(_00854_),
    .Y(_00185_));
 XOR2x2_ASAP7_75t_R _16021_ (.A(_00576_),
    .B(_00855_),
    .Y(_00186_));
 XOR2x2_ASAP7_75t_R _16023_ (.A(_00577_),
    .B(_00856_),
    .Y(_00187_));
 XOR2x2_ASAP7_75t_R _16024_ (.A(_00578_),
    .B(_00857_),
    .Y(_00188_));
 XOR2x2_ASAP7_75t_R _16025_ (.A(_00579_),
    .B(_00858_),
    .Y(_00189_));
 XOR2x2_ASAP7_75t_R _16026_ (.A(_00580_),
    .B(_00859_),
    .Y(_00190_));
 XOR2x2_ASAP7_75t_R _16027_ (.A(_00581_),
    .B(_00861_),
    .Y(_00191_));
 XOR2x2_ASAP7_75t_R _16029_ (.A(_00582_),
    .B(_00862_),
    .Y(_00192_));
 INVx1_ASAP7_75t_SL _16030_ (.A(ld),
    .Y(_08005_));
 INVx1_ASAP7_75t_R _16036_ (.A(_00572_),
    .Y(_08011_));
 AND5x1_ASAP7_75t_R _16037_ (.A(_00411_),
    .B(_08005_),
    .C(_08011_),
    .D(_00570_),
    .E(_00571_),
    .Y(_00160_));
 INVx1_ASAP7_75t_R _16038_ (.A(_00965_),
    .Y(\u0.r0.rcnt[1] ));
 INVx1_ASAP7_75t_R _16039_ (.A(\u0.r0.rcnt_next[0] ),
    .Y(\u0.r0.rcnt[0] ));
 XOR2x2_ASAP7_75t_SL _16040_ (.A(_00440_),
    .B(_00914_),
    .Y(_08012_));
 XOR2x2_ASAP7_75t_R _16041_ (.A(_08012_),
    .B(_00946_),
    .Y(_08013_));
 XOR2x2_ASAP7_75t_R _16042_ (.A(_00850_),
    .B(_00882_),
    .Y(_08014_));
 XOR2x2_ASAP7_75t_SL _16043_ (.A(_08013_),
    .B(_08014_),
    .Y(_08015_));
 NOR2x1_ASAP7_75t_SL _16045_ (.A(key[20]),
    .B(_08005_),
    .Y(_08017_));
 AO21x1_ASAP7_75t_SL _16046_ (.A1(_08015_),
    .A2(_08005_),
    .B(_08017_),
    .Y(_08018_));
 INVx1_ASAP7_75t_SL _16048_ (.A(_08018_),
    .Y(_08020_));
 XOR2x2_ASAP7_75t_R _16051_ (.A(_00441_),
    .B(_00915_),
    .Y(_08022_));
 INVx1_ASAP7_75t_R _16052_ (.A(_00947_),
    .Y(_08023_));
 XOR2x2_ASAP7_75t_R _16053_ (.A(_08022_),
    .B(_08023_),
    .Y(_08024_));
 XNOR2x2_ASAP7_75t_R _16054_ (.A(_00851_),
    .B(_00883_),
    .Y(_08025_));
 XOR2x2_ASAP7_75t_R _16055_ (.A(_08024_),
    .B(_08025_),
    .Y(_08026_));
 NAND2x1_ASAP7_75t_R _16056_ (.A(_08005_),
    .B(_08026_),
    .Y(_08027_));
 OA21x2_ASAP7_75t_R _16057_ (.A1(_08005_),
    .A2(key[21]),
    .B(_08027_),
    .Y(_08028_));
 XOR2x2_ASAP7_75t_SL _16060_ (.A(_00439_),
    .B(_00912_),
    .Y(_08030_));
 INVx1_ASAP7_75t_R _16061_ (.A(_00944_),
    .Y(_08031_));
 XOR2x2_ASAP7_75t_SL _16062_ (.A(_08030_),
    .B(_08031_),
    .Y(_08032_));
 XNOR2x2_ASAP7_75t_R _16063_ (.A(_00848_),
    .B(_00880_),
    .Y(_08033_));
 XOR2x2_ASAP7_75t_SL _16064_ (.A(_08032_),
    .B(_08033_),
    .Y(_08034_));
 NAND2x1_ASAP7_75t_SL _16065_ (.A(_08005_),
    .B(_08034_),
    .Y(_08035_));
 OAI21x1_ASAP7_75t_R _16066_ (.A1(_08005_),
    .A2(key[19]),
    .B(_08035_),
    .Y(_08036_));
 INVx2_ASAP7_75t_SL _16067_ (.A(_08036_),
    .Y(_08037_));
 XOR2x1_ASAP7_75t_SL _16070_ (.A(_00437_),
    .Y(_08039_),
    .B(_00909_));
 INVx1_ASAP7_75t_SL _16071_ (.A(_00941_),
    .Y(_08040_));
 XOR2x2_ASAP7_75t_R _16072_ (.A(_08039_),
    .B(_08040_),
    .Y(_08041_));
 XNOR2x2_ASAP7_75t_R _16073_ (.A(_00845_),
    .B(_00877_),
    .Y(_08042_));
 XOR2x2_ASAP7_75t_SL _16074_ (.A(_08041_),
    .B(_08042_),
    .Y(_08043_));
 NOR2x1_ASAP7_75t_R _16075_ (.A(key[16]),
    .B(_08005_),
    .Y(_08044_));
 AO21x1_ASAP7_75t_R _16076_ (.A1(_08043_),
    .A2(_08005_),
    .B(_08044_),
    .Y(_08045_));
 XOR2x2_ASAP7_75t_SL _16078_ (.A(_00438_),
    .B(_00910_),
    .Y(_08046_));
 INVx1_ASAP7_75t_R _16079_ (.A(_00942_),
    .Y(_08047_));
 XOR2x2_ASAP7_75t_SL _16080_ (.A(_08046_),
    .B(_08047_),
    .Y(_08048_));
 XNOR2x2_ASAP7_75t_R _16081_ (.A(_00846_),
    .B(_00878_),
    .Y(_08049_));
 XOR2x2_ASAP7_75t_SL _16082_ (.A(_08048_),
    .B(_08049_),
    .Y(_08050_));
 NOR2x1_ASAP7_75t_R _16083_ (.A(key[17]),
    .B(_08005_),
    .Y(_08051_));
 AO21x1_ASAP7_75t_SL _16084_ (.A1(_08050_),
    .A2(_08005_),
    .B(_08051_),
    .Y(_08052_));
 AND2x2_ASAP7_75t_R _16087_ (.A(ld),
    .B(key[18]),
    .Y(_08054_));
 INVx1_ASAP7_75t_R _16088_ (.A(_00412_),
    .Y(_08055_));
 XOR2x2_ASAP7_75t_R _16089_ (.A(_00847_),
    .B(_00879_),
    .Y(_08056_));
 XOR2x2_ASAP7_75t_R _16090_ (.A(_00911_),
    .B(_00943_),
    .Y(_08057_));
 XNOR2x1_ASAP7_75t_SL _16091_ (.B(_08057_),
    .Y(_08058_),
    .A(_08056_));
 NOR2x1_ASAP7_75t_R _16092_ (.A(_08055_),
    .B(_08058_),
    .Y(_08059_));
 XOR2x1_ASAP7_75t_L _16093_ (.A(_08056_),
    .Y(_08060_),
    .B(_08057_));
 NOR2x1_ASAP7_75t_SL _16094_ (.A(_00412_),
    .B(_08060_),
    .Y(_08061_));
 OA21x2_ASAP7_75t_SL _16095_ (.A1(_08059_),
    .A2(_08061_),
    .B(_08005_),
    .Y(_08062_));
 NOR2x1_ASAP7_75t_SL _16096_ (.A(_08054_),
    .B(_08062_),
    .Y(_08063_));
 INVx3_ASAP7_75t_SL _16098_ (.A(_08063_),
    .Y(_00989_));
 XOR2x2_ASAP7_75t_R _16100_ (.A(_00442_),
    .B(_00916_),
    .Y(_08066_));
 XOR2x2_ASAP7_75t_R _16101_ (.A(_08066_),
    .B(_00948_),
    .Y(_08067_));
 XOR2x2_ASAP7_75t_R _16102_ (.A(_00852_),
    .B(_00884_),
    .Y(_08068_));
 XOR2x2_ASAP7_75t_R _16103_ (.A(_08067_),
    .B(_08068_),
    .Y(_08069_));
 NAND2x1_ASAP7_75t_R _16104_ (.A(_08005_),
    .B(_08069_),
    .Y(_08070_));
 OA21x2_ASAP7_75t_R _16105_ (.A1(_08005_),
    .A2(key[22]),
    .B(_08070_),
    .Y(_08071_));
 XOR2x2_ASAP7_75t_R _16108_ (.A(_00443_),
    .B(_00917_),
    .Y(_08073_));
 XOR2x2_ASAP7_75t_R _16109_ (.A(_08073_),
    .B(_00949_),
    .Y(_08074_));
 XOR2x2_ASAP7_75t_R _16110_ (.A(_00853_),
    .B(_00885_),
    .Y(_08075_));
 XOR2x2_ASAP7_75t_R _16111_ (.A(_08074_),
    .B(_08075_),
    .Y(_08076_));
 NAND2x1_ASAP7_75t_R _16112_ (.A(_08005_),
    .B(_08076_),
    .Y(_08077_));
 OA21x2_ASAP7_75t_R _16113_ (.A1(_08005_),
    .A2(key[23]),
    .B(_08077_),
    .Y(_08078_));
 INVx4_ASAP7_75t_SL _16115_ (.A(_08052_),
    .Y(_00972_));
 INVx3_ASAP7_75t_SL _16117_ (.A(_08045_),
    .Y(_00973_));
 INVx1_ASAP7_75t_R _16118_ (.A(_00978_),
    .Y(_08079_));
 NAND2x2_ASAP7_75t_SL _16120_ (.A(_08079_),
    .B(_08063_),
    .Y(_08081_));
 INVx1_ASAP7_75t_R _16122_ (.A(_00979_),
    .Y(_08083_));
 NOR2x1_ASAP7_75t_R _16123_ (.A(_08083_),
    .B(_08063_),
    .Y(_08084_));
 NOR2x1_ASAP7_75t_SL _16124_ (.A(_08036_),
    .B(_08084_),
    .Y(_08085_));
 NAND2x1_ASAP7_75t_SL _16125_ (.A(_08081_),
    .B(_08085_),
    .Y(_08086_));
 NAND2x1_ASAP7_75t_SL _16127_ (.A(_08045_),
    .B(_08063_),
    .Y(_08088_));
 NAND2x1_ASAP7_75t_SL _16128_ (.A(_08036_),
    .B(_08088_),
    .Y(_08089_));
 AND2x2_ASAP7_75t_SL _16130_ (.A(_08089_),
    .B(_08018_),
    .Y(_08091_));
 INVx1_ASAP7_75t_SL _16131_ (.A(_08071_),
    .Y(_08092_));
 AOI21x1_ASAP7_75t_SL _16132_ (.A1(_08086_),
    .A2(_08091_),
    .B(_08092_),
    .Y(_08093_));
 INVx1_ASAP7_75t_SL _16133_ (.A(_00975_),
    .Y(_08094_));
 NOR2x1_ASAP7_75t_SL _16134_ (.A(_08094_),
    .B(_08063_),
    .Y(_08095_));
 NOR2x1_ASAP7_75t_SL _16135_ (.A(_08036_),
    .B(_08095_),
    .Y(_08096_));
 INVx1_ASAP7_75t_SL _16136_ (.A(_08096_),
    .Y(_08097_));
 NAND2x2_ASAP7_75t_SL _16137_ (.A(_00976_),
    .B(_08063_),
    .Y(_08098_));
 INVx1_ASAP7_75t_SL _16138_ (.A(_08098_),
    .Y(_08099_));
 NAND2x1_ASAP7_75t_SL _16139_ (.A(_08045_),
    .B(_00989_),
    .Y(_08100_));
 AND2x2_ASAP7_75t_SL _16140_ (.A(_08081_),
    .B(_08036_),
    .Y(_08101_));
 AOI21x1_ASAP7_75t_SL _16142_ (.A1(_08100_),
    .A2(_08101_),
    .B(_08018_),
    .Y(_08103_));
 OAI21x1_ASAP7_75t_SL _16143_ (.A1(_08097_),
    .A2(_08099_),
    .B(_08103_),
    .Y(_08104_));
 INVx1_ASAP7_75t_SL _16144_ (.A(_08028_),
    .Y(_08105_));
 AOI21x1_ASAP7_75t_SL _16146_ (.A1(_08093_),
    .A2(_08104_),
    .B(_08105_),
    .Y(_08107_));
 INVx1_ASAP7_75t_R _16147_ (.A(_00974_),
    .Y(_08108_));
 NAND2x1_ASAP7_75t_SL _16149_ (.A(_08108_),
    .B(_08063_),
    .Y(_08110_));
 INVx1_ASAP7_75t_SL _16150_ (.A(_08110_),
    .Y(_08111_));
 AO21x1_ASAP7_75t_SL _16152_ (.A1(_00989_),
    .A2(_00975_),
    .B(_08037_),
    .Y(_08113_));
 AND2x2_ASAP7_75t_SL _16153_ (.A(_08063_),
    .B(_00983_),
    .Y(_08114_));
 INVx1_ASAP7_75t_R _16154_ (.A(_08114_),
    .Y(_08115_));
 INVx1_ASAP7_75t_SL _16155_ (.A(_00981_),
    .Y(_08116_));
 NOR2x1_ASAP7_75t_SL _16156_ (.A(_08116_),
    .B(_08063_),
    .Y(_08117_));
 INVx1_ASAP7_75t_SL _16157_ (.A(_08117_),
    .Y(_08118_));
 AO21x1_ASAP7_75t_SL _16159_ (.A1(_08115_),
    .A2(_08118_),
    .B(_08036_),
    .Y(_08120_));
 OAI21x1_ASAP7_75t_SL _16160_ (.A1(_08111_),
    .A2(_08113_),
    .B(_08120_),
    .Y(_08121_));
 NAND2x1_ASAP7_75t_SL _16161_ (.A(_08045_),
    .B(_08052_),
    .Y(_08122_));
 NOR2x2_ASAP7_75t_SL _16162_ (.A(_08045_),
    .B(_08063_),
    .Y(_08123_));
 NOR2x1_ASAP7_75t_SL _16163_ (.A(_08037_),
    .B(_08123_),
    .Y(_08124_));
 NAND2x1_ASAP7_75t_SL _16164_ (.A(_08122_),
    .B(_08124_),
    .Y(_08125_));
 INVx1_ASAP7_75t_SL _16166_ (.A(_08123_),
    .Y(_08127_));
 NAND2x1_ASAP7_75t_SL _16167_ (.A(_08122_),
    .B(_08127_),
    .Y(_08128_));
 AOI21x1_ASAP7_75t_SL _16168_ (.A1(_08037_),
    .A2(_08128_),
    .B(_08018_),
    .Y(_08129_));
 AOI21x1_ASAP7_75t_SL _16169_ (.A1(_08125_),
    .A2(_08129_),
    .B(_08071_),
    .Y(_08130_));
 OAI21x1_ASAP7_75t_SL _16170_ (.A1(_08020_),
    .A2(_08121_),
    .B(_08130_),
    .Y(_08131_));
 AOI21x1_ASAP7_75t_SL _16171_ (.A1(_08107_),
    .A2(_08131_),
    .B(_08078_),
    .Y(_08132_));
 NOR2x1_ASAP7_75t_SL _16172_ (.A(_00975_),
    .B(_08063_),
    .Y(_08133_));
 INVx1_ASAP7_75t_R _16173_ (.A(_08133_),
    .Y(_08134_));
 AO21x1_ASAP7_75t_SL _16175_ (.A1(_08115_),
    .A2(_08134_),
    .B(_08036_),
    .Y(_08136_));
 AND2x2_ASAP7_75t_SL _16176_ (.A(_08063_),
    .B(_00981_),
    .Y(_08137_));
 INVx1_ASAP7_75t_SL _16177_ (.A(_08137_),
    .Y(_08138_));
 OA21x2_ASAP7_75t_SL _16178_ (.A1(_08062_),
    .A2(_08054_),
    .B(_00983_),
    .Y(_08139_));
 INVx1_ASAP7_75t_SL _16179_ (.A(_08139_),
    .Y(_08140_));
 AO21x1_ASAP7_75t_SL _16182_ (.A1(_08138_),
    .A2(_08140_),
    .B(_08037_),
    .Y(_08143_));
 AOI21x1_ASAP7_75t_SL _16185_ (.A1(_08136_),
    .A2(_08143_),
    .B(_08020_),
    .Y(_08146_));
 NAND2x1_ASAP7_75t_SL _16186_ (.A(_08036_),
    .B(_08095_),
    .Y(_08147_));
 NAND2x1_ASAP7_75t_SL _16187_ (.A(_00975_),
    .B(_08063_),
    .Y(_08148_));
 NAND2x1_ASAP7_75t_R _16188_ (.A(_08037_),
    .B(_08148_),
    .Y(_08149_));
 AND2x2_ASAP7_75t_SL _16189_ (.A(_08147_),
    .B(_08149_),
    .Y(_08150_));
 NAND2x2_ASAP7_75t_SL _16190_ (.A(_08052_),
    .B(_08063_),
    .Y(_08151_));
 NOR2x1_ASAP7_75t_SL _16191_ (.A(_08037_),
    .B(_08151_),
    .Y(_08152_));
 NOR2x1_ASAP7_75t_SL _16192_ (.A(_08018_),
    .B(_08152_),
    .Y(_08153_));
 AO21x1_ASAP7_75t_SL _16193_ (.A1(_08150_),
    .A2(_08153_),
    .B(_08071_),
    .Y(_08154_));
 NOR2x1_ASAP7_75t_SL _16194_ (.A(_08146_),
    .B(_08154_),
    .Y(_08155_));
 INVx1_ASAP7_75t_SL _16195_ (.A(_08152_),
    .Y(_08156_));
 NOR2x1_ASAP7_75t_SL _16196_ (.A(_00984_),
    .B(_08063_),
    .Y(_08157_));
 NAND2x1_ASAP7_75t_SL _16197_ (.A(_08036_),
    .B(_08157_),
    .Y(_08158_));
 AND2x2_ASAP7_75t_SL _16198_ (.A(_08156_),
    .B(_08158_),
    .Y(_08159_));
 AND3x1_ASAP7_75t_SL _16199_ (.A(_08037_),
    .B(_00973_),
    .C(_08063_),
    .Y(_08160_));
 NOR2x1_ASAP7_75t_SL _16200_ (.A(_08108_),
    .B(_08063_),
    .Y(_08161_));
 AO21x1_ASAP7_75t_SL _16201_ (.A1(_08161_),
    .A2(_08037_),
    .B(_08020_),
    .Y(_08162_));
 NOR2x1_ASAP7_75t_SL _16202_ (.A(_08160_),
    .B(_08162_),
    .Y(_08163_));
 NAND2x1_ASAP7_75t_SL _16203_ (.A(_08159_),
    .B(_08163_),
    .Y(_08164_));
 NOR2x1_ASAP7_75t_SL _16204_ (.A(_08063_),
    .B(_00972_),
    .Y(_08165_));
 NOR2x1_ASAP7_75t_SL _16205_ (.A(_08037_),
    .B(_08165_),
    .Y(_08166_));
 INVx1_ASAP7_75t_SL _16206_ (.A(_00976_),
    .Y(_08167_));
 NOR2x1_ASAP7_75t_SL _16207_ (.A(_08167_),
    .B(_08063_),
    .Y(_08168_));
 NAND2x1_ASAP7_75t_SL _16208_ (.A(_08037_),
    .B(_08088_),
    .Y(_08169_));
 OAI21x1_ASAP7_75t_SL _16209_ (.A1(_08168_),
    .A2(_08169_),
    .B(_08020_),
    .Y(_08170_));
 AO21x1_ASAP7_75t_SL _16210_ (.A1(_08166_),
    .A2(_08081_),
    .B(_08170_),
    .Y(_08171_));
 AOI21x1_ASAP7_75t_SL _16211_ (.A1(_08164_),
    .A2(_08171_),
    .B(_08092_),
    .Y(_08172_));
 OAI21x1_ASAP7_75t_SL _16213_ (.A1(_08155_),
    .A2(_08172_),
    .B(_08105_),
    .Y(_08174_));
 NAND2x1_ASAP7_75t_SL _16214_ (.A(_08132_),
    .B(_08174_),
    .Y(_08175_));
 INVx1_ASAP7_75t_SL _16215_ (.A(_00991_),
    .Y(_08176_));
 NAND2x1_ASAP7_75t_SL _16217_ (.A(_08094_),
    .B(_08063_),
    .Y(_08178_));
 NAND2x1_ASAP7_75t_SL _16219_ (.A(_08036_),
    .B(_08178_),
    .Y(_08180_));
 OAI21x1_ASAP7_75t_SL _16220_ (.A1(_08176_),
    .A2(_08036_),
    .B(_08180_),
    .Y(_08181_));
 AOI21x1_ASAP7_75t_SL _16221_ (.A1(_08020_),
    .A2(_08181_),
    .B(_08028_),
    .Y(_08182_));
 NOR2x1_ASAP7_75t_SL _16222_ (.A(_08079_),
    .B(_08063_),
    .Y(_08183_));
 INVx1_ASAP7_75t_SL _16223_ (.A(_08183_),
    .Y(_08184_));
 AO21x1_ASAP7_75t_SL _16224_ (.A1(_08184_),
    .A2(_08088_),
    .B(_08037_),
    .Y(_08185_));
 AO21x1_ASAP7_75t_SL _16225_ (.A1(_08139_),
    .A2(_08037_),
    .B(_08020_),
    .Y(_08186_));
 NOR2x1_ASAP7_75t_SL _16226_ (.A(_08160_),
    .B(_08186_),
    .Y(_08187_));
 NAND2x1_ASAP7_75t_SL _16227_ (.A(_08185_),
    .B(_08187_),
    .Y(_08188_));
 NAND2x1_ASAP7_75t_SL _16228_ (.A(_08182_),
    .B(_08188_),
    .Y(_08189_));
 NAND2x1_ASAP7_75t_SL _16230_ (.A(_08037_),
    .B(_08157_),
    .Y(_08191_));
 OAI21x1_ASAP7_75t_SL _16232_ (.A1(_08183_),
    .A2(_08137_),
    .B(_08036_),
    .Y(_08193_));
 AOI21x1_ASAP7_75t_SL _16234_ (.A1(_08191_),
    .A2(_08193_),
    .B(_08018_),
    .Y(_08195_));
 NAND2x2_ASAP7_75t_SL _16235_ (.A(_00982_),
    .B(_08063_),
    .Y(_08196_));
 AND2x2_ASAP7_75t_SL _16236_ (.A(_08196_),
    .B(_08037_),
    .Y(_08197_));
 OAI21x1_ASAP7_75t_SL _16237_ (.A1(_00978_),
    .A2(_08063_),
    .B(_08197_),
    .Y(_08198_));
 AOI21x1_ASAP7_75t_SL _16239_ (.A1(_08158_),
    .A2(_08198_),
    .B(_08020_),
    .Y(_08200_));
 OAI21x1_ASAP7_75t_SL _16241_ (.A1(_08195_),
    .A2(_08200_),
    .B(_08028_),
    .Y(_08202_));
 AOI21x1_ASAP7_75t_SL _16242_ (.A1(_08189_),
    .A2(_08202_),
    .B(_08071_),
    .Y(_08203_));
 NAND2x2_ASAP7_75t_SL _16243_ (.A(_08083_),
    .B(_08063_),
    .Y(_08204_));
 INVx1_ASAP7_75t_SL _16244_ (.A(_08204_),
    .Y(_08205_));
 NAND2x1_ASAP7_75t_SL _16245_ (.A(_08036_),
    .B(_08205_),
    .Y(_08206_));
 INVx1_ASAP7_75t_R _16246_ (.A(_08161_),
    .Y(_08207_));
 NAND2x1_ASAP7_75t_SL _16247_ (.A(_08063_),
    .B(_00973_),
    .Y(_08208_));
 AO21x1_ASAP7_75t_SL _16249_ (.A1(_08207_),
    .A2(_08208_),
    .B(_08036_),
    .Y(_08210_));
 AOI21x1_ASAP7_75t_SL _16250_ (.A1(_08206_),
    .A2(_08210_),
    .B(_08020_),
    .Y(_08211_));
 NOR2x1_ASAP7_75t_SL _16251_ (.A(_00982_),
    .B(_08063_),
    .Y(_08212_));
 INVx1_ASAP7_75t_R _16252_ (.A(_08212_),
    .Y(_08213_));
 AO21x1_ASAP7_75t_SL _16253_ (.A1(_08213_),
    .A2(_08204_),
    .B(_08037_),
    .Y(_08214_));
 AOI21x1_ASAP7_75t_SL _16255_ (.A1(_08097_),
    .A2(_08214_),
    .B(_08018_),
    .Y(_08216_));
 OAI21x1_ASAP7_75t_SL _16256_ (.A1(_08211_),
    .A2(_08216_),
    .B(_08105_),
    .Y(_08217_));
 INVx1_ASAP7_75t_SL _16257_ (.A(_08085_),
    .Y(_08218_));
 OAI21x1_ASAP7_75t_SL _16258_ (.A1(_08157_),
    .A2(_08114_),
    .B(_08036_),
    .Y(_08219_));
 AOI21x1_ASAP7_75t_SL _16259_ (.A1(_08218_),
    .A2(_08219_),
    .B(_08018_),
    .Y(_08220_));
 NOR2x1_ASAP7_75t_SL _16260_ (.A(_08036_),
    .B(_08123_),
    .Y(_08221_));
 AND2x2_ASAP7_75t_SL _16261_ (.A(_08221_),
    .B(_08138_),
    .Y(_08222_));
 AO21x1_ASAP7_75t_SL _16262_ (.A1(_08166_),
    .A2(_08148_),
    .B(_08020_),
    .Y(_08223_));
 NOR2x1_ASAP7_75t_SL _16263_ (.A(_08222_),
    .B(_08223_),
    .Y(_08224_));
 OAI21x1_ASAP7_75t_SL _16264_ (.A1(_08220_),
    .A2(_08224_),
    .B(_08028_),
    .Y(_08225_));
 AOI21x1_ASAP7_75t_SL _16266_ (.A1(_08217_),
    .A2(_08225_),
    .B(_08092_),
    .Y(_08227_));
 OAI21x1_ASAP7_75t_SL _16267_ (.A1(_08203_),
    .A2(_08227_),
    .B(_08078_),
    .Y(_08228_));
 NAND2x1_ASAP7_75t_SL _16268_ (.A(_08175_),
    .B(_08228_),
    .Y(_00000_));
 NAND2x1_ASAP7_75t_SL _16269_ (.A(_08151_),
    .B(_08085_),
    .Y(_08229_));
 NAND2x2_ASAP7_75t_SL _16270_ (.A(_08063_),
    .B(_00972_),
    .Y(_08230_));
 NAND2x1_ASAP7_75t_R _16271_ (.A(_08230_),
    .B(_08124_),
    .Y(_08231_));
 AND3x1_ASAP7_75t_SL _16273_ (.A(_08229_),
    .B(_08231_),
    .C(_08105_),
    .Y(_08233_));
 AO21x1_ASAP7_75t_SL _16274_ (.A1(_08115_),
    .A2(_08127_),
    .B(_08037_),
    .Y(_08234_));
 AND2x2_ASAP7_75t_SL _16275_ (.A(_08063_),
    .B(_00978_),
    .Y(_08235_));
 INVx2_ASAP7_75t_SL _16276_ (.A(_08235_),
    .Y(_08236_));
 AO21x1_ASAP7_75t_SL _16277_ (.A1(_08236_),
    .A2(_08207_),
    .B(_08036_),
    .Y(_08237_));
 NAND2x1_ASAP7_75t_SL _16278_ (.A(_08234_),
    .B(_08237_),
    .Y(_08238_));
 OAI21x1_ASAP7_75t_SL _16279_ (.A1(_08105_),
    .A2(_08238_),
    .B(_08020_),
    .Y(_08239_));
 INVx1_ASAP7_75t_SL _16280_ (.A(_00992_),
    .Y(_08240_));
 OR3x1_ASAP7_75t_SL _16282_ (.A(_08028_),
    .B(_08240_),
    .C(_08036_),
    .Y(_08242_));
 OAI21x1_ASAP7_75t_SL _16283_ (.A1(_08161_),
    .A2(_08137_),
    .B(_08036_),
    .Y(_08243_));
 AO21x1_ASAP7_75t_SL _16284_ (.A1(_08242_),
    .A2(_08243_),
    .B(_08020_),
    .Y(_08244_));
 OAI21x1_ASAP7_75t_SL _16285_ (.A1(_08233_),
    .A2(_08239_),
    .B(_08244_),
    .Y(_08245_));
 NOR2x1_ASAP7_75t_SL _16286_ (.A(_08071_),
    .B(_08245_),
    .Y(_08246_));
 AO21x1_ASAP7_75t_SL _16287_ (.A1(_08207_),
    .A2(_08208_),
    .B(_08037_),
    .Y(_08247_));
 AO21x1_ASAP7_75t_SL _16288_ (.A1(_08247_),
    .A2(_08097_),
    .B(_08020_),
    .Y(_08248_));
 NAND2x1_ASAP7_75t_SL _16289_ (.A(_00984_),
    .B(_08063_),
    .Y(_08249_));
 NOR2x1_ASAP7_75t_SL _16290_ (.A(_08037_),
    .B(_08168_),
    .Y(_08250_));
 NAND2x1_ASAP7_75t_R _16291_ (.A(_08037_),
    .B(_08110_),
    .Y(_08251_));
 NOR2x1_ASAP7_75t_SL _16292_ (.A(_08133_),
    .B(_08251_),
    .Y(_08252_));
 AO21x1_ASAP7_75t_SL _16293_ (.A1(_08249_),
    .A2(_08250_),
    .B(_08252_),
    .Y(_08253_));
 NAND2x1_ASAP7_75t_SL _16294_ (.A(_08020_),
    .B(_08253_),
    .Y(_08254_));
 AOI21x1_ASAP7_75t_SL _16295_ (.A1(_08248_),
    .A2(_08254_),
    .B(_08028_),
    .Y(_08255_));
 OAI21x1_ASAP7_75t_SL _16296_ (.A1(_08036_),
    .A2(_08140_),
    .B(_08158_),
    .Y(_08256_));
 OA21x2_ASAP7_75t_SL _16297_ (.A1(_08208_),
    .A2(_08037_),
    .B(_08020_),
    .Y(_08257_));
 OAI21x1_ASAP7_75t_SL _16298_ (.A1(_08036_),
    .A2(_08178_),
    .B(_08257_),
    .Y(_08258_));
 OAI21x1_ASAP7_75t_SL _16299_ (.A1(_08256_),
    .A2(_08258_),
    .B(_08028_),
    .Y(_08259_));
 AO21x1_ASAP7_75t_SL _16300_ (.A1(_08115_),
    .A2(_08100_),
    .B(_08037_),
    .Y(_08260_));
 AND3x1_ASAP7_75t_SL _16301_ (.A(_08260_),
    .B(_08018_),
    .C(_08229_),
    .Y(_08261_));
 OAI21x1_ASAP7_75t_SL _16302_ (.A1(_08259_),
    .A2(_08261_),
    .B(_08071_),
    .Y(_08262_));
 INVx1_ASAP7_75t_SL _16303_ (.A(_08078_),
    .Y(_08263_));
 OAI21x1_ASAP7_75t_SL _16305_ (.A1(_08255_),
    .A2(_08262_),
    .B(_08263_),
    .Y(_08265_));
 INVx2_ASAP7_75t_SL _16306_ (.A(_08165_),
    .Y(_08266_));
 AND2x2_ASAP7_75t_SL _16307_ (.A(_08098_),
    .B(_08037_),
    .Y(_08267_));
 AOI21x1_ASAP7_75t_SL _16308_ (.A1(_08266_),
    .A2(_08267_),
    .B(_08018_),
    .Y(_08268_));
 OAI21x1_ASAP7_75t_SL _16309_ (.A1(_08037_),
    .A2(_08207_),
    .B(_08268_),
    .Y(_08269_));
 NAND2x1_ASAP7_75t_R _16310_ (.A(_08083_),
    .B(_00989_),
    .Y(_08270_));
 OAI21x1_ASAP7_75t_SL _16312_ (.A1(_08037_),
    .A2(_08270_),
    .B(_08018_),
    .Y(_08272_));
 OA21x2_ASAP7_75t_SL _16313_ (.A1(_08252_),
    .A2(_08272_),
    .B(_08028_),
    .Y(_08273_));
 AO21x1_ASAP7_75t_SL _16314_ (.A1(_08269_),
    .A2(_08273_),
    .B(_08092_),
    .Y(_08274_));
 AND3x1_ASAP7_75t_SL _16315_ (.A(_08100_),
    .B(_08036_),
    .C(_08178_),
    .Y(_08275_));
 NAND2x1_ASAP7_75t_R _16316_ (.A(_08052_),
    .B(_00973_),
    .Y(_08276_));
 AND3x1_ASAP7_75t_SL _16317_ (.A(_08088_),
    .B(_08037_),
    .C(_08276_),
    .Y(_08277_));
 OA21x2_ASAP7_75t_SL _16318_ (.A1(_08275_),
    .A2(_08277_),
    .B(_08018_),
    .Y(_08278_));
 AND3x1_ASAP7_75t_SL _16319_ (.A(_08140_),
    .B(_08036_),
    .C(_08208_),
    .Y(_08279_));
 AO21x1_ASAP7_75t_SL _16320_ (.A1(_08096_),
    .A2(_08204_),
    .B(_08018_),
    .Y(_08280_));
 NOR2x1_ASAP7_75t_SL _16321_ (.A(_08279_),
    .B(_08280_),
    .Y(_08281_));
 OA21x2_ASAP7_75t_SL _16322_ (.A1(_08278_),
    .A2(_08281_),
    .B(_08105_),
    .Y(_08282_));
 NAND2x1_ASAP7_75t_SL _16323_ (.A(_08037_),
    .B(_08235_),
    .Y(_08283_));
 AO21x1_ASAP7_75t_SL _16324_ (.A1(_08230_),
    .A2(_08276_),
    .B(_08037_),
    .Y(_08284_));
 AOI21x1_ASAP7_75t_SL _16325_ (.A1(_08283_),
    .A2(_08284_),
    .B(_08020_),
    .Y(_08285_));
 AO21x1_ASAP7_75t_SL _16326_ (.A1(_08270_),
    .A2(_08088_),
    .B(_08037_),
    .Y(_08286_));
 AO21x1_ASAP7_75t_SL _16327_ (.A1(_08134_),
    .A2(_08208_),
    .B(_08036_),
    .Y(_08287_));
 AOI21x1_ASAP7_75t_SL _16328_ (.A1(_08286_),
    .A2(_08287_),
    .B(_08018_),
    .Y(_08288_));
 OAI21x1_ASAP7_75t_SL _16329_ (.A1(_08285_),
    .A2(_08288_),
    .B(_08028_),
    .Y(_08289_));
 OA21x2_ASAP7_75t_SL _16330_ (.A1(_08204_),
    .A2(_08037_),
    .B(_08020_),
    .Y(_08290_));
 AND2x2_ASAP7_75t_SL _16331_ (.A(_08037_),
    .B(_00986_),
    .Y(_08291_));
 AOI21x1_ASAP7_75t_SL _16332_ (.A1(_08036_),
    .A2(_08165_),
    .B(_08291_),
    .Y(_08292_));
 AOI21x1_ASAP7_75t_SL _16333_ (.A1(_08290_),
    .A2(_08292_),
    .B(_08028_),
    .Y(_08293_));
 AO21x1_ASAP7_75t_SL _16334_ (.A1(_08184_),
    .A2(_08204_),
    .B(_08037_),
    .Y(_08294_));
 OA21x2_ASAP7_75t_SL _16335_ (.A1(_08149_),
    .A2(_08168_),
    .B(_08018_),
    .Y(_08295_));
 NAND2x1_ASAP7_75t_SL _16336_ (.A(_08294_),
    .B(_08295_),
    .Y(_08296_));
 AOI21x1_ASAP7_75t_SL _16337_ (.A1(_08293_),
    .A2(_08296_),
    .B(_08071_),
    .Y(_08297_));
 AOI21x1_ASAP7_75t_SL _16338_ (.A1(_08289_),
    .A2(_08297_),
    .B(_08263_),
    .Y(_08298_));
 OAI21x1_ASAP7_75t_SL _16339_ (.A1(_08274_),
    .A2(_08282_),
    .B(_08298_),
    .Y(_08299_));
 OAI21x1_ASAP7_75t_SL _16340_ (.A1(_08246_),
    .A2(_08265_),
    .B(_08299_),
    .Y(_00001_));
 NAND2x1_ASAP7_75t_SL _16341_ (.A(_08167_),
    .B(_08063_),
    .Y(_08300_));
 AOI21x1_ASAP7_75t_SL _16342_ (.A1(_08300_),
    .A2(_08124_),
    .B(_08018_),
    .Y(_08301_));
 INVx1_ASAP7_75t_R _16343_ (.A(_08151_),
    .Y(_08302_));
 OR3x1_ASAP7_75t_SL _16344_ (.A(_08302_),
    .B(_08036_),
    .C(_08212_),
    .Y(_08303_));
 NAND2x1_ASAP7_75t_SL _16345_ (.A(_08301_),
    .B(_08303_),
    .Y(_08304_));
 AO21x1_ASAP7_75t_SL _16346_ (.A1(_08134_),
    .A2(_08148_),
    .B(_08036_),
    .Y(_08305_));
 NAND3x1_ASAP7_75t_SL _16347_ (.A(_08100_),
    .B(_08036_),
    .C(_08196_),
    .Y(_08306_));
 AO21x1_ASAP7_75t_SL _16348_ (.A1(_08305_),
    .A2(_08306_),
    .B(_08020_),
    .Y(_08307_));
 AOI21x1_ASAP7_75t_SL _16349_ (.A1(_08304_),
    .A2(_08307_),
    .B(_08105_),
    .Y(_08308_));
 NOR2x2_ASAP7_75t_SL _16350_ (.A(_08052_),
    .B(_08063_),
    .Y(_08309_));
 INVx1_ASAP7_75t_R _16351_ (.A(_08309_),
    .Y(_08310_));
 AO21x1_ASAP7_75t_SL _16352_ (.A1(_08310_),
    .A2(_08204_),
    .B(_08036_),
    .Y(_08311_));
 AND3x1_ASAP7_75t_SL _16353_ (.A(_08214_),
    .B(_08311_),
    .C(_08018_),
    .Y(_08312_));
 AND2x2_ASAP7_75t_SL _16355_ (.A(_08300_),
    .B(_08036_),
    .Y(_08314_));
 AOI22x1_ASAP7_75t_SL _16356_ (.A1(_08221_),
    .A2(_08204_),
    .B1(_08314_),
    .B2(_08213_),
    .Y(_08315_));
 OAI21x1_ASAP7_75t_SL _16357_ (.A1(_08018_),
    .A2(_08315_),
    .B(_08105_),
    .Y(_08316_));
 OAI21x1_ASAP7_75t_SL _16358_ (.A1(_08312_),
    .A2(_08316_),
    .B(_08071_),
    .Y(_08317_));
 NOR2x1_ASAP7_75t_SL _16359_ (.A(_08308_),
    .B(_08317_),
    .Y(_08318_));
 NOR2x1_ASAP7_75t_SL _16360_ (.A(_08168_),
    .B(_08251_),
    .Y(_08319_));
 AO21x1_ASAP7_75t_SL _16361_ (.A1(_08081_),
    .A2(_08036_),
    .B(_08020_),
    .Y(_08320_));
 OA21x2_ASAP7_75t_SL _16362_ (.A1(_08319_),
    .A2(_08320_),
    .B(_08028_),
    .Y(_08321_));
 NOR2x1_ASAP7_75t_SL _16363_ (.A(_08037_),
    .B(_08133_),
    .Y(_08322_));
 NAND2x1_ASAP7_75t_SL _16364_ (.A(_08151_),
    .B(_08322_),
    .Y(_08323_));
 INVx1_ASAP7_75t_R _16365_ (.A(_00984_),
    .Y(_08324_));
 NAND2x1_ASAP7_75t_R _16366_ (.A(_08324_),
    .B(_08063_),
    .Y(_08325_));
 NAND2x1_ASAP7_75t_SL _16367_ (.A(_08325_),
    .B(_08221_),
    .Y(_08326_));
 AO21x1_ASAP7_75t_SL _16368_ (.A1(_08323_),
    .A2(_08326_),
    .B(_08018_),
    .Y(_08327_));
 AO21x1_ASAP7_75t_SL _16369_ (.A1(_08321_),
    .A2(_08327_),
    .B(_08071_),
    .Y(_08328_));
 NAND2x1_ASAP7_75t_R _16370_ (.A(_08037_),
    .B(_08204_),
    .Y(_08329_));
 OA21x2_ASAP7_75t_SL _16371_ (.A1(_08329_),
    .A2(_08183_),
    .B(_08018_),
    .Y(_08330_));
 OAI21x1_ASAP7_75t_SL _16372_ (.A1(_08309_),
    .A2(_08180_),
    .B(_08330_),
    .Y(_08331_));
 AO21x1_ASAP7_75t_SL _16373_ (.A1(_08236_),
    .A2(_08266_),
    .B(_08036_),
    .Y(_08332_));
 AO21x1_ASAP7_75t_SL _16374_ (.A1(_08270_),
    .A2(_08300_),
    .B(_08037_),
    .Y(_08333_));
 AO21x1_ASAP7_75t_SL _16375_ (.A1(_08332_),
    .A2(_08333_),
    .B(_08018_),
    .Y(_08334_));
 AOI21x1_ASAP7_75t_SL _16376_ (.A1(_08331_),
    .A2(_08334_),
    .B(_08028_),
    .Y(_08335_));
 OAI21x1_ASAP7_75t_SL _16377_ (.A1(_08328_),
    .A2(_08335_),
    .B(_08263_),
    .Y(_08336_));
 AND3x1_ASAP7_75t_SL _16378_ (.A(_08115_),
    .B(_08036_),
    .C(_08310_),
    .Y(_08337_));
 AND2x2_ASAP7_75t_R _16379_ (.A(_08178_),
    .B(_08037_),
    .Y(_08338_));
 AO21x1_ASAP7_75t_SL _16380_ (.A1(_08338_),
    .A2(_08118_),
    .B(_08018_),
    .Y(_08339_));
 NOR2x1_ASAP7_75t_SL _16381_ (.A(_08337_),
    .B(_08339_),
    .Y(_08340_));
 NAND2x1_ASAP7_75t_SL _16382_ (.A(_00992_),
    .B(_08036_),
    .Y(_08341_));
 AO21x1_ASAP7_75t_SL _16383_ (.A1(_08230_),
    .A2(_08276_),
    .B(_08036_),
    .Y(_08342_));
 AOI21x1_ASAP7_75t_SL _16384_ (.A1(_08341_),
    .A2(_08342_),
    .B(_08020_),
    .Y(_08343_));
 OA21x2_ASAP7_75t_SL _16385_ (.A1(_08340_),
    .A2(_08343_),
    .B(_08105_),
    .Y(_08344_));
 OA21x2_ASAP7_75t_SL _16386_ (.A1(_08063_),
    .A2(_08045_),
    .B(_00988_),
    .Y(_08345_));
 NOR2x1_ASAP7_75t_SL _16387_ (.A(_08036_),
    .B(_08345_),
    .Y(_08346_));
 NOR2x1_ASAP7_75t_SL _16388_ (.A(_08309_),
    .B(_08180_),
    .Y(_08347_));
 OR3x1_ASAP7_75t_SL _16389_ (.A(_08346_),
    .B(_08018_),
    .C(_08347_),
    .Y(_08348_));
 NOR2x1_ASAP7_75t_SL _16390_ (.A(_00978_),
    .B(_08063_),
    .Y(_08349_));
 NAND2x1_ASAP7_75t_R _16391_ (.A(_08176_),
    .B(_08036_),
    .Y(_08350_));
 OA21x2_ASAP7_75t_SL _16392_ (.A1(_08149_),
    .A2(_08349_),
    .B(_08350_),
    .Y(_08351_));
 AOI21x1_ASAP7_75t_SL _16393_ (.A1(_08018_),
    .A2(_08351_),
    .B(_08105_),
    .Y(_08352_));
 AO21x1_ASAP7_75t_SL _16394_ (.A1(_08348_),
    .A2(_08352_),
    .B(_08092_),
    .Y(_08353_));
 OA21x2_ASAP7_75t_SL _16395_ (.A1(_08037_),
    .A2(_00988_),
    .B(_08020_),
    .Y(_08354_));
 AND2x2_ASAP7_75t_SL _16396_ (.A(_08037_),
    .B(_00990_),
    .Y(_08355_));
 OAI21x1_ASAP7_75t_SL _16397_ (.A1(_08355_),
    .A2(_08320_),
    .B(_08105_),
    .Y(_08356_));
 AO21x1_ASAP7_75t_SL _16398_ (.A1(_08332_),
    .A2(_08354_),
    .B(_08356_),
    .Y(_08357_));
 NAND2x1_ASAP7_75t_SL _16399_ (.A(_00979_),
    .B(_08063_),
    .Y(_08358_));
 NAND2x1_ASAP7_75t_SL _16400_ (.A(_08358_),
    .B(_08096_),
    .Y(_08359_));
 NAND2x1_ASAP7_75t_SL _16401_ (.A(_08036_),
    .B(_08139_),
    .Y(_08360_));
 AND2x2_ASAP7_75t_SL _16402_ (.A(_08360_),
    .B(_08018_),
    .Y(_08361_));
 AOI21x1_ASAP7_75t_SL _16403_ (.A1(_08359_),
    .A2(_08361_),
    .B(_08105_),
    .Y(_08362_));
 NAND2x1_ASAP7_75t_SL _16404_ (.A(_08110_),
    .B(_08221_),
    .Y(_08363_));
 NAND3x1_ASAP7_75t_SL _16405_ (.A(_08363_),
    .B(_08020_),
    .C(_08243_),
    .Y(_08364_));
 AOI21x1_ASAP7_75t_SL _16406_ (.A1(_08362_),
    .A2(_08364_),
    .B(_08071_),
    .Y(_08365_));
 AOI21x1_ASAP7_75t_SL _16407_ (.A1(_08357_),
    .A2(_08365_),
    .B(_08263_),
    .Y(_08366_));
 OAI21x1_ASAP7_75t_SL _16408_ (.A1(_08344_),
    .A2(_08353_),
    .B(_08366_),
    .Y(_08367_));
 OAI21x1_ASAP7_75t_SL _16409_ (.A1(_08318_),
    .A2(_08336_),
    .B(_08367_),
    .Y(_00002_));
 AO21x1_ASAP7_75t_SL _16410_ (.A1(_08208_),
    .A2(_08122_),
    .B(_08037_),
    .Y(_08368_));
 NAND2x1_ASAP7_75t_SL _16411_ (.A(_08037_),
    .B(_08081_),
    .Y(_08369_));
 AND2x2_ASAP7_75t_SL _16412_ (.A(_08369_),
    .B(_08018_),
    .Y(_08370_));
 AOI21x1_ASAP7_75t_SL _16413_ (.A1(_08368_),
    .A2(_08370_),
    .B(_08028_),
    .Y(_08371_));
 NAND2x1_ASAP7_75t_SL _16414_ (.A(_08196_),
    .B(_08322_),
    .Y(_08372_));
 NAND2x1_ASAP7_75t_SL _16415_ (.A(_08372_),
    .B(_08268_),
    .Y(_08373_));
 NAND2x1_ASAP7_75t_SL _16416_ (.A(_08371_),
    .B(_08373_),
    .Y(_08374_));
 OAI21x1_ASAP7_75t_SL _16417_ (.A1(_08095_),
    .A2(_08137_),
    .B(_08036_),
    .Y(_08375_));
 NAND3x1_ASAP7_75t_SL _16418_ (.A(_08127_),
    .B(_08037_),
    .C(_08122_),
    .Y(_08376_));
 AOI21x1_ASAP7_75t_SL _16419_ (.A1(_08375_),
    .A2(_08376_),
    .B(_08018_),
    .Y(_08377_));
 OAI21x1_ASAP7_75t_SL _16420_ (.A1(_08117_),
    .A2(_08235_),
    .B(_08037_),
    .Y(_08378_));
 AO21x1_ASAP7_75t_SL _16421_ (.A1(_08207_),
    .A2(_08178_),
    .B(_08037_),
    .Y(_08379_));
 AOI21x1_ASAP7_75t_SL _16422_ (.A1(_08378_),
    .A2(_08379_),
    .B(_08020_),
    .Y(_08380_));
 OAI21x1_ASAP7_75t_SL _16423_ (.A1(_08377_),
    .A2(_08380_),
    .B(_08028_),
    .Y(_08381_));
 AOI21x1_ASAP7_75t_SL _16424_ (.A1(_08374_),
    .A2(_08381_),
    .B(_08092_),
    .Y(_08382_));
 NAND2x1_ASAP7_75t_SL _16425_ (.A(_08167_),
    .B(_00989_),
    .Y(_08383_));
 AO21x1_ASAP7_75t_SL _16426_ (.A1(_08383_),
    .A2(_08204_),
    .B(_08036_),
    .Y(_08384_));
 AOI21x1_ASAP7_75t_SL _16427_ (.A1(_08151_),
    .A2(_08322_),
    .B(_08020_),
    .Y(_08385_));
 AOI21x1_ASAP7_75t_SL _16428_ (.A1(_08384_),
    .A2(_08385_),
    .B(_08105_),
    .Y(_08386_));
 NOR2x1_ASAP7_75t_SL _16429_ (.A(_08139_),
    .B(_08149_),
    .Y(_08387_));
 AND3x1_ASAP7_75t_SL _16430_ (.A(_08118_),
    .B(_08036_),
    .C(_08208_),
    .Y(_08388_));
 OAI21x1_ASAP7_75t_SL _16431_ (.A1(_08387_),
    .A2(_08388_),
    .B(_08020_),
    .Y(_08389_));
 NAND2x1_ASAP7_75t_SL _16432_ (.A(_08386_),
    .B(_08389_),
    .Y(_08390_));
 NAND2x1_ASAP7_75t_SL _16433_ (.A(_08151_),
    .B(_08096_),
    .Y(_08391_));
 AOI21x1_ASAP7_75t_SL _16434_ (.A1(_08391_),
    .A2(_08368_),
    .B(_08020_),
    .Y(_08392_));
 OA21x2_ASAP7_75t_SL _16435_ (.A1(_08345_),
    .A2(_08037_),
    .B(_08149_),
    .Y(_08393_));
 NOR2x1_ASAP7_75t_SL _16436_ (.A(_08018_),
    .B(_08393_),
    .Y(_08394_));
 OAI21x1_ASAP7_75t_SL _16437_ (.A1(_08392_),
    .A2(_08394_),
    .B(_08105_),
    .Y(_08395_));
 AOI21x1_ASAP7_75t_SL _16438_ (.A1(_08390_),
    .A2(_08395_),
    .B(_08071_),
    .Y(_08396_));
 OAI21x1_ASAP7_75t_SL _16439_ (.A1(_08382_),
    .A2(_08396_),
    .B(_08078_),
    .Y(_08397_));
 AOI21x1_ASAP7_75t_SL _16440_ (.A1(_08191_),
    .A2(_08147_),
    .B(_08018_),
    .Y(_08398_));
 NAND2x1_ASAP7_75t_SL _16441_ (.A(_08037_),
    .B(_08212_),
    .Y(_08399_));
 AOI21x1_ASAP7_75t_SL _16442_ (.A1(_08399_),
    .A2(_08306_),
    .B(_08020_),
    .Y(_08400_));
 OAI21x1_ASAP7_75t_SL _16443_ (.A1(_08398_),
    .A2(_08400_),
    .B(_08028_),
    .Y(_08401_));
 NAND2x1_ASAP7_75t_SL _16444_ (.A(_08098_),
    .B(_08221_),
    .Y(_08402_));
 AO21x1_ASAP7_75t_SL _16445_ (.A1(_08134_),
    .A2(_08208_),
    .B(_08037_),
    .Y(_08403_));
 AOI21x1_ASAP7_75t_SL _16446_ (.A1(_08402_),
    .A2(_08403_),
    .B(_08020_),
    .Y(_08404_));
 INVx1_ASAP7_75t_SL _16447_ (.A(_08148_),
    .Y(_08405_));
 OAI21x1_ASAP7_75t_SL _16448_ (.A1(_08157_),
    .A2(_08405_),
    .B(_08037_),
    .Y(_08406_));
 AND2x2_ASAP7_75t_R _16449_ (.A(_08063_),
    .B(_08116_),
    .Y(_08407_));
 NOR2x1_ASAP7_75t_SL _16450_ (.A(_08037_),
    .B(_08407_),
    .Y(_08408_));
 NAND2x1_ASAP7_75t_SL _16451_ (.A(_08310_),
    .B(_08408_),
    .Y(_08409_));
 AOI21x1_ASAP7_75t_SL _16452_ (.A1(_08406_),
    .A2(_08409_),
    .B(_08018_),
    .Y(_08410_));
 OAI21x1_ASAP7_75t_SL _16453_ (.A1(_08404_),
    .A2(_08410_),
    .B(_08105_),
    .Y(_08411_));
 AOI21x1_ASAP7_75t_SL _16454_ (.A1(_08401_),
    .A2(_08411_),
    .B(_08071_),
    .Y(_08412_));
 NAND2x1_ASAP7_75t_SL _16455_ (.A(_08196_),
    .B(_08221_),
    .Y(_08413_));
 AOI21x1_ASAP7_75t_SL _16456_ (.A1(_08243_),
    .A2(_08413_),
    .B(_08020_),
    .Y(_08414_));
 OAI21x1_ASAP7_75t_SL _16457_ (.A1(_08301_),
    .A2(_08414_),
    .B(_08105_),
    .Y(_08415_));
 AOI21x1_ASAP7_75t_SL _16458_ (.A1(_08284_),
    .A2(_08187_),
    .B(_08105_),
    .Y(_08416_));
 NOR2x1_ASAP7_75t_SL _16459_ (.A(_08036_),
    .B(_00989_),
    .Y(_08417_));
 NAND2x1_ASAP7_75t_SL _16460_ (.A(_08045_),
    .B(_08417_),
    .Y(_08418_));
 NAND2x1_ASAP7_75t_SL _16461_ (.A(_08399_),
    .B(_08418_),
    .Y(_08419_));
 INVx2_ASAP7_75t_SL _16462_ (.A(_08419_),
    .Y(_08420_));
 AO21x1_ASAP7_75t_SL _16463_ (.A1(_08134_),
    .A2(_08300_),
    .B(_08037_),
    .Y(_08421_));
 NAND3x1_ASAP7_75t_SL _16464_ (.A(_08420_),
    .B(_08020_),
    .C(_08421_),
    .Y(_08422_));
 NAND2x1_ASAP7_75t_SL _16465_ (.A(_08416_),
    .B(_08422_),
    .Y(_08423_));
 AOI21x1_ASAP7_75t_SL _16466_ (.A1(_08415_),
    .A2(_08423_),
    .B(_08092_),
    .Y(_08424_));
 OAI21x1_ASAP7_75t_SL _16467_ (.A1(_08412_),
    .A2(_08424_),
    .B(_08263_),
    .Y(_08425_));
 NAND2x1_ASAP7_75t_SL _16468_ (.A(_08397_),
    .B(_08425_),
    .Y(_00003_));
 NAND2x1_ASAP7_75t_SL _16469_ (.A(_08018_),
    .B(_08342_),
    .Y(_08426_));
 INVx1_ASAP7_75t_SL _16470_ (.A(_08231_),
    .Y(_08427_));
 OA21x2_ASAP7_75t_SL _16471_ (.A1(_08426_),
    .A2(_08427_),
    .B(_08105_),
    .Y(_08428_));
 OR3x1_ASAP7_75t_SL _16472_ (.A(_08114_),
    .B(_08036_),
    .C(_08309_),
    .Y(_08429_));
 NAND2x1_ASAP7_75t_R _16473_ (.A(_00973_),
    .B(_00972_),
    .Y(_08430_));
 AO21x1_ASAP7_75t_SL _16474_ (.A1(_08266_),
    .A2(_08430_),
    .B(_08037_),
    .Y(_08431_));
 AO21x1_ASAP7_75t_SL _16475_ (.A1(_08429_),
    .A2(_08431_),
    .B(_08018_),
    .Y(_08432_));
 AND2x2_ASAP7_75t_SL _16476_ (.A(_08428_),
    .B(_08432_),
    .Y(_08433_));
 OAI21x1_ASAP7_75t_SL _16477_ (.A1(_00993_),
    .A2(_08036_),
    .B(_08018_),
    .Y(_08434_));
 AO221x1_ASAP7_75t_SL _16478_ (.A1(_00973_),
    .A2(_00989_),
    .B1(_08036_),
    .B2(_08114_),
    .C(_08434_),
    .Y(_08435_));
 AO21x1_ASAP7_75t_SL _16479_ (.A1(_00989_),
    .A2(_08324_),
    .B(_08018_),
    .Y(_08436_));
 OA21x2_ASAP7_75t_SL _16480_ (.A1(_08197_),
    .A2(_08436_),
    .B(_08028_),
    .Y(_08437_));
 AO21x1_ASAP7_75t_SL _16481_ (.A1(_08435_),
    .A2(_08437_),
    .B(_08263_),
    .Y(_08438_));
 NAND2x1_ASAP7_75t_SL _16482_ (.A(_08036_),
    .B(_08249_),
    .Y(_08439_));
 AND3x1_ASAP7_75t_SL _16483_ (.A(_08251_),
    .B(_08439_),
    .C(_08020_),
    .Y(_08440_));
 NOR2x1_ASAP7_75t_SL _16484_ (.A(_08105_),
    .B(_08440_),
    .Y(_08441_));
 INVx1_ASAP7_75t_R _16485_ (.A(_08178_),
    .Y(_08442_));
 AO21x1_ASAP7_75t_R _16486_ (.A1(_00989_),
    .A2(_00979_),
    .B(_08037_),
    .Y(_08443_));
 OAI21x1_ASAP7_75t_SL _16487_ (.A1(_08442_),
    .A2(_08443_),
    .B(_08163_),
    .Y(_08444_));
 NAND2x1_ASAP7_75t_SL _16488_ (.A(_08441_),
    .B(_08444_),
    .Y(_08445_));
 NOR2x1_ASAP7_75t_R _16489_ (.A(_08020_),
    .B(_08417_),
    .Y(_08446_));
 NAND2x1_ASAP7_75t_SL _16490_ (.A(_08098_),
    .B(_08124_),
    .Y(_08447_));
 AOI21x1_ASAP7_75t_SL _16491_ (.A1(_08446_),
    .A2(_08447_),
    .B(_08028_),
    .Y(_08448_));
 NAND3x1_ASAP7_75t_SL _16492_ (.A(_08153_),
    .B(_08229_),
    .C(_08360_),
    .Y(_08449_));
 AOI21x1_ASAP7_75t_SL _16493_ (.A1(_08448_),
    .A2(_08449_),
    .B(_08078_),
    .Y(_08450_));
 AOI21x1_ASAP7_75t_SL _16494_ (.A1(_08445_),
    .A2(_08450_),
    .B(_08092_),
    .Y(_08451_));
 OAI21x1_ASAP7_75t_SL _16495_ (.A1(_08433_),
    .A2(_08438_),
    .B(_08451_),
    .Y(_08452_));
 NAND2x1_ASAP7_75t_SL _16496_ (.A(_08148_),
    .B(_08250_),
    .Y(_08453_));
 AOI21x1_ASAP7_75t_SL _16497_ (.A1(_08453_),
    .A2(_08198_),
    .B(_08020_),
    .Y(_08454_));
 AO21x1_ASAP7_75t_SL _16498_ (.A1(_08213_),
    .A2(_08178_),
    .B(_08036_),
    .Y(_08455_));
 AOI21x1_ASAP7_75t_SL _16499_ (.A1(_08214_),
    .A2(_08455_),
    .B(_08018_),
    .Y(_08456_));
 OA21x2_ASAP7_75t_SL _16500_ (.A1(_08454_),
    .A2(_08456_),
    .B(_08028_),
    .Y(_08457_));
 NOR2x1_ASAP7_75t_SL _16501_ (.A(_08036_),
    .B(_08349_),
    .Y(_08458_));
 NAND2x1_ASAP7_75t_SL _16502_ (.A(_08151_),
    .B(_08458_),
    .Y(_08459_));
 AND3x1_ASAP7_75t_SL _16503_ (.A(_08333_),
    .B(_08020_),
    .C(_08459_),
    .Y(_08460_));
 AOI21x1_ASAP7_75t_SL _16504_ (.A1(_00972_),
    .A2(_08417_),
    .B(_08186_),
    .Y(_08461_));
 AO21x1_ASAP7_75t_SL _16505_ (.A1(_08461_),
    .A2(_08294_),
    .B(_08028_),
    .Y(_08462_));
 OAI21x1_ASAP7_75t_SL _16506_ (.A1(_08460_),
    .A2(_08462_),
    .B(_08078_),
    .Y(_08463_));
 AOI21x1_ASAP7_75t_SL _16507_ (.A1(_08036_),
    .A2(_08183_),
    .B(_08018_),
    .Y(_08464_));
 NAND2x1_ASAP7_75t_SL _16508_ (.A(_08266_),
    .B(_08197_),
    .Y(_08465_));
 NAND2x1_ASAP7_75t_SL _16509_ (.A(_08464_),
    .B(_08465_),
    .Y(_08466_));
 AO21x1_ASAP7_75t_SL _16510_ (.A1(_08036_),
    .A2(_00974_),
    .B(_08020_),
    .Y(_08467_));
 OA21x2_ASAP7_75t_SL _16511_ (.A1(_08338_),
    .A2(_08467_),
    .B(_08028_),
    .Y(_08468_));
 AOI21x1_ASAP7_75t_SL _16512_ (.A1(_08466_),
    .A2(_08468_),
    .B(_08078_),
    .Y(_08469_));
 AO21x1_ASAP7_75t_SL _16513_ (.A1(_08127_),
    .A2(_08122_),
    .B(_08036_),
    .Y(_08470_));
 AOI21x1_ASAP7_75t_SL _16514_ (.A1(_08219_),
    .A2(_08470_),
    .B(_08020_),
    .Y(_08471_));
 AOI21x1_ASAP7_75t_SL _16515_ (.A1(_08413_),
    .A2(_08431_),
    .B(_08018_),
    .Y(_08472_));
 OAI21x1_ASAP7_75t_SL _16516_ (.A1(_08471_),
    .A2(_08472_),
    .B(_08105_),
    .Y(_08473_));
 AOI21x1_ASAP7_75t_SL _16517_ (.A1(_08469_),
    .A2(_08473_),
    .B(_08071_),
    .Y(_08474_));
 OAI21x1_ASAP7_75t_SL _16518_ (.A1(_08457_),
    .A2(_08463_),
    .B(_08474_),
    .Y(_08475_));
 NAND2x1_ASAP7_75t_SL _16519_ (.A(_08452_),
    .B(_08475_),
    .Y(_00004_));
 INVx1_ASAP7_75t_SL _16520_ (.A(_08267_),
    .Y(_08476_));
 AOI21x1_ASAP7_75t_SL _16521_ (.A1(_08476_),
    .A2(_08290_),
    .B(_08105_),
    .Y(_08477_));
 NOR2x1_ASAP7_75t_SL _16522_ (.A(_08020_),
    .B(_08221_),
    .Y(_08478_));
 AO21x1_ASAP7_75t_SL _16523_ (.A1(_08236_),
    .A2(_08207_),
    .B(_08037_),
    .Y(_08479_));
 NAND2x1_ASAP7_75t_SL _16524_ (.A(_08478_),
    .B(_08479_),
    .Y(_08480_));
 AOI21x1_ASAP7_75t_SL _16525_ (.A1(_08477_),
    .A2(_08480_),
    .B(_08071_),
    .Y(_08481_));
 OA21x2_ASAP7_75t_SL _16526_ (.A1(_08097_),
    .A2(_08407_),
    .B(_08020_),
    .Y(_08482_));
 NAND2x1_ASAP7_75t_SL _16527_ (.A(_08098_),
    .B(_08322_),
    .Y(_08483_));
 AO21x1_ASAP7_75t_SL _16528_ (.A1(_08108_),
    .A2(_00989_),
    .B(_08037_),
    .Y(_08484_));
 OA21x2_ASAP7_75t_SL _16529_ (.A1(_08036_),
    .A2(_08116_),
    .B(_08018_),
    .Y(_08485_));
 AO21x1_ASAP7_75t_SL _16530_ (.A1(_08484_),
    .A2(_08485_),
    .B(_08028_),
    .Y(_08486_));
 AO21x1_ASAP7_75t_SL _16531_ (.A1(_08482_),
    .A2(_08483_),
    .B(_08486_),
    .Y(_08487_));
 AOI21x1_ASAP7_75t_SL _16532_ (.A1(_08481_),
    .A2(_08487_),
    .B(_08078_),
    .Y(_08488_));
 NAND2x1_ASAP7_75t_SL _16533_ (.A(_08196_),
    .B(_08166_),
    .Y(_08489_));
 OA211x2_ASAP7_75t_SL _16534_ (.A1(_08095_),
    .A2(_08369_),
    .B(_08489_),
    .C(_08020_),
    .Y(_08490_));
 OA21x2_ASAP7_75t_SL _16535_ (.A1(_08036_),
    .A2(_08045_),
    .B(_08125_),
    .Y(_08491_));
 AO21x1_ASAP7_75t_SL _16536_ (.A1(_08491_),
    .A2(_08018_),
    .B(_08105_),
    .Y(_08492_));
 AO21x1_ASAP7_75t_SL _16537_ (.A1(_08127_),
    .A2(_08204_),
    .B(_08037_),
    .Y(_08493_));
 NAND2x1_ASAP7_75t_SL _16538_ (.A(_08493_),
    .B(_08163_),
    .Y(_08494_));
 NOR2x1_ASAP7_75t_SL _16539_ (.A(_08099_),
    .B(_08484_),
    .Y(_08495_));
 AO21x1_ASAP7_75t_SL _16540_ (.A1(_08137_),
    .A2(_08037_),
    .B(_08018_),
    .Y(_08496_));
 OA21x2_ASAP7_75t_SL _16541_ (.A1(_08495_),
    .A2(_08496_),
    .B(_08105_),
    .Y(_08497_));
 AOI21x1_ASAP7_75t_SL _16542_ (.A1(_08494_),
    .A2(_08497_),
    .B(_08092_),
    .Y(_08498_));
 OAI21x1_ASAP7_75t_SL _16543_ (.A1(_08490_),
    .A2(_08492_),
    .B(_08498_),
    .Y(_08499_));
 NAND2x1_ASAP7_75t_SL _16544_ (.A(_08488_),
    .B(_08499_),
    .Y(_08500_));
 NOR2x1_ASAP7_75t_SL _16545_ (.A(_08037_),
    .B(_08349_),
    .Y(_08501_));
 AOI221x1_ASAP7_75t_SL _16546_ (.A1(_08196_),
    .A2(_08501_),
    .B1(_08221_),
    .B2(_08358_),
    .C(_08018_),
    .Y(_08502_));
 OAI21x1_ASAP7_75t_SL _16547_ (.A1(_08218_),
    .A2(_08099_),
    .B(_08159_),
    .Y(_08503_));
 OAI21x1_ASAP7_75t_SL _16548_ (.A1(_08020_),
    .A2(_08503_),
    .B(_08028_),
    .Y(_08504_));
 NAND2x1_ASAP7_75t_SL _16549_ (.A(_08236_),
    .B(_08443_),
    .Y(_08505_));
 OA21x2_ASAP7_75t_SL _16550_ (.A1(_08505_),
    .A2(_08018_),
    .B(_08105_),
    .Y(_08506_));
 NAND3x1_ASAP7_75t_SL _16551_ (.A(_08420_),
    .B(_08018_),
    .C(_08113_),
    .Y(_08507_));
 AOI21x1_ASAP7_75t_SL _16552_ (.A1(_08506_),
    .A2(_08507_),
    .B(_08092_),
    .Y(_08508_));
 OAI21x1_ASAP7_75t_SL _16553_ (.A1(_08502_),
    .A2(_08504_),
    .B(_08508_),
    .Y(_08509_));
 AO21x1_ASAP7_75t_SL _16554_ (.A1(_08115_),
    .A2(_08096_),
    .B(_08314_),
    .Y(_08510_));
 NAND2x1_ASAP7_75t_SL _16555_ (.A(_08018_),
    .B(_08510_),
    .Y(_08511_));
 AO21x1_ASAP7_75t_SL _16556_ (.A1(_08442_),
    .A2(_08037_),
    .B(_08018_),
    .Y(_08512_));
 NOR2x1_ASAP7_75t_SL _16557_ (.A(_08309_),
    .B(_08439_),
    .Y(_08513_));
 OA21x2_ASAP7_75t_SL _16558_ (.A1(_08512_),
    .A2(_08513_),
    .B(_08105_),
    .Y(_08514_));
 AOI21x1_ASAP7_75t_SL _16559_ (.A1(_08511_),
    .A2(_08514_),
    .B(_08071_),
    .Y(_08515_));
 AO21x1_ASAP7_75t_SL _16560_ (.A1(_00973_),
    .A2(_00972_),
    .B(_08089_),
    .Y(_08516_));
 OR3x1_ASAP7_75t_SL _16561_ (.A(_08137_),
    .B(_08036_),
    .C(_08161_),
    .Y(_08517_));
 AO21x1_ASAP7_75t_SL _16562_ (.A1(_08516_),
    .A2(_08517_),
    .B(_08018_),
    .Y(_08518_));
 NAND2x1_ASAP7_75t_SL _16563_ (.A(_08036_),
    .B(_00973_),
    .Y(_08519_));
 AO21x1_ASAP7_75t_SL _16564_ (.A1(_00972_),
    .A2(_08519_),
    .B(_08152_),
    .Y(_08520_));
 OA21x2_ASAP7_75t_SL _16565_ (.A1(_08520_),
    .A2(_08020_),
    .B(_08028_),
    .Y(_08521_));
 NAND2x1_ASAP7_75t_SL _16566_ (.A(_08518_),
    .B(_08521_),
    .Y(_08522_));
 AOI21x1_ASAP7_75t_SL _16567_ (.A1(_08515_),
    .A2(_08522_),
    .B(_08263_),
    .Y(_08523_));
 NAND2x1_ASAP7_75t_SL _16568_ (.A(_08509_),
    .B(_08523_),
    .Y(_08524_));
 NAND2x1_ASAP7_75t_SL _16569_ (.A(_08500_),
    .B(_08524_),
    .Y(_00005_));
 AO21x1_ASAP7_75t_SL _16570_ (.A1(_08197_),
    .A2(_08266_),
    .B(_08408_),
    .Y(_08525_));
 AOI21x1_ASAP7_75t_SL _16571_ (.A1(_08020_),
    .A2(_08525_),
    .B(_08330_),
    .Y(_08526_));
 INVx1_ASAP7_75t_SL _16572_ (.A(_08095_),
    .Y(_08527_));
 AO21x1_ASAP7_75t_SL _16573_ (.A1(_08527_),
    .A2(_08300_),
    .B(_08036_),
    .Y(_08528_));
 NAND2x1_ASAP7_75t_SL _16574_ (.A(_08257_),
    .B(_08528_),
    .Y(_08529_));
 AOI21x1_ASAP7_75t_SL _16575_ (.A1(_00987_),
    .A2(_08037_),
    .B(_08020_),
    .Y(_08530_));
 AOI21x1_ASAP7_75t_SL _16576_ (.A1(_08530_),
    .A2(_08489_),
    .B(_08105_),
    .Y(_08531_));
 NAND2x1_ASAP7_75t_SL _16577_ (.A(_08529_),
    .B(_08531_),
    .Y(_08532_));
 OAI21x1_ASAP7_75t_SL _16578_ (.A1(_08028_),
    .A2(_08526_),
    .B(_08532_),
    .Y(_08533_));
 OAI21x1_ASAP7_75t_SL _16579_ (.A1(_08071_),
    .A2(_08533_),
    .B(_08263_),
    .Y(_08534_));
 NAND2x1_ASAP7_75t_SL _16580_ (.A(_00986_),
    .B(_08037_),
    .Y(_08535_));
 AND2x2_ASAP7_75t_SL _16581_ (.A(_08133_),
    .B(_08036_),
    .Y(_08536_));
 NOR2x1_ASAP7_75t_SL _16582_ (.A(_08536_),
    .B(_08419_),
    .Y(_08537_));
 AOI22x1_ASAP7_75t_SL _16583_ (.A1(_08103_),
    .A2(_08535_),
    .B1(_08537_),
    .B2(_08018_),
    .Y(_08538_));
 NAND2x1_ASAP7_75t_SL _16584_ (.A(_08122_),
    .B(_08208_),
    .Y(_08539_));
 NOR2x1_ASAP7_75t_SL _16585_ (.A(_08036_),
    .B(_08539_),
    .Y(_08540_));
 AND2x2_ASAP7_75t_SL _16586_ (.A(_08250_),
    .B(_08208_),
    .Y(_08541_));
 OAI21x1_ASAP7_75t_SL _16587_ (.A1(_08540_),
    .A2(_08541_),
    .B(_08020_),
    .Y(_08542_));
 OAI21x1_ASAP7_75t_SL _16588_ (.A1(_08036_),
    .A2(_08539_),
    .B(_08018_),
    .Y(_08543_));
 AO21x1_ASAP7_75t_SL _16589_ (.A1(_08166_),
    .A2(_08236_),
    .B(_08543_),
    .Y(_08544_));
 AOI21x1_ASAP7_75t_SL _16590_ (.A1(_08542_),
    .A2(_08544_),
    .B(_08105_),
    .Y(_08545_));
 AOI211x1_ASAP7_75t_SL _16591_ (.A1(_08538_),
    .A2(_08105_),
    .B(_08545_),
    .C(_08092_),
    .Y(_08546_));
 AOI211x1_ASAP7_75t_SL _16592_ (.A1(_08178_),
    .A2(_08124_),
    .B(_08419_),
    .C(_08018_),
    .Y(_08547_));
 AND2x2_ASAP7_75t_SL _16593_ (.A(_08063_),
    .B(_00974_),
    .Y(_08548_));
 OA21x2_ASAP7_75t_SL _16594_ (.A1(_08548_),
    .A2(_08157_),
    .B(_08037_),
    .Y(_08549_));
 AND2x2_ASAP7_75t_SL _16595_ (.A(_08250_),
    .B(_08196_),
    .Y(_08550_));
 NOR2x1_ASAP7_75t_SL _16596_ (.A(_08549_),
    .B(_08550_),
    .Y(_08551_));
 AO21x1_ASAP7_75t_SL _16597_ (.A1(_08551_),
    .A2(_08018_),
    .B(_08028_),
    .Y(_08552_));
 OA21x2_ASAP7_75t_SL _16598_ (.A1(_08037_),
    .A2(_00972_),
    .B(_08018_),
    .Y(_08553_));
 AO21x1_ASAP7_75t_SL _16599_ (.A1(_08266_),
    .A2(_08430_),
    .B(_08036_),
    .Y(_08554_));
 AOI21x1_ASAP7_75t_SL _16600_ (.A1(_08553_),
    .A2(_08554_),
    .B(_08105_),
    .Y(_08555_));
 AO21x1_ASAP7_75t_SL _16601_ (.A1(_08213_),
    .A2(_08325_),
    .B(_08036_),
    .Y(_08556_));
 NAND3x1_ASAP7_75t_SL _16602_ (.A(_08556_),
    .B(_08020_),
    .C(_08360_),
    .Y(_08557_));
 AOI21x1_ASAP7_75t_SL _16603_ (.A1(_08555_),
    .A2(_08557_),
    .B(_08092_),
    .Y(_08558_));
 OAI21x1_ASAP7_75t_SL _16604_ (.A1(_08547_),
    .A2(_08552_),
    .B(_08558_),
    .Y(_08559_));
 NOR2x1_ASAP7_75t_SL _16605_ (.A(_08018_),
    .B(_08355_),
    .Y(_08560_));
 NAND2x1_ASAP7_75t_SL _16606_ (.A(_08527_),
    .B(_08101_),
    .Y(_08561_));
 AOI21x1_ASAP7_75t_SL _16607_ (.A1(_08560_),
    .A2(_08561_),
    .B(_08105_),
    .Y(_08562_));
 AOI21x1_ASAP7_75t_SL _16608_ (.A1(_08249_),
    .A2(_08322_),
    .B(_08020_),
    .Y(_08563_));
 OAI21x1_ASAP7_75t_SL _16609_ (.A1(_08165_),
    .A2(_08369_),
    .B(_08563_),
    .Y(_08564_));
 AOI21x1_ASAP7_75t_SL _16610_ (.A1(_08562_),
    .A2(_08564_),
    .B(_08071_),
    .Y(_08565_));
 AOI22x1_ASAP7_75t_SL _16611_ (.A1(_08124_),
    .A2(_08178_),
    .B1(_08458_),
    .B2(_08208_),
    .Y(_08566_));
 NAND2x1_ASAP7_75t_SL _16612_ (.A(_08018_),
    .B(_08566_),
    .Y(_08567_));
 AND2x2_ASAP7_75t_SL _16613_ (.A(_08458_),
    .B(_08230_),
    .Y(_08568_));
 AO21x1_ASAP7_75t_SL _16614_ (.A1(_08137_),
    .A2(_08036_),
    .B(_08018_),
    .Y(_08569_));
 OA21x2_ASAP7_75t_SL _16615_ (.A1(_08568_),
    .A2(_08569_),
    .B(_08105_),
    .Y(_08570_));
 NAND2x1_ASAP7_75t_SL _16616_ (.A(_08567_),
    .B(_08570_),
    .Y(_08571_));
 AOI21x1_ASAP7_75t_SL _16617_ (.A1(_08565_),
    .A2(_08571_),
    .B(_08263_),
    .Y(_08572_));
 NAND2x1_ASAP7_75t_SL _16618_ (.A(_08559_),
    .B(_08572_),
    .Y(_08573_));
 OAI21x1_ASAP7_75t_SL _16619_ (.A1(_08534_),
    .A2(_08546_),
    .B(_08573_),
    .Y(_00006_));
 AO21x1_ASAP7_75t_SL _16620_ (.A1(_08197_),
    .A2(_08266_),
    .B(_08250_),
    .Y(_08574_));
 OA21x2_ASAP7_75t_SL _16621_ (.A1(_08574_),
    .A2(_08020_),
    .B(_08028_),
    .Y(_08575_));
 OA21x2_ASAP7_75t_SL _16622_ (.A1(_08548_),
    .A2(_08139_),
    .B(_08037_),
    .Y(_08576_));
 NOR2x1_ASAP7_75t_SL _16623_ (.A(_08349_),
    .B(_08089_),
    .Y(_08577_));
 OR3x1_ASAP7_75t_SL _16624_ (.A(_08576_),
    .B(_08018_),
    .C(_08577_),
    .Y(_08578_));
 OAI21x1_ASAP7_75t_SL _16625_ (.A1(_08346_),
    .A2(_08550_),
    .B(_08018_),
    .Y(_08579_));
 AO21x1_ASAP7_75t_SL _16626_ (.A1(_08383_),
    .A2(_08178_),
    .B(_08036_),
    .Y(_08580_));
 AO21x1_ASAP7_75t_SL _16627_ (.A1(_08403_),
    .A2(_08580_),
    .B(_08018_),
    .Y(_08581_));
 AOI21x1_ASAP7_75t_SL _16628_ (.A1(_08579_),
    .A2(_08581_),
    .B(_08028_),
    .Y(_08582_));
 AOI211x1_ASAP7_75t_SL _16629_ (.A1(_08575_),
    .A2(_08578_),
    .B(_08582_),
    .C(_08092_),
    .Y(_08583_));
 INVx1_ASAP7_75t_SL _16630_ (.A(_08519_),
    .Y(_08584_));
 AO21x1_ASAP7_75t_SL _16631_ (.A1(_08221_),
    .A2(_08151_),
    .B(_08584_),
    .Y(_08585_));
 OAI21x1_ASAP7_75t_SL _16632_ (.A1(_08018_),
    .A2(_08585_),
    .B(_08028_),
    .Y(_08586_));
 AOI21x1_ASAP7_75t_SL _16633_ (.A1(_08166_),
    .A2(_08110_),
    .B(_08426_),
    .Y(_08587_));
 NAND2x1_ASAP7_75t_SL _16634_ (.A(_08110_),
    .B(_08322_),
    .Y(_08588_));
 NOR2x1_ASAP7_75t_SL _16635_ (.A(_08018_),
    .B(_08458_),
    .Y(_08589_));
 INVx1_ASAP7_75t_SL _16636_ (.A(_08147_),
    .Y(_08590_));
 OAI21x1_ASAP7_75t_SL _16637_ (.A1(_08590_),
    .A2(_08162_),
    .B(_08105_),
    .Y(_08591_));
 AO21x1_ASAP7_75t_SL _16638_ (.A1(_08588_),
    .A2(_08589_),
    .B(_08591_),
    .Y(_08592_));
 OAI21x1_ASAP7_75t_SL _16639_ (.A1(_08586_),
    .A2(_08587_),
    .B(_08592_),
    .Y(_08593_));
 OAI21x1_ASAP7_75t_SL _16640_ (.A1(_08071_),
    .A2(_08593_),
    .B(_08263_),
    .Y(_08594_));
 AO21x1_ASAP7_75t_SL _16641_ (.A1(_08527_),
    .A2(_08178_),
    .B(_08036_),
    .Y(_08595_));
 AND3x1_ASAP7_75t_SL _16642_ (.A(_08595_),
    .B(_08257_),
    .C(_08350_),
    .Y(_08596_));
 NOR2x1_ASAP7_75t_SL _16643_ (.A(_08037_),
    .B(_08148_),
    .Y(_08597_));
 AO21x1_ASAP7_75t_SL _16644_ (.A1(_08036_),
    .A2(_08212_),
    .B(_08434_),
    .Y(_08598_));
 OAI21x1_ASAP7_75t_SL _16645_ (.A1(_08597_),
    .A2(_08598_),
    .B(_08105_),
    .Y(_08599_));
 NAND2x1_ASAP7_75t_SL _16646_ (.A(_00974_),
    .B(_08037_),
    .Y(_08600_));
 OA21x2_ASAP7_75t_SL _16647_ (.A1(_08325_),
    .A2(_08037_),
    .B(_08018_),
    .Y(_08601_));
 AOI21x1_ASAP7_75t_SL _16648_ (.A1(_08600_),
    .A2(_08601_),
    .B(_08105_),
    .Y(_08602_));
 NAND3x1_ASAP7_75t_SL _16649_ (.A(_08229_),
    .B(_08464_),
    .C(_08156_),
    .Y(_08603_));
 AOI21x1_ASAP7_75t_SL _16650_ (.A1(_08602_),
    .A2(_08603_),
    .B(_08071_),
    .Y(_08604_));
 OAI21x1_ASAP7_75t_SL _16651_ (.A1(_08596_),
    .A2(_08599_),
    .B(_08604_),
    .Y(_08605_));
 OA21x2_ASAP7_75t_SL _16652_ (.A1(_08037_),
    .A2(_00979_),
    .B(_08020_),
    .Y(_08606_));
 NAND2x1_ASAP7_75t_SL _16653_ (.A(_08606_),
    .B(_08554_),
    .Y(_08607_));
 OA21x2_ASAP7_75t_SL _16654_ (.A1(_08036_),
    .A2(_08151_),
    .B(_08140_),
    .Y(_08608_));
 AOI21x1_ASAP7_75t_SL _16655_ (.A1(_08601_),
    .A2(_08608_),
    .B(_08028_),
    .Y(_08609_));
 AOI21x1_ASAP7_75t_SL _16656_ (.A1(_08607_),
    .A2(_08609_),
    .B(_08092_),
    .Y(_08610_));
 AO21x1_ASAP7_75t_SL _16657_ (.A1(_08138_),
    .A2(_08527_),
    .B(_08036_),
    .Y(_08611_));
 INVx1_ASAP7_75t_SL _16658_ (.A(_08548_),
    .Y(_08612_));
 AO21x1_ASAP7_75t_SL _16659_ (.A1(_08612_),
    .A2(_08140_),
    .B(_08037_),
    .Y(_08613_));
 NAND2x1_ASAP7_75t_SL _16660_ (.A(_08611_),
    .B(_08613_),
    .Y(_08614_));
 AOI21x1_ASAP7_75t_SL _16661_ (.A1(_08196_),
    .A2(_08221_),
    .B(_08018_),
    .Y(_08615_));
 AO21x1_ASAP7_75t_SL _16662_ (.A1(_08612_),
    .A2(_08266_),
    .B(_08037_),
    .Y(_08616_));
 AOI21x1_ASAP7_75t_SL _16663_ (.A1(_08615_),
    .A2(_08616_),
    .B(_08105_),
    .Y(_08617_));
 OAI21x1_ASAP7_75t_SL _16664_ (.A1(_08020_),
    .A2(_08614_),
    .B(_08617_),
    .Y(_08618_));
 AOI21x1_ASAP7_75t_SL _16665_ (.A1(_08610_),
    .A2(_08618_),
    .B(_08263_),
    .Y(_08619_));
 NAND2x1_ASAP7_75t_SL _16666_ (.A(_08605_),
    .B(_08619_),
    .Y(_08620_));
 OAI21x1_ASAP7_75t_SL _16667_ (.A1(_08583_),
    .A2(_08594_),
    .B(_08620_),
    .Y(_00007_));
 XOR2x1_ASAP7_75t_SL _16668_ (.A(_00838_),
    .Y(_08621_),
    .B(_00421_));
 AND2x2_ASAP7_75t_R _16674_ (.A(ld),
    .B(key[96]),
    .Y(_08627_));
 AO21x1_ASAP7_75t_R _16675_ (.A1(_08621_),
    .A2(_08005_),
    .B(_08627_),
    .Y(_00289_));
 XOR2x2_ASAP7_75t_SL _16676_ (.A(_00849_),
    .B(_00422_),
    .Y(_08628_));
 AND2x2_ASAP7_75t_R _16677_ (.A(ld),
    .B(key[97]),
    .Y(_08629_));
 AO21x1_ASAP7_75t_R _16678_ (.A1(_08628_),
    .A2(_08005_),
    .B(_08629_),
    .Y(_00300_));
 XOR2x2_ASAP7_75t_R _16679_ (.A(_00423_),
    .B(_00860_),
    .Y(_08630_));
 AND2x2_ASAP7_75t_R _16680_ (.A(ld),
    .B(key[98]),
    .Y(_08631_));
 AO21x1_ASAP7_75t_R _16681_ (.A1(_08630_),
    .A2(_08005_),
    .B(_08631_),
    .Y(_00311_));
 XOR2x2_ASAP7_75t_R _16682_ (.A(_00424_),
    .B(_00863_),
    .Y(_08632_));
 AND2x2_ASAP7_75t_R _16683_ (.A(ld),
    .B(key[99]),
    .Y(_08633_));
 AO21x1_ASAP7_75t_R _16684_ (.A1(_08632_),
    .A2(_08005_),
    .B(_08633_),
    .Y(_00314_));
 XOR2x2_ASAP7_75t_SL _16685_ (.A(_00425_),
    .B(_00864_),
    .Y(_08634_));
 AND2x2_ASAP7_75t_R _16686_ (.A(ld),
    .B(key[100]),
    .Y(_08635_));
 AO21x1_ASAP7_75t_R _16687_ (.A1(_08634_),
    .A2(_08005_),
    .B(_08635_),
    .Y(_00315_));
 XOR2x2_ASAP7_75t_SL _16688_ (.A(_00426_),
    .B(_00865_),
    .Y(_08636_));
 AND2x2_ASAP7_75t_R _16689_ (.A(ld),
    .B(key[101]),
    .Y(_08637_));
 AO21x1_ASAP7_75t_R _16690_ (.A1(_08636_),
    .A2(_08005_),
    .B(_08637_),
    .Y(_00316_));
 XOR2x2_ASAP7_75t_SL _16691_ (.A(_00427_),
    .B(_00866_),
    .Y(_08638_));
 AND2x2_ASAP7_75t_R _16692_ (.A(ld),
    .B(key[102]),
    .Y(_08639_));
 AO21x1_ASAP7_75t_R _16693_ (.A1(_08638_),
    .A2(_08005_),
    .B(_08639_),
    .Y(_00317_));
 XOR2x2_ASAP7_75t_R _16694_ (.A(_00428_),
    .B(_00867_),
    .Y(_08640_));
 AND2x2_ASAP7_75t_R _16696_ (.A(ld),
    .B(key[103]),
    .Y(_08642_));
 AO21x1_ASAP7_75t_R _16697_ (.A1(_08640_),
    .A2(_08005_),
    .B(_08642_),
    .Y(_00318_));
 XOR2x2_ASAP7_75t_SL _16698_ (.A(_00429_),
    .B(_00868_),
    .Y(_08643_));
 AND2x2_ASAP7_75t_R _16699_ (.A(ld),
    .B(key[104]),
    .Y(_08644_));
 AO21x1_ASAP7_75t_R _16700_ (.A1(_08643_),
    .A2(_08005_),
    .B(_08644_),
    .Y(_00319_));
 XOR2x2_ASAP7_75t_R _16701_ (.A(_00430_),
    .B(_00869_),
    .Y(_08645_));
 AND2x2_ASAP7_75t_R _16703_ (.A(ld),
    .B(key[105]),
    .Y(_08647_));
 AO21x1_ASAP7_75t_R _16704_ (.A1(_08645_),
    .A2(_08005_),
    .B(_08647_),
    .Y(_00320_));
 XOR2x2_ASAP7_75t_R _16705_ (.A(_00431_),
    .B(_00839_),
    .Y(_08648_));
 AND2x2_ASAP7_75t_R _16706_ (.A(ld),
    .B(key[106]),
    .Y(_08649_));
 AO21x1_ASAP7_75t_R _16707_ (.A1(_08648_),
    .A2(_08005_),
    .B(_08649_),
    .Y(_00290_));
 XOR2x2_ASAP7_75t_R _16708_ (.A(_00432_),
    .B(_00840_),
    .Y(_08650_));
 AND2x2_ASAP7_75t_R _16709_ (.A(ld),
    .B(key[107]),
    .Y(_08651_));
 AO21x1_ASAP7_75t_R _16710_ (.A1(_08650_),
    .A2(_08005_),
    .B(_08651_),
    .Y(_00291_));
 XOR2x2_ASAP7_75t_SL _16711_ (.A(_00433_),
    .B(_00841_),
    .Y(_08652_));
 AND2x2_ASAP7_75t_R _16712_ (.A(ld),
    .B(key[108]),
    .Y(_08653_));
 AO21x1_ASAP7_75t_R _16713_ (.A1(_08652_),
    .A2(_08005_),
    .B(_08653_),
    .Y(_00292_));
 XOR2x2_ASAP7_75t_SL _16714_ (.A(_00434_),
    .B(_00842_),
    .Y(_08654_));
 AND2x2_ASAP7_75t_R _16715_ (.A(ld),
    .B(key[109]),
    .Y(_08655_));
 AO21x1_ASAP7_75t_R _16716_ (.A1(_08654_),
    .A2(_08005_),
    .B(_08655_),
    .Y(_00293_));
 XOR2x2_ASAP7_75t_SL _16717_ (.A(_00435_),
    .B(_00843_),
    .Y(_08656_));
 AND2x2_ASAP7_75t_R _16718_ (.A(ld),
    .B(key[110]),
    .Y(_08657_));
 AO21x1_ASAP7_75t_R _16719_ (.A1(_08656_),
    .A2(_08005_),
    .B(_08657_),
    .Y(_00294_));
 XOR2x2_ASAP7_75t_SL _16720_ (.A(_00436_),
    .B(_00844_),
    .Y(_08658_));
 AND2x2_ASAP7_75t_R _16721_ (.A(ld),
    .B(key[111]),
    .Y(_08659_));
 AO21x1_ASAP7_75t_R _16722_ (.A1(_08658_),
    .A2(_08005_),
    .B(_08659_),
    .Y(_00295_));
 XOR2x2_ASAP7_75t_R _16723_ (.A(_00437_),
    .B(_00845_),
    .Y(_08660_));
 AND2x2_ASAP7_75t_R _16724_ (.A(ld),
    .B(key[112]),
    .Y(_08661_));
 AO21x1_ASAP7_75t_R _16725_ (.A1(_08660_),
    .A2(_08005_),
    .B(_08661_),
    .Y(_00296_));
 XOR2x2_ASAP7_75t_R _16726_ (.A(_00438_),
    .B(_00846_),
    .Y(_08662_));
 AND2x2_ASAP7_75t_R _16728_ (.A(ld),
    .B(key[113]),
    .Y(_08664_));
 AO21x1_ASAP7_75t_R _16729_ (.A1(_08662_),
    .A2(_08005_),
    .B(_08664_),
    .Y(_00297_));
 XNOR2x2_ASAP7_75t_R _16733_ (.A(_00412_),
    .B(_00847_),
    .Y(_08668_));
 NOR2x1_ASAP7_75t_R _16734_ (.A(ld),
    .B(_08668_),
    .Y(_08669_));
 AO21x1_ASAP7_75t_R _16735_ (.A1(ld),
    .A2(key[114]),
    .B(_08669_),
    .Y(_00298_));
 XOR2x2_ASAP7_75t_R _16736_ (.A(_00439_),
    .B(_00848_),
    .Y(_08670_));
 AND2x2_ASAP7_75t_R _16737_ (.A(ld),
    .B(key[115]),
    .Y(_08671_));
 AO21x1_ASAP7_75t_R _16738_ (.A1(_08670_),
    .A2(_08005_),
    .B(_08671_),
    .Y(_00299_));
 XOR2x2_ASAP7_75t_R _16739_ (.A(_00440_),
    .B(_00850_),
    .Y(_08672_));
 AND2x2_ASAP7_75t_R _16741_ (.A(ld),
    .B(key[116]),
    .Y(_08674_));
 AO21x1_ASAP7_75t_R _16742_ (.A1(_08672_),
    .A2(_08005_),
    .B(_08674_),
    .Y(_00301_));
 XOR2x2_ASAP7_75t_R _16743_ (.A(_00441_),
    .B(_00851_),
    .Y(_08675_));
 AND2x2_ASAP7_75t_R _16744_ (.A(ld),
    .B(key[117]),
    .Y(_08676_));
 AO21x1_ASAP7_75t_R _16745_ (.A1(_08675_),
    .A2(_08005_),
    .B(_08676_),
    .Y(_00302_));
 XOR2x2_ASAP7_75t_R _16746_ (.A(_00442_),
    .B(_00852_),
    .Y(_08677_));
 AND2x2_ASAP7_75t_R _16747_ (.A(ld),
    .B(key[118]),
    .Y(_08678_));
 AO21x1_ASAP7_75t_R _16748_ (.A1(_08677_),
    .A2(_08005_),
    .B(_08678_),
    .Y(_00303_));
 XOR2x2_ASAP7_75t_R _16749_ (.A(_00443_),
    .B(_00853_),
    .Y(_08679_));
 AND2x2_ASAP7_75t_R _16750_ (.A(ld),
    .B(key[119]),
    .Y(_08680_));
 AO21x1_ASAP7_75t_R _16751_ (.A1(_08679_),
    .A2(_08005_),
    .B(_08680_),
    .Y(_00304_));
 XOR2x2_ASAP7_75t_SL _16754_ (.A(_00830_),
    .B(_00854_),
    .Y(_08683_));
 XOR2x2_ASAP7_75t_SL _16755_ (.A(_08683_),
    .B(_00413_),
    .Y(_08684_));
 NOR2x1_ASAP7_75t_R _16756_ (.A(ld),
    .B(_08684_),
    .Y(_08685_));
 AO21x1_ASAP7_75t_R _16757_ (.A1(ld),
    .A2(key[120]),
    .B(_08685_),
    .Y(_00305_));
 XOR2x2_ASAP7_75t_SL _16758_ (.A(_00855_),
    .B(_00831_),
    .Y(_08686_));
 XOR2x2_ASAP7_75t_SL _16759_ (.A(_08686_),
    .B(_00414_),
    .Y(_08687_));
 NOR2x1_ASAP7_75t_R _16760_ (.A(ld),
    .B(_08687_),
    .Y(_08688_));
 AO21x1_ASAP7_75t_R _16761_ (.A1(ld),
    .A2(key[121]),
    .B(_08688_),
    .Y(_00306_));
 XOR2x1_ASAP7_75t_SL _16762_ (.A(_00832_),
    .Y(_08689_),
    .B(_00856_));
 XOR2x2_ASAP7_75t_SL _16763_ (.A(_08689_),
    .B(_00415_),
    .Y(_08690_));
 NOR2x1_ASAP7_75t_R _16764_ (.A(ld),
    .B(_08690_),
    .Y(_08691_));
 AO21x1_ASAP7_75t_R _16765_ (.A1(ld),
    .A2(key[122]),
    .B(_08691_),
    .Y(_00307_));
 XOR2x2_ASAP7_75t_SL _16766_ (.A(_00833_),
    .B(_00857_),
    .Y(_08692_));
 XOR2x2_ASAP7_75t_SL _16767_ (.A(_08692_),
    .B(_00416_),
    .Y(_08693_));
 NOR2x1_ASAP7_75t_R _16768_ (.A(ld),
    .B(_08693_),
    .Y(_08694_));
 AO21x1_ASAP7_75t_R _16769_ (.A1(ld),
    .A2(key[123]),
    .B(_08694_),
    .Y(_00308_));
 XOR2x1_ASAP7_75t_SL _16770_ (.A(_00834_),
    .Y(_08695_),
    .B(_00858_));
 XOR2x2_ASAP7_75t_R _16771_ (.A(_08695_),
    .B(_00417_),
    .Y(_08696_));
 NOR2x1_ASAP7_75t_R _16772_ (.A(ld),
    .B(_08696_),
    .Y(_08697_));
 AO21x1_ASAP7_75t_R _16773_ (.A1(ld),
    .A2(key[124]),
    .B(_08697_),
    .Y(_00309_));
 XOR2x2_ASAP7_75t_SL _16774_ (.A(_00835_),
    .B(_00859_),
    .Y(_08698_));
 XOR2x2_ASAP7_75t_R _16775_ (.A(_08698_),
    .B(_00418_),
    .Y(_08699_));
 NOR2x1_ASAP7_75t_R _16776_ (.A(ld),
    .B(_08699_),
    .Y(_08700_));
 AO21x1_ASAP7_75t_R _16777_ (.A1(ld),
    .A2(key[125]),
    .B(_08700_),
    .Y(_00310_));
 XOR2x2_ASAP7_75t_SL _16778_ (.A(_00836_),
    .B(_00861_),
    .Y(_08701_));
 XOR2x2_ASAP7_75t_R _16779_ (.A(_08701_),
    .B(_00419_),
    .Y(_08702_));
 NOR2x1_ASAP7_75t_R _16780_ (.A(ld),
    .B(_08702_),
    .Y(_08703_));
 AO21x1_ASAP7_75t_R _16781_ (.A1(ld),
    .A2(key[126]),
    .B(_08703_),
    .Y(_00312_));
 XOR2x2_ASAP7_75t_SL _16782_ (.A(_00837_),
    .B(_00862_),
    .Y(_08704_));
 XOR2x2_ASAP7_75t_R _16783_ (.A(_08704_),
    .B(_00420_),
    .Y(_08705_));
 NOR2x1_ASAP7_75t_R _16784_ (.A(ld),
    .B(_08705_),
    .Y(_08706_));
 AO21x1_ASAP7_75t_R _16785_ (.A1(ld),
    .A2(key[127]),
    .B(_08706_),
    .Y(_00313_));
 XOR2x2_ASAP7_75t_SL _16788_ (.A(_00870_),
    .B(_08621_),
    .Y(_08709_));
 NOR2x1_ASAP7_75t_R _16789_ (.A(ld),
    .B(_08709_),
    .Y(_08710_));
 AO21x1_ASAP7_75t_R _16790_ (.A1(ld),
    .A2(key[64]),
    .B(_08710_),
    .Y(_00321_));
 XOR2x2_ASAP7_75t_SL _16791_ (.A(_00881_),
    .B(_08628_),
    .Y(_08711_));
 NOR2x1_ASAP7_75t_R _16792_ (.A(ld),
    .B(_08711_),
    .Y(_08712_));
 AO21x1_ASAP7_75t_R _16793_ (.A1(ld),
    .A2(key[65]),
    .B(_08712_),
    .Y(_00332_));
 XOR2x2_ASAP7_75t_R _16795_ (.A(_08630_),
    .B(_00892_),
    .Y(_08714_));
 NOR2x1_ASAP7_75t_R _16796_ (.A(ld),
    .B(_08714_),
    .Y(_08715_));
 AO21x1_ASAP7_75t_R _16797_ (.A1(ld),
    .A2(key[66]),
    .B(_08715_),
    .Y(_00343_));
 XOR2x2_ASAP7_75t_SL _16798_ (.A(_00863_),
    .B(_00895_),
    .Y(_08716_));
 XOR2x2_ASAP7_75t_R _16799_ (.A(_08716_),
    .B(_00424_),
    .Y(_08717_));
 NOR2x1_ASAP7_75t_R _16800_ (.A(ld),
    .B(_08717_),
    .Y(_08718_));
 AO21x1_ASAP7_75t_R _16801_ (.A1(ld),
    .A2(key[67]),
    .B(_08718_),
    .Y(_00346_));
 XOR2x2_ASAP7_75t_SL _16802_ (.A(_08634_),
    .B(_00896_),
    .Y(_08719_));
 NOR2x1_ASAP7_75t_R _16803_ (.A(ld),
    .B(_08719_),
    .Y(_08720_));
 AO21x1_ASAP7_75t_R _16804_ (.A1(ld),
    .A2(key[68]),
    .B(_08720_),
    .Y(_00347_));
 XOR2x2_ASAP7_75t_R _16805_ (.A(_08636_),
    .B(_00897_),
    .Y(_08721_));
 NOR2x1_ASAP7_75t_R _16806_ (.A(ld),
    .B(_08721_),
    .Y(_08722_));
 AO21x1_ASAP7_75t_R _16807_ (.A1(ld),
    .A2(key[69]),
    .B(_08722_),
    .Y(_00348_));
 XOR2x2_ASAP7_75t_R _16808_ (.A(_08638_),
    .B(_00898_),
    .Y(_08723_));
 NOR2x1_ASAP7_75t_R _16809_ (.A(ld),
    .B(_08723_),
    .Y(_08724_));
 AO21x1_ASAP7_75t_R _16810_ (.A1(ld),
    .A2(key[70]),
    .B(_08724_),
    .Y(_00349_));
 XOR2x2_ASAP7_75t_R _16811_ (.A(_08640_),
    .B(_00899_),
    .Y(_08725_));
 NOR2x1_ASAP7_75t_R _16812_ (.A(ld),
    .B(_08725_),
    .Y(_08726_));
 AO21x1_ASAP7_75t_R _16813_ (.A1(ld),
    .A2(key[71]),
    .B(_08726_),
    .Y(_00350_));
 XOR2x2_ASAP7_75t_SL _16814_ (.A(_08643_),
    .B(_00900_),
    .Y(_08727_));
 NOR2x1_ASAP7_75t_R _16815_ (.A(ld),
    .B(_08727_),
    .Y(_08728_));
 AO21x1_ASAP7_75t_R _16816_ (.A1(ld),
    .A2(key[72]),
    .B(_08728_),
    .Y(_00351_));
 INVx1_ASAP7_75t_R _16817_ (.A(_00901_),
    .Y(_08729_));
 OA21x2_ASAP7_75t_R _16818_ (.A1(_08645_),
    .A2(_08729_),
    .B(_08005_),
    .Y(_08730_));
 NAND2x1_ASAP7_75t_R _16819_ (.A(_08729_),
    .B(_08645_),
    .Y(_08731_));
 AO22x1_ASAP7_75t_R _16821_ (.A1(_08730_),
    .A2(_08731_),
    .B1(ld),
    .B2(key[73]),
    .Y(_00352_));
 XOR2x2_ASAP7_75t_R _16822_ (.A(_08648_),
    .B(_00871_),
    .Y(_08733_));
 NOR2x1_ASAP7_75t_R _16823_ (.A(ld),
    .B(_08733_),
    .Y(_08734_));
 AO21x1_ASAP7_75t_R _16824_ (.A1(ld),
    .A2(key[74]),
    .B(_08734_),
    .Y(_00322_));
 XOR2x2_ASAP7_75t_L _16826_ (.A(_00840_),
    .B(_00872_),
    .Y(_08736_));
 XOR2x2_ASAP7_75t_R _16827_ (.A(_08736_),
    .B(_00432_),
    .Y(_08737_));
 NOR2x1_ASAP7_75t_R _16828_ (.A(ld),
    .B(_08737_),
    .Y(_08738_));
 AO21x1_ASAP7_75t_R _16829_ (.A1(ld),
    .A2(key[75]),
    .B(_08738_),
    .Y(_00323_));
 XOR2x2_ASAP7_75t_SL _16830_ (.A(_08652_),
    .B(_00873_),
    .Y(_08739_));
 NOR2x1_ASAP7_75t_R _16831_ (.A(ld),
    .B(_08739_),
    .Y(_08740_));
 AO21x1_ASAP7_75t_R _16832_ (.A1(ld),
    .A2(key[76]),
    .B(_08740_),
    .Y(_00324_));
 XOR2x2_ASAP7_75t_R _16834_ (.A(_08654_),
    .B(_00874_),
    .Y(_08742_));
 NOR2x1_ASAP7_75t_R _16835_ (.A(ld),
    .B(_08742_),
    .Y(_08743_));
 AO21x1_ASAP7_75t_R _16836_ (.A1(ld),
    .A2(key[77]),
    .B(_08743_),
    .Y(_00325_));
 XOR2x2_ASAP7_75t_R _16837_ (.A(_08656_),
    .B(_00875_),
    .Y(_08744_));
 NOR2x1_ASAP7_75t_R _16838_ (.A(ld),
    .B(_08744_),
    .Y(_08745_));
 AO21x1_ASAP7_75t_R _16839_ (.A1(ld),
    .A2(key[78]),
    .B(_08745_),
    .Y(_00326_));
 XOR2x2_ASAP7_75t_R _16840_ (.A(_08658_),
    .B(_00876_),
    .Y(_08746_));
 NOR2x1_ASAP7_75t_R _16841_ (.A(ld),
    .B(_08746_),
    .Y(_08747_));
 AO21x1_ASAP7_75t_R _16842_ (.A1(ld),
    .A2(key[79]),
    .B(_08747_),
    .Y(_00327_));
 XOR2x2_ASAP7_75t_R _16843_ (.A(_08660_),
    .B(_00877_),
    .Y(_08748_));
 NOR2x1_ASAP7_75t_R _16844_ (.A(ld),
    .B(_08748_),
    .Y(_08749_));
 AO21x1_ASAP7_75t_R _16845_ (.A1(ld),
    .A2(key[80]),
    .B(_08749_),
    .Y(_00328_));
 XOR2x2_ASAP7_75t_R _16846_ (.A(_08662_),
    .B(_00878_),
    .Y(_08750_));
 NOR2x1_ASAP7_75t_R _16847_ (.A(ld),
    .B(_08750_),
    .Y(_08751_));
 AO21x1_ASAP7_75t_R _16848_ (.A1(ld),
    .A2(key[81]),
    .B(_08751_),
    .Y(_00329_));
 XOR2x2_ASAP7_75t_R _16849_ (.A(_08056_),
    .B(_00412_),
    .Y(_08752_));
 NOR2x1_ASAP7_75t_R _16850_ (.A(ld),
    .B(_08752_),
    .Y(_08753_));
 AO21x1_ASAP7_75t_R _16851_ (.A1(ld),
    .A2(key[82]),
    .B(_08753_),
    .Y(_00330_));
 XOR2x2_ASAP7_75t_R _16852_ (.A(_08670_),
    .B(_00880_),
    .Y(_08754_));
 NOR2x1_ASAP7_75t_R _16853_ (.A(ld),
    .B(_08754_),
    .Y(_08755_));
 AO21x1_ASAP7_75t_R _16854_ (.A1(ld),
    .A2(key[83]),
    .B(_08755_),
    .Y(_00331_));
 XOR2x2_ASAP7_75t_R _16855_ (.A(_08014_),
    .B(_00440_),
    .Y(_08756_));
 NOR2x1_ASAP7_75t_R _16856_ (.A(ld),
    .B(_08756_),
    .Y(_08757_));
 AO21x1_ASAP7_75t_R _16857_ (.A1(ld),
    .A2(key[84]),
    .B(_08757_),
    .Y(_00333_));
 XOR2x2_ASAP7_75t_R _16859_ (.A(_08675_),
    .B(_00883_),
    .Y(_08759_));
 NOR2x1_ASAP7_75t_R _16860_ (.A(ld),
    .B(_08759_),
    .Y(_08760_));
 AO21x1_ASAP7_75t_R _16861_ (.A1(ld),
    .A2(key[85]),
    .B(_08760_),
    .Y(_00334_));
 XOR2x2_ASAP7_75t_R _16862_ (.A(_08068_),
    .B(_00442_),
    .Y(_08761_));
 NOR2x1_ASAP7_75t_R _16863_ (.A(ld),
    .B(_08761_),
    .Y(_08762_));
 AO21x1_ASAP7_75t_R _16864_ (.A1(ld),
    .A2(key[86]),
    .B(_08762_),
    .Y(_00335_));
 XOR2x2_ASAP7_75t_R _16866_ (.A(_08075_),
    .B(_00443_),
    .Y(_08764_));
 NOR2x1_ASAP7_75t_R _16867_ (.A(ld),
    .B(_08764_),
    .Y(_08765_));
 AO21x1_ASAP7_75t_R _16868_ (.A1(ld),
    .A2(key[87]),
    .B(_08765_),
    .Y(_00336_));
 XOR2x2_ASAP7_75t_SL _16869_ (.A(_08684_),
    .B(_00886_),
    .Y(_08766_));
 AND2x2_ASAP7_75t_R _16870_ (.A(ld),
    .B(key[88]),
    .Y(_08767_));
 AO21x1_ASAP7_75t_R _16871_ (.A1(_08766_),
    .A2(_08005_),
    .B(_08767_),
    .Y(_00337_));
 INVx1_ASAP7_75t_R _16872_ (.A(_00887_),
    .Y(_08768_));
 XOR2x2_ASAP7_75t_SL _16873_ (.A(_08768_),
    .B(_08687_),
    .Y(_08769_));
 NOR2x1_ASAP7_75t_R _16874_ (.A(ld),
    .B(_08769_),
    .Y(_08770_));
 AO21x1_ASAP7_75t_R _16875_ (.A1(ld),
    .A2(key[89]),
    .B(_08770_),
    .Y(_00338_));
 XOR2x1_ASAP7_75t_SL _16876_ (.A(_08690_),
    .Y(_08771_),
    .B(_00888_));
 AND2x2_ASAP7_75t_R _16877_ (.A(ld),
    .B(key[90]),
    .Y(_08772_));
 AO21x1_ASAP7_75t_R _16878_ (.A1(_08771_),
    .A2(_08005_),
    .B(_08772_),
    .Y(_00339_));
 XOR2x2_ASAP7_75t_SL _16879_ (.A(_08693_),
    .B(_00889_),
    .Y(_08773_));
 AND2x2_ASAP7_75t_R _16880_ (.A(ld),
    .B(key[91]),
    .Y(_08774_));
 AO21x1_ASAP7_75t_R _16881_ (.A1(_08773_),
    .A2(_08005_),
    .B(_08774_),
    .Y(_00340_));
 INVx1_ASAP7_75t_R _16882_ (.A(_00890_),
    .Y(_08775_));
 XOR2x2_ASAP7_75t_R _16883_ (.A(_08696_),
    .B(_08775_),
    .Y(_08776_));
 NOR2x1_ASAP7_75t_R _16884_ (.A(ld),
    .B(_08776_),
    .Y(_08777_));
 AO21x1_ASAP7_75t_R _16885_ (.A1(ld),
    .A2(key[92]),
    .B(_08777_),
    .Y(_00341_));
 INVx1_ASAP7_75t_R _16886_ (.A(_00891_),
    .Y(_08778_));
 XOR2x2_ASAP7_75t_SL _16887_ (.A(_08699_),
    .B(_08778_),
    .Y(_08779_));
 NOR2x1_ASAP7_75t_R _16888_ (.A(ld),
    .B(_08779_),
    .Y(_08780_));
 AO21x1_ASAP7_75t_R _16889_ (.A1(ld),
    .A2(key[93]),
    .B(_08780_),
    .Y(_00342_));
 XNOR2x2_ASAP7_75t_SL _16890_ (.A(_00893_),
    .B(_08702_),
    .Y(_08781_));
 NOR2x1_ASAP7_75t_R _16891_ (.A(ld),
    .B(_08781_),
    .Y(_08782_));
 AO21x1_ASAP7_75t_R _16892_ (.A1(ld),
    .A2(key[94]),
    .B(_08782_),
    .Y(_00344_));
 XNOR2x2_ASAP7_75t_R _16893_ (.A(_00894_),
    .B(_08705_),
    .Y(_08783_));
 NOR2x1_ASAP7_75t_R _16894_ (.A(ld),
    .B(_08783_),
    .Y(_08784_));
 AO21x1_ASAP7_75t_R _16895_ (.A1(ld),
    .A2(key[95]),
    .B(_08784_),
    .Y(_00345_));
 XOR2x2_ASAP7_75t_SL _16896_ (.A(_00902_),
    .B(_08709_),
    .Y(_08785_));
 AND2x2_ASAP7_75t_R _16897_ (.A(ld),
    .B(key[32]),
    .Y(_08786_));
 AO21x1_ASAP7_75t_R _16898_ (.A1(_08785_),
    .A2(_08005_),
    .B(_08786_),
    .Y(_00353_));
 XOR2x2_ASAP7_75t_SL _16899_ (.A(_00913_),
    .B(_08711_),
    .Y(_08787_));
 AND2x2_ASAP7_75t_R _16901_ (.A(ld),
    .B(key[33]),
    .Y(_08789_));
 AO21x1_ASAP7_75t_R _16902_ (.A1(_08787_),
    .A2(_08005_),
    .B(_08789_),
    .Y(_00364_));
 INVx1_ASAP7_75t_R _16903_ (.A(_00924_),
    .Y(_08790_));
 AO21x1_ASAP7_75t_R _16905_ (.A1(_08714_),
    .A2(_08790_),
    .B(ld),
    .Y(_08792_));
 NOR2x1_ASAP7_75t_R _16906_ (.A(_08790_),
    .B(_08714_),
    .Y(_08793_));
 OA22x2_ASAP7_75t_R _16907_ (.A1(_08005_),
    .A2(key[34]),
    .B1(_08792_),
    .B2(_08793_),
    .Y(_00375_));
 XOR2x2_ASAP7_75t_R _16908_ (.A(_00424_),
    .B(_00927_),
    .Y(_08794_));
 XOR2x2_ASAP7_75t_SL _16909_ (.A(_08716_),
    .B(_08794_),
    .Y(_08795_));
 AND2x2_ASAP7_75t_R _16910_ (.A(ld),
    .B(key[35]),
    .Y(_08796_));
 AO21x1_ASAP7_75t_R _16911_ (.A1(_08795_),
    .A2(_08005_),
    .B(_08796_),
    .Y(_00378_));
 XOR2x2_ASAP7_75t_SL _16912_ (.A(_08719_),
    .B(_00928_),
    .Y(_08797_));
 AND2x2_ASAP7_75t_R _16914_ (.A(ld),
    .B(key[36]),
    .Y(_08799_));
 AO21x1_ASAP7_75t_R _16915_ (.A1(_08797_),
    .A2(_08005_),
    .B(_08799_),
    .Y(_00379_));
 XOR2x2_ASAP7_75t_R _16916_ (.A(_08721_),
    .B(_00929_),
    .Y(_08800_));
 AND2x2_ASAP7_75t_R _16917_ (.A(ld),
    .B(key[37]),
    .Y(_08801_));
 AO21x1_ASAP7_75t_R _16918_ (.A1(_08800_),
    .A2(_08005_),
    .B(_08801_),
    .Y(_00380_));
 XOR2x2_ASAP7_75t_R _16919_ (.A(_08723_),
    .B(_00930_),
    .Y(_08802_));
 AND2x2_ASAP7_75t_R _16920_ (.A(ld),
    .B(key[38]),
    .Y(_08803_));
 AO21x1_ASAP7_75t_R _16921_ (.A1(_08802_),
    .A2(_08005_),
    .B(_08803_),
    .Y(_00381_));
 XOR2x2_ASAP7_75t_R _16922_ (.A(_08725_),
    .B(_00931_),
    .Y(_08804_));
 AND2x2_ASAP7_75t_R _16923_ (.A(ld),
    .B(key[39]),
    .Y(_08805_));
 AO21x1_ASAP7_75t_R _16924_ (.A1(_08804_),
    .A2(_08005_),
    .B(_08805_),
    .Y(_00382_));
 XOR2x2_ASAP7_75t_SL _16925_ (.A(_08727_),
    .B(_00932_),
    .Y(_08806_));
 AND2x2_ASAP7_75t_R _16926_ (.A(ld),
    .B(key[40]),
    .Y(_08807_));
 AO21x1_ASAP7_75t_R _16927_ (.A1(_08806_),
    .A2(_08005_),
    .B(_08807_),
    .Y(_00383_));
 XOR2x2_ASAP7_75t_SL _16928_ (.A(_00933_),
    .B(_00901_),
    .Y(_08808_));
 XOR2x2_ASAP7_75t_R _16929_ (.A(_08645_),
    .B(_08808_),
    .Y(_08809_));
 AND2x2_ASAP7_75t_R _16930_ (.A(ld),
    .B(key[41]),
    .Y(_08810_));
 AO21x1_ASAP7_75t_R _16931_ (.A1(_08809_),
    .A2(_08005_),
    .B(_08810_),
    .Y(_00384_));
 INVx1_ASAP7_75t_R _16932_ (.A(_00903_),
    .Y(_08811_));
 AO21x1_ASAP7_75t_R _16933_ (.A1(_08733_),
    .A2(_08811_),
    .B(ld),
    .Y(_08812_));
 NOR2x1_ASAP7_75t_R _16934_ (.A(_08811_),
    .B(_08733_),
    .Y(_08813_));
 OA22x2_ASAP7_75t_R _16935_ (.A1(_08005_),
    .A2(key[42]),
    .B1(_08812_),
    .B2(_08813_),
    .Y(_00354_));
 XOR2x2_ASAP7_75t_L _16936_ (.A(_00432_),
    .B(_00904_),
    .Y(_08814_));
 XOR2x2_ASAP7_75t_SL _16937_ (.A(_08736_),
    .B(_08814_),
    .Y(_08815_));
 AND2x2_ASAP7_75t_R _16938_ (.A(ld),
    .B(key[43]),
    .Y(_08816_));
 AO21x1_ASAP7_75t_R _16939_ (.A1(_08815_),
    .A2(_08005_),
    .B(_08816_),
    .Y(_00355_));
 XOR2x2_ASAP7_75t_SL _16940_ (.A(_08739_),
    .B(_00905_),
    .Y(_08817_));
 AND2x2_ASAP7_75t_R _16941_ (.A(ld),
    .B(key[44]),
    .Y(_08818_));
 AO21x1_ASAP7_75t_R _16942_ (.A1(_08817_),
    .A2(_08005_),
    .B(_08818_),
    .Y(_00356_));
 XOR2x2_ASAP7_75t_SL _16943_ (.A(_08742_),
    .B(_00906_),
    .Y(_08819_));
 AND2x2_ASAP7_75t_R _16945_ (.A(ld),
    .B(key[45]),
    .Y(_08821_));
 AO21x1_ASAP7_75t_R _16946_ (.A1(_08819_),
    .A2(_08005_),
    .B(_08821_),
    .Y(_00357_));
 XOR2x2_ASAP7_75t_SL _16947_ (.A(_08744_),
    .B(_00907_),
    .Y(_08822_));
 AND2x2_ASAP7_75t_R _16948_ (.A(ld),
    .B(key[46]),
    .Y(_08823_));
 AO21x1_ASAP7_75t_R _16949_ (.A1(_08822_),
    .A2(_08005_),
    .B(_08823_),
    .Y(_00358_));
 XOR2x2_ASAP7_75t_SL _16950_ (.A(_08746_),
    .B(_00908_),
    .Y(_08824_));
 AND2x2_ASAP7_75t_R _16952_ (.A(ld),
    .B(key[47]),
    .Y(_08826_));
 AO21x1_ASAP7_75t_R _16953_ (.A1(_08824_),
    .A2(_08005_),
    .B(_08826_),
    .Y(_00359_));
 XOR2x2_ASAP7_75t_R _16954_ (.A(_08748_),
    .B(_00909_),
    .Y(_08827_));
 AND2x2_ASAP7_75t_R _16955_ (.A(ld),
    .B(key[48]),
    .Y(_08828_));
 AO21x1_ASAP7_75t_R _16956_ (.A1(_08827_),
    .A2(_08005_),
    .B(_08828_),
    .Y(_00360_));
 XOR2x2_ASAP7_75t_R _16957_ (.A(_08750_),
    .B(_00910_),
    .Y(_08829_));
 AND2x2_ASAP7_75t_R _16958_ (.A(ld),
    .B(key[49]),
    .Y(_08830_));
 AO21x1_ASAP7_75t_R _16959_ (.A1(_08829_),
    .A2(_08005_),
    .B(_08830_),
    .Y(_00361_));
 XOR2x2_ASAP7_75t_R _16960_ (.A(_08752_),
    .B(_00911_),
    .Y(_08831_));
 AND2x2_ASAP7_75t_R _16961_ (.A(ld),
    .B(key[50]),
    .Y(_08832_));
 AO21x1_ASAP7_75t_R _16962_ (.A1(_08831_),
    .A2(_08005_),
    .B(_08832_),
    .Y(_00362_));
 XOR2x2_ASAP7_75t_R _16963_ (.A(_08754_),
    .B(_00912_),
    .Y(_08833_));
 AND2x2_ASAP7_75t_R _16964_ (.A(ld),
    .B(key[51]),
    .Y(_08834_));
 AO21x1_ASAP7_75t_R _16965_ (.A1(_08833_),
    .A2(_08005_),
    .B(_08834_),
    .Y(_00363_));
 XOR2x2_ASAP7_75t_R _16966_ (.A(_08756_),
    .B(_00914_),
    .Y(_08835_));
 AND2x2_ASAP7_75t_R _16967_ (.A(ld),
    .B(key[52]),
    .Y(_08836_));
 AO21x1_ASAP7_75t_R _16968_ (.A1(_08835_),
    .A2(_08005_),
    .B(_08836_),
    .Y(_00365_));
 XOR2x2_ASAP7_75t_R _16969_ (.A(_08759_),
    .B(_00915_),
    .Y(_08837_));
 AND2x2_ASAP7_75t_R _16970_ (.A(ld),
    .B(key[53]),
    .Y(_08838_));
 AO21x1_ASAP7_75t_R _16971_ (.A1(_08837_),
    .A2(_08005_),
    .B(_08838_),
    .Y(_00366_));
 XOR2x2_ASAP7_75t_R _16972_ (.A(_08761_),
    .B(_00916_),
    .Y(_08839_));
 AND2x2_ASAP7_75t_R _16973_ (.A(ld),
    .B(key[54]),
    .Y(_08840_));
 AO21x1_ASAP7_75t_R _16974_ (.A1(_08839_),
    .A2(_08005_),
    .B(_08840_),
    .Y(_00367_));
 XOR2x2_ASAP7_75t_R _16975_ (.A(_08764_),
    .B(_00917_),
    .Y(_08841_));
 AND2x2_ASAP7_75t_R _16976_ (.A(ld),
    .B(key[55]),
    .Y(_08842_));
 AO21x1_ASAP7_75t_R _16977_ (.A1(_08841_),
    .A2(_08005_),
    .B(_08842_),
    .Y(_00368_));
 INVx1_ASAP7_75t_R _16978_ (.A(_00918_),
    .Y(_08843_));
 OA21x2_ASAP7_75t_R _16979_ (.A1(_08766_),
    .A2(_08843_),
    .B(_08005_),
    .Y(_08844_));
 NAND2x1_ASAP7_75t_R _16980_ (.A(_08843_),
    .B(_08766_),
    .Y(_08845_));
 AO22x1_ASAP7_75t_R _16981_ (.A1(_08844_),
    .A2(_08845_),
    .B1(ld),
    .B2(key[56]),
    .Y(_00369_));
 XOR2x2_ASAP7_75t_R _16982_ (.A(_08769_),
    .B(_00919_),
    .Y(_08846_));
 AND2x2_ASAP7_75t_R _16983_ (.A(ld),
    .B(key[57]),
    .Y(_08847_));
 AO21x1_ASAP7_75t_R _16984_ (.A1(_08846_),
    .A2(_08005_),
    .B(_08847_),
    .Y(_00370_));
 INVx1_ASAP7_75t_R _16985_ (.A(_00920_),
    .Y(_08848_));
 OA21x2_ASAP7_75t_R _16986_ (.A1(_08771_),
    .A2(_08848_),
    .B(_08005_),
    .Y(_08849_));
 NAND2x1_ASAP7_75t_R _16987_ (.A(_08848_),
    .B(_08771_),
    .Y(_08850_));
 AO22x1_ASAP7_75t_R _16988_ (.A1(_08849_),
    .A2(_08850_),
    .B1(ld),
    .B2(key[58]),
    .Y(_00371_));
 INVx1_ASAP7_75t_R _16989_ (.A(_00921_),
    .Y(_08851_));
 OA21x2_ASAP7_75t_R _16990_ (.A1(_08773_),
    .A2(_08851_),
    .B(_08005_),
    .Y(_08852_));
 NAND2x1_ASAP7_75t_R _16991_ (.A(_08851_),
    .B(_08773_),
    .Y(_08853_));
 AO22x1_ASAP7_75t_R _16992_ (.A1(_08852_),
    .A2(_08853_),
    .B1(ld),
    .B2(key[59]),
    .Y(_00372_));
 XOR2x2_ASAP7_75t_R _16993_ (.A(_08776_),
    .B(_00922_),
    .Y(_08854_));
 AND2x2_ASAP7_75t_R _16994_ (.A(ld),
    .B(key[60]),
    .Y(_08855_));
 AO21x1_ASAP7_75t_R _16995_ (.A1(_08854_),
    .A2(_08005_),
    .B(_08855_),
    .Y(_00373_));
 XOR2x2_ASAP7_75t_R _16996_ (.A(_08779_),
    .B(_00923_),
    .Y(_08856_));
 AND2x2_ASAP7_75t_R _16997_ (.A(ld),
    .B(key[61]),
    .Y(_08857_));
 AO21x1_ASAP7_75t_R _16998_ (.A1(_08856_),
    .A2(_08005_),
    .B(_08857_),
    .Y(_00374_));
 XNOR2x2_ASAP7_75t_R _16999_ (.A(_00925_),
    .B(_08781_),
    .Y(_08858_));
 NOR2x1_ASAP7_75t_R _17000_ (.A(ld),
    .B(_08858_),
    .Y(_08859_));
 AO21x1_ASAP7_75t_R _17001_ (.A1(ld),
    .A2(key[62]),
    .B(_08859_),
    .Y(_00376_));
 XNOR2x2_ASAP7_75t_SL _17002_ (.A(_00926_),
    .B(_08783_),
    .Y(_08860_));
 NOR2x1_ASAP7_75t_R _17003_ (.A(ld),
    .B(_08860_),
    .Y(_08861_));
 AO21x1_ASAP7_75t_R _17004_ (.A1(ld),
    .A2(key[63]),
    .B(_08861_),
    .Y(_00377_));
 INVx1_ASAP7_75t_R _17005_ (.A(_00934_),
    .Y(_08862_));
 XOR2x2_ASAP7_75t_SL _17006_ (.A(_08785_),
    .B(_08862_),
    .Y(_08863_));
 NOR2x1_ASAP7_75t_R _17007_ (.A(key[0]),
    .B(_08005_),
    .Y(_08864_));
 INVx1_ASAP7_75t_R _17008_ (.A(_08864_),
    .Y(_08865_));
 OAI21x1_ASAP7_75t_R _17009_ (.A1(ld),
    .A2(_08863_),
    .B(_08865_),
    .Y(_08866_));
 INVx1_ASAP7_75t_R _17011_ (.A(_00945_),
    .Y(_08867_));
 XOR2x2_ASAP7_75t_SL _17012_ (.A(_08787_),
    .B(_08867_),
    .Y(_08868_));
 NOR2x1_ASAP7_75t_R _17013_ (.A(key[1]),
    .B(_08005_),
    .Y(_08869_));
 INVx1_ASAP7_75t_R _17014_ (.A(_08869_),
    .Y(_08870_));
 OAI21x1_ASAP7_75t_R _17015_ (.A1(ld),
    .A2(_08868_),
    .B(_08870_),
    .Y(_08871_));
 OR2x2_ASAP7_75t_SL _17017_ (.A(_08005_),
    .B(key[2]),
    .Y(_08872_));
 XOR2x1_ASAP7_75t_SL _17018_ (.A(_00924_),
    .Y(_08873_),
    .B(_00956_));
 XOR2x2_ASAP7_75t_SL _17019_ (.A(_08873_),
    .B(_00423_),
    .Y(_08874_));
 XOR2x2_ASAP7_75t_R _17020_ (.A(_00860_),
    .B(_00892_),
    .Y(_08875_));
 XOR2x2_ASAP7_75t_SL _17021_ (.A(_08874_),
    .B(_08875_),
    .Y(_08876_));
 NAND2x2_ASAP7_75t_SL _17022_ (.A(_08005_),
    .B(_08876_),
    .Y(_08877_));
 NAND2x2_ASAP7_75t_SL _17023_ (.A(_08872_),
    .B(_08877_),
    .Y(_08878_));
 INVx2_ASAP7_75t_SL _17024_ (.A(_08878_),
    .Y(_08879_));
 INVx1_ASAP7_75t_R _17026_ (.A(_00959_),
    .Y(_08880_));
 NOR2x1_ASAP7_75t_R _17027_ (.A(_08880_),
    .B(_08795_),
    .Y(_08881_));
 AND2x2_ASAP7_75t_SL _17028_ (.A(_08795_),
    .B(_08880_),
    .Y(_08882_));
 OAI21x1_ASAP7_75t_SL _17029_ (.A1(_08881_),
    .A2(_08882_),
    .B(_08005_),
    .Y(_08883_));
 OAI21x1_ASAP7_75t_SL _17030_ (.A1(_08005_),
    .A2(key[3]),
    .B(_08883_),
    .Y(_08884_));
 INVx2_ASAP7_75t_SL _17031_ (.A(_08884_),
    .Y(_08885_));
 XOR2x2_ASAP7_75t_R _17035_ (.A(_08797_),
    .B(_00960_),
    .Y(_08888_));
 NAND2x1_ASAP7_75t_R _17036_ (.A(ld),
    .B(key[4]),
    .Y(_08889_));
 OAI21x1_ASAP7_75t_SL _17037_ (.A1(ld),
    .A2(_08888_),
    .B(_08889_),
    .Y(_08890_));
 XOR2x2_ASAP7_75t_SL _17040_ (.A(_08800_),
    .B(_00961_),
    .Y(_08892_));
 NAND2x1_ASAP7_75t_R _17041_ (.A(ld),
    .B(key[5]),
    .Y(_08893_));
 OAI21x1_ASAP7_75t_R _17042_ (.A1(ld),
    .A2(_08892_),
    .B(_08893_),
    .Y(_08894_));
 XOR2x2_ASAP7_75t_SL _17045_ (.A(_08802_),
    .B(_00962_),
    .Y(_08896_));
 NAND2x1_ASAP7_75t_R _17046_ (.A(_08005_),
    .B(_08896_),
    .Y(_08897_));
 OAI21x1_ASAP7_75t_SL _17047_ (.A1(_08005_),
    .A2(key[6]),
    .B(_08897_),
    .Y(_08898_));
 INVx1_ASAP7_75t_SL _17048_ (.A(_08898_),
    .Y(_08899_));
 XOR2x2_ASAP7_75t_R _17050_ (.A(_08804_),
    .B(_00963_),
    .Y(_08900_));
 NAND2x1_ASAP7_75t_SL _17051_ (.A(_08005_),
    .B(_08900_),
    .Y(_08901_));
 OA21x2_ASAP7_75t_SL _17052_ (.A1(_08005_),
    .A2(key[7]),
    .B(_08901_),
    .Y(_08902_));
 INVx1_ASAP7_75t_R _17054_ (.A(_00964_),
    .Y(_08903_));
 XOR2x2_ASAP7_75t_SL _17055_ (.A(_08806_),
    .B(_08903_),
    .Y(_08904_));
 NOR2x1_ASAP7_75t_R _17056_ (.A(key[8]),
    .B(_08005_),
    .Y(_08905_));
 INVx1_ASAP7_75t_R _17057_ (.A(_08905_),
    .Y(_08906_));
 OAI21x1_ASAP7_75t_R _17058_ (.A1(ld),
    .A2(_08904_),
    .B(_08906_),
    .Y(_08907_));
 XOR2x2_ASAP7_75t_SL _17060_ (.A(_08808_),
    .B(_00430_),
    .Y(_08908_));
 XNOR2x2_ASAP7_75t_R _17061_ (.A(_00486_),
    .B(_00869_),
    .Y(_08909_));
 XOR2x2_ASAP7_75t_SL _17062_ (.A(_08908_),
    .B(_08909_),
    .Y(_08910_));
 OR2x2_ASAP7_75t_R _17063_ (.A(_08005_),
    .B(key[9]),
    .Y(_08911_));
 OAI21x1_ASAP7_75t_SL _17064_ (.A1(_08910_),
    .A2(ld),
    .B(_08911_),
    .Y(_01002_));
 OR2x2_ASAP7_75t_SL _17065_ (.A(_08005_),
    .B(key[10]),
    .Y(_08912_));
 XOR2x1_ASAP7_75t_SL _17066_ (.A(_00903_),
    .Y(_08913_),
    .B(_00935_));
 XOR2x2_ASAP7_75t_SL _17067_ (.A(_08913_),
    .B(_00431_),
    .Y(_08914_));
 XOR2x2_ASAP7_75t_SL _17068_ (.A(_00839_),
    .B(_00871_),
    .Y(_08915_));
 XOR2x1_ASAP7_75t_SL _17069_ (.A(_08914_),
    .Y(_08916_),
    .B(_08915_));
 NAND2x1_ASAP7_75t_SL _17070_ (.A(_08005_),
    .B(_08916_),
    .Y(_08917_));
 NAND2x1_ASAP7_75t_SL _17071_ (.A(_08912_),
    .B(_08917_),
    .Y(_08918_));
 INVx1_ASAP7_75t_SL _17072_ (.A(_08918_),
    .Y(_08919_));
 INVx1_ASAP7_75t_R _17074_ (.A(_00936_),
    .Y(_08920_));
 NOR2x1_ASAP7_75t_R _17075_ (.A(_08920_),
    .B(_08815_),
    .Y(_08921_));
 AND2x2_ASAP7_75t_R _17076_ (.A(_08815_),
    .B(_08920_),
    .Y(_08922_));
 OAI21x1_ASAP7_75t_SL _17077_ (.A1(_08921_),
    .A2(_08922_),
    .B(_08005_),
    .Y(_08923_));
 OAI21x1_ASAP7_75t_SL _17078_ (.A1(_08005_),
    .A2(key[11]),
    .B(_08923_),
    .Y(_08924_));
 INVx2_ASAP7_75t_SL _17079_ (.A(_08924_),
    .Y(_08925_));
 XOR2x2_ASAP7_75t_SL _17082_ (.A(_08817_),
    .B(_00937_),
    .Y(_08927_));
 NAND2x1_ASAP7_75t_R _17083_ (.A(ld),
    .B(key[12]),
    .Y(_08928_));
 OAI21x1_ASAP7_75t_R _17084_ (.A1(ld),
    .A2(_08927_),
    .B(_08928_),
    .Y(_08929_));
 XOR2x2_ASAP7_75t_R _17087_ (.A(_08819_),
    .B(_00938_),
    .Y(_08931_));
 NAND2x1_ASAP7_75t_R _17088_ (.A(_08005_),
    .B(_08931_),
    .Y(_08932_));
 OAI21x1_ASAP7_75t_SL _17089_ (.A1(_08005_),
    .A2(key[13]),
    .B(_08932_),
    .Y(_08933_));
 INVx2_ASAP7_75t_SL _17090_ (.A(_08933_),
    .Y(_08934_));
 XOR2x2_ASAP7_75t_R _17092_ (.A(_08822_),
    .B(_00939_),
    .Y(_08935_));
 NAND2x1_ASAP7_75t_SL _17093_ (.A(_08005_),
    .B(_08935_),
    .Y(_08936_));
 OAI21x1_ASAP7_75t_SL _17094_ (.A1(_08005_),
    .A2(key[14]),
    .B(_08936_),
    .Y(_08937_));
 INVx1_ASAP7_75t_SL _17095_ (.A(_08937_),
    .Y(_08938_));
 XOR2x2_ASAP7_75t_R _17097_ (.A(_08824_),
    .B(_00940_),
    .Y(_08939_));
 NAND2x1_ASAP7_75t_R _17098_ (.A(_08005_),
    .B(_08939_),
    .Y(_08940_));
 OA21x2_ASAP7_75t_SL _17099_ (.A1(_08005_),
    .A2(key[15]),
    .B(_08940_),
    .Y(_08941_));
 XOR2x2_ASAP7_75t_R _17101_ (.A(_00918_),
    .B(_00950_),
    .Y(_08942_));
 AOI21x1_ASAP7_75t_R _17102_ (.A1(_08942_),
    .A2(_08766_),
    .B(ld),
    .Y(_08943_));
 NOR2x1_ASAP7_75t_SL _17103_ (.A(_08942_),
    .B(_08766_),
    .Y(_08944_));
 INVx1_ASAP7_75t_R _17104_ (.A(_08944_),
    .Y(_08945_));
 AND2x2_ASAP7_75t_R _17105_ (.A(ld),
    .B(key[24]),
    .Y(_08946_));
 AOI21x1_ASAP7_75t_SL _17106_ (.A1(_08945_),
    .A2(_08943_),
    .B(_08946_),
    .Y(_01043_));
 XNOR2x2_ASAP7_75t_R _17107_ (.A(_00919_),
    .B(_00951_),
    .Y(_08947_));
 XOR2x2_ASAP7_75t_SL _17108_ (.A(_08769_),
    .B(_08947_),
    .Y(_08948_));
 NOR2x1_ASAP7_75t_R _17109_ (.A(key[25]),
    .B(_08005_),
    .Y(_08949_));
 INVx1_ASAP7_75t_R _17110_ (.A(_08949_),
    .Y(_08950_));
 OAI21x1_ASAP7_75t_SL _17111_ (.A1(_08948_),
    .A2(ld),
    .B(_08950_),
    .Y(_01046_));
 XOR2x2_ASAP7_75t_R _17112_ (.A(_00920_),
    .B(_00952_),
    .Y(_08951_));
 INVx1_ASAP7_75t_R _17113_ (.A(_08951_),
    .Y(_08952_));
 INVx1_ASAP7_75t_SL _17114_ (.A(_00888_),
    .Y(_08953_));
 XOR2x2_ASAP7_75t_SL _17115_ (.A(_08690_),
    .B(_08953_),
    .Y(_08954_));
 NAND2x1_ASAP7_75t_SL _17116_ (.A(_08952_),
    .B(_08954_),
    .Y(_08955_));
 AOI21x1_ASAP7_75t_L _17117_ (.A1(_08951_),
    .A2(_08771_),
    .B(ld),
    .Y(_08956_));
 AND2x2_ASAP7_75t_R _17118_ (.A(ld),
    .B(key[26]),
    .Y(_08957_));
 AOI21x1_ASAP7_75t_SL _17119_ (.A1(_08955_),
    .A2(_08956_),
    .B(_08957_),
    .Y(_08958_));
 XOR2x2_ASAP7_75t_R _17122_ (.A(_00921_),
    .B(_00953_),
    .Y(_08960_));
 NOR2x1_ASAP7_75t_R _17123_ (.A(_08960_),
    .B(_08773_),
    .Y(_08961_));
 INVx1_ASAP7_75t_R _17124_ (.A(_08960_),
    .Y(_08962_));
 INVx1_ASAP7_75t_R _17125_ (.A(_00889_),
    .Y(_08963_));
 XOR2x2_ASAP7_75t_R _17126_ (.A(_08693_),
    .B(_08963_),
    .Y(_08964_));
 OAI21x1_ASAP7_75t_R _17127_ (.A1(_08962_),
    .A2(_08964_),
    .B(_08005_),
    .Y(_08965_));
 AND2x2_ASAP7_75t_R _17128_ (.A(ld),
    .B(key[27]),
    .Y(_08966_));
 INVx1_ASAP7_75t_R _17129_ (.A(_08966_),
    .Y(_08967_));
 OAI21x1_ASAP7_75t_SL _17130_ (.A1(_08961_),
    .A2(_08965_),
    .B(_08967_),
    .Y(_08968_));
 XNOR2x2_ASAP7_75t_R _17134_ (.A(_00922_),
    .B(_00954_),
    .Y(_08971_));
 XOR2x2_ASAP7_75t_SL _17135_ (.A(_08776_),
    .B(_08971_),
    .Y(_08972_));
 NOR2x1_ASAP7_75t_R _17136_ (.A(key[28]),
    .B(_08005_),
    .Y(_08973_));
 INVx1_ASAP7_75t_R _17137_ (.A(_08973_),
    .Y(_08974_));
 OAI21x1_ASAP7_75t_R _17138_ (.A1(ld),
    .A2(_08972_),
    .B(_08974_),
    .Y(_08975_));
 INVx1_ASAP7_75t_SL _17139_ (.A(_08975_),
    .Y(_08976_));
 XNOR2x2_ASAP7_75t_R _17142_ (.A(_00923_),
    .B(_00955_),
    .Y(_08978_));
 XOR2x2_ASAP7_75t_R _17143_ (.A(_08779_),
    .B(_08978_),
    .Y(_08979_));
 NOR2x1_ASAP7_75t_R _17144_ (.A(key[29]),
    .B(_08005_),
    .Y(_08980_));
 INVx1_ASAP7_75t_R _17145_ (.A(_08980_),
    .Y(_08981_));
 OA21x2_ASAP7_75t_SL _17146_ (.A1(_08979_),
    .A2(ld),
    .B(_08981_),
    .Y(_08982_));
 XOR2x2_ASAP7_75t_SL _17149_ (.A(_08858_),
    .B(_00957_),
    .Y(_08984_));
 NOR2x1_ASAP7_75t_R _17150_ (.A(key[30]),
    .B(_08005_),
    .Y(_08985_));
 INVx1_ASAP7_75t_R _17151_ (.A(_08985_),
    .Y(_08986_));
 OAI21x1_ASAP7_75t_R _17152_ (.A1(ld),
    .A2(_08984_),
    .B(_08986_),
    .Y(_08987_));
 INVx1_ASAP7_75t_SL _17153_ (.A(_08987_),
    .Y(_08988_));
 XOR2x2_ASAP7_75t_R _17155_ (.A(_08860_),
    .B(_00958_),
    .Y(_08989_));
 NOR2x1_ASAP7_75t_R _17156_ (.A(key[31]),
    .B(_08005_),
    .Y(_08990_));
 INVx1_ASAP7_75t_R _17157_ (.A(_08990_),
    .Y(_08991_));
 OA21x2_ASAP7_75t_SL _17158_ (.A1(_08989_),
    .A2(ld),
    .B(_08991_),
    .Y(_08992_));
 INVx4_ASAP7_75t_SL _17160_ (.A(_01002_),
    .Y(_00994_));
 XOR2x2_ASAP7_75t_SL _17163_ (.A(_08806_),
    .B(_00964_),
    .Y(_08994_));
 AOI21x1_ASAP7_75t_R _17164_ (.A1(_08005_),
    .A2(_08994_),
    .B(_08905_),
    .Y(_08995_));
 NAND2x1_ASAP7_75t_SL _17167_ (.A(_01003_),
    .B(_08919_),
    .Y(_08997_));
 INVx1_ASAP7_75t_SL _17170_ (.A(_01005_),
    .Y(_09000_));
 AO21x1_ASAP7_75t_SL _17171_ (.A1(_08917_),
    .A2(_08912_),
    .B(_09000_),
    .Y(_09001_));
 AO21x1_ASAP7_75t_SL _17174_ (.A1(_08997_),
    .A2(_09001_),
    .B(_08924_),
    .Y(_09004_));
 INVx2_ASAP7_75t_R _17176_ (.A(_00996_),
    .Y(_09006_));
 AND2x2_ASAP7_75t_SL _17177_ (.A(_08918_),
    .B(_09006_),
    .Y(_09007_));
 INVx1_ASAP7_75t_SL _17178_ (.A(_09007_),
    .Y(_09008_));
 INVx1_ASAP7_75t_SL _17179_ (.A(_00997_),
    .Y(_09009_));
 NOR2x1p5_ASAP7_75t_SL _17180_ (.A(_09009_),
    .B(_08918_),
    .Y(_09010_));
 NOR2x1p5_ASAP7_75t_SL _17181_ (.A(_09010_),
    .B(_08925_),
    .Y(_09011_));
 AOI21x1_ASAP7_75t_SL _17182_ (.A1(_09008_),
    .A2(_09011_),
    .B(_08929_),
    .Y(_09012_));
 NAND2x1_ASAP7_75t_SL _17183_ (.A(_00994_),
    .B(_08907_),
    .Y(_09013_));
 NAND2x1_ASAP7_75t_SL _17184_ (.A(_08918_),
    .B(_08995_),
    .Y(_09014_));
 AOI21x1_ASAP7_75t_SL _17185_ (.A1(_09013_),
    .A2(_09014_),
    .B(_08925_),
    .Y(_09015_));
 INVx1_ASAP7_75t_SL _17186_ (.A(_09015_),
    .Y(_09016_));
 NAND2x1_ASAP7_75t_SL _17187_ (.A(_01002_),
    .B(_08907_),
    .Y(_09017_));
 NAND2x1_ASAP7_75t_SL _17188_ (.A(_08919_),
    .B(_08995_),
    .Y(_09018_));
 NAND2x1_ASAP7_75t_SL _17189_ (.A(_09017_),
    .B(_09018_),
    .Y(_09019_));
 INVx1_ASAP7_75t_SL _17190_ (.A(_08929_),
    .Y(_09020_));
 AOI21x1_ASAP7_75t_SL _17193_ (.A1(_08925_),
    .A2(_09019_),
    .B(_09020_),
    .Y(_09023_));
 AOI221x1_ASAP7_75t_SL _17194_ (.A1(_09004_),
    .A2(_09012_),
    .B1(_09016_),
    .B2(_09023_),
    .C(_08938_),
    .Y(_09024_));
 INVx1_ASAP7_75t_SL _17195_ (.A(_08941_),
    .Y(_09025_));
 NOR2x1p5_ASAP7_75t_SL _17196_ (.A(_08924_),
    .B(_09010_),
    .Y(_09026_));
 INVx1_ASAP7_75t_SL _17197_ (.A(_00998_),
    .Y(_09027_));
 AO21x2_ASAP7_75t_R _17198_ (.A1(_08917_),
    .A2(_08912_),
    .B(_09027_),
    .Y(_09028_));
 AND2x2_ASAP7_75t_SL _17199_ (.A(_09028_),
    .B(_09026_),
    .Y(_09029_));
 NAND2x1_ASAP7_75t_SL _17200_ (.A(_08919_),
    .B(_08907_),
    .Y(_09030_));
 INVx1_ASAP7_75t_SL _17201_ (.A(_01000_),
    .Y(_09031_));
 AND2x2_ASAP7_75t_R _17202_ (.A(_08918_),
    .B(_09031_),
    .Y(_09032_));
 NOR2x1_ASAP7_75t_L _17203_ (.A(_08925_),
    .B(_09032_),
    .Y(_09033_));
 NAND2x1_ASAP7_75t_R _17204_ (.A(_09030_),
    .B(_09033_),
    .Y(_09034_));
 INVx1_ASAP7_75t_SL _17205_ (.A(_09034_),
    .Y(_09035_));
 OAI21x1_ASAP7_75t_SL _17207_ (.A1(_09029_),
    .A2(_09035_),
    .B(_08929_),
    .Y(_09037_));
 AOI21x1_ASAP7_75t_SL _17209_ (.A1(_08918_),
    .A2(_08907_),
    .B(_08925_),
    .Y(_09039_));
 AO21x1_ASAP7_75t_R _17211_ (.A1(_08919_),
    .A2(_01001_),
    .B(_08924_),
    .Y(_09041_));
 NOR2x1_ASAP7_75t_SL _17212_ (.A(_09032_),
    .B(_09041_),
    .Y(_09042_));
 OAI21x1_ASAP7_75t_SL _17214_ (.A1(_09039_),
    .A2(_09042_),
    .B(_09020_),
    .Y(_09044_));
 AO21x1_ASAP7_75t_SL _17216_ (.A1(_09044_),
    .A2(_09037_),
    .B(_08937_),
    .Y(_09046_));
 NAND2x1_ASAP7_75t_SL _17217_ (.A(_09046_),
    .B(_09025_),
    .Y(_09047_));
 NOR2x1_ASAP7_75t_SL _17218_ (.A(_01006_),
    .B(_08918_),
    .Y(_09048_));
 INVx1_ASAP7_75t_SL _17219_ (.A(_09048_),
    .Y(_09049_));
 AO21x1_ASAP7_75t_SL _17221_ (.A1(_09049_),
    .A2(_09001_),
    .B(_08925_),
    .Y(_09051_));
 AND2x2_ASAP7_75t_SL _17223_ (.A(_09041_),
    .B(_08929_),
    .Y(_09053_));
 AOI21x1_ASAP7_75t_SL _17224_ (.A1(_09051_),
    .A2(_09053_),
    .B(_08937_),
    .Y(_09054_));
 NAND2x1_ASAP7_75t_SL _17225_ (.A(_00994_),
    .B(_08919_),
    .Y(_09055_));
 AO21x1_ASAP7_75t_SL _17226_ (.A1(_08917_),
    .A2(_08912_),
    .B(_00997_),
    .Y(_09056_));
 AO21x1_ASAP7_75t_R _17228_ (.A1(_09055_),
    .A2(_09056_),
    .B(_08925_),
    .Y(_09058_));
 INVx1_ASAP7_75t_SL _17229_ (.A(_09058_),
    .Y(_09059_));
 INVx1_ASAP7_75t_R _17230_ (.A(_01003_),
    .Y(_09060_));
 AO21x2_ASAP7_75t_SL _17231_ (.A1(_08917_),
    .A2(_08912_),
    .B(_09060_),
    .Y(_09061_));
 INVx1_ASAP7_75t_SL _17232_ (.A(_09061_),
    .Y(_09062_));
 OAI21x1_ASAP7_75t_SL _17234_ (.A1(_08918_),
    .A2(_08907_),
    .B(_08925_),
    .Y(_09064_));
 NOR2x1_ASAP7_75t_SL _17235_ (.A(_09062_),
    .B(_09064_),
    .Y(_09065_));
 OAI21x1_ASAP7_75t_SL _17237_ (.A1(_09059_),
    .A2(_09065_),
    .B(_09020_),
    .Y(_09067_));
 AOI21x1_ASAP7_75t_SL _17238_ (.A1(_09054_),
    .A2(_09067_),
    .B(_09025_),
    .Y(_09068_));
 NOR2x1_ASAP7_75t_L _17239_ (.A(_08925_),
    .B(_09061_),
    .Y(_09069_));
 NAND2x1_ASAP7_75t_SL _17240_ (.A(_08925_),
    .B(_09048_),
    .Y(_09070_));
 INVx1_ASAP7_75t_SL _17241_ (.A(_09070_),
    .Y(_09071_));
 NOR2x1_ASAP7_75t_SL _17242_ (.A(_09069_),
    .B(_09071_),
    .Y(_09072_));
 NOR2x1_ASAP7_75t_R _17243_ (.A(_09031_),
    .B(_08918_),
    .Y(_09073_));
 INVx1_ASAP7_75t_R _17244_ (.A(_09073_),
    .Y(_09074_));
 OA21x2_ASAP7_75t_SL _17245_ (.A1(_09074_),
    .A2(_08925_),
    .B(_08929_),
    .Y(_09075_));
 AOI21x1_ASAP7_75t_SL _17246_ (.A1(_09072_),
    .A2(_09075_),
    .B(_08938_),
    .Y(_09076_));
 AO21x1_ASAP7_75t_SL _17247_ (.A1(_08919_),
    .A2(_09031_),
    .B(_08924_),
    .Y(_09077_));
 AND2x2_ASAP7_75t_R _17248_ (.A(_08918_),
    .B(_01004_),
    .Y(_09078_));
 OA21x2_ASAP7_75t_SL _17249_ (.A1(_09077_),
    .A2(_09078_),
    .B(_09020_),
    .Y(_09079_));
 OAI21x1_ASAP7_75t_SL _17250_ (.A1(_08925_),
    .A2(_09049_),
    .B(_09079_),
    .Y(_09080_));
 NAND2x1_ASAP7_75t_SL _17251_ (.A(_09076_),
    .B(_09080_),
    .Y(_09081_));
 AOI21x1_ASAP7_75t_SL _17254_ (.A1(_09068_),
    .A2(_09081_),
    .B(_08933_),
    .Y(_09084_));
 OAI21x1_ASAP7_75t_SL _17255_ (.A1(_09047_),
    .A2(_09024_),
    .B(_09084_),
    .Y(_09085_));
 NOR2x1_ASAP7_75t_R _17257_ (.A(_01000_),
    .B(_08918_),
    .Y(_09087_));
 INVx1_ASAP7_75t_R _17258_ (.A(_09087_),
    .Y(_09088_));
 AOI21x1_ASAP7_75t_R _17259_ (.A1(_08918_),
    .A2(_08995_),
    .B(_08925_),
    .Y(_09089_));
 NAND2x1_ASAP7_75t_SL _17260_ (.A(_09088_),
    .B(_09089_),
    .Y(_09090_));
 OAI21x1_ASAP7_75t_R _17261_ (.A1(_08919_),
    .A2(_08995_),
    .B(_08925_),
    .Y(_09091_));
 NOR2x1_ASAP7_75t_R _17262_ (.A(_01005_),
    .B(_08918_),
    .Y(_09092_));
 OA21x2_ASAP7_75t_SL _17263_ (.A1(_09091_),
    .A2(_09092_),
    .B(_09020_),
    .Y(_09093_));
 AND2x4_ASAP7_75t_L _17264_ (.A(_09056_),
    .B(_08924_),
    .Y(_09094_));
 INVx1_ASAP7_75t_SL _17265_ (.A(_01013_),
    .Y(_09095_));
 NOR2x1_ASAP7_75t_R _17266_ (.A(_09095_),
    .B(_08924_),
    .Y(_09096_));
 OA21x2_ASAP7_75t_SL _17267_ (.A1(_09094_),
    .A2(_09096_),
    .B(_08929_),
    .Y(_09097_));
 AOI21x1_ASAP7_75t_SL _17268_ (.A1(_09090_),
    .A2(_09093_),
    .B(_09097_),
    .Y(_09098_));
 INVx2_ASAP7_75t_SL _17269_ (.A(_09026_),
    .Y(_09099_));
 NOR2x1_ASAP7_75t_R _17270_ (.A(_01004_),
    .B(_08918_),
    .Y(_09100_));
 NAND2x1_ASAP7_75t_SL _17271_ (.A(_08924_),
    .B(_09100_),
    .Y(_09101_));
 AND2x2_ASAP7_75t_R _17272_ (.A(_09101_),
    .B(_08929_),
    .Y(_09102_));
 NAND2x1_ASAP7_75t_SL _17273_ (.A(_09099_),
    .B(_09102_),
    .Y(_09103_));
 NOR2x1_ASAP7_75t_R _17274_ (.A(_00996_),
    .B(_08918_),
    .Y(_09104_));
 OAI21x1_ASAP7_75t_SL _17275_ (.A1(_09104_),
    .A2(_09091_),
    .B(_09020_),
    .Y(_09105_));
 AO21x1_ASAP7_75t_SL _17277_ (.A1(_08917_),
    .A2(_08912_),
    .B(_01001_),
    .Y(_09107_));
 INVx1_ASAP7_75t_R _17278_ (.A(_09107_),
    .Y(_09108_));
 AO21x1_ASAP7_75t_SL _17279_ (.A1(_08924_),
    .A2(_09108_),
    .B(_08937_),
    .Y(_09109_));
 AO21x1_ASAP7_75t_SL _17280_ (.A1(_09103_),
    .A2(_09105_),
    .B(_09109_),
    .Y(_09110_));
 OA21x2_ASAP7_75t_SL _17281_ (.A1(_09098_),
    .A2(_08938_),
    .B(_09110_),
    .Y(_09111_));
 NAND2x1_ASAP7_75t_SL _17283_ (.A(_01002_),
    .B(_08918_),
    .Y(_09113_));
 NOR2x1_ASAP7_75t_SL _17284_ (.A(_08925_),
    .B(_09113_),
    .Y(_09114_));
 AOI211x1_ASAP7_75t_R _17285_ (.A1(_08924_),
    .A2(_09048_),
    .B(_09114_),
    .C(_08929_),
    .Y(_09115_));
 NOR2x1_ASAP7_75t_SL _17286_ (.A(_09006_),
    .B(_08918_),
    .Y(_09116_));
 INVx2_ASAP7_75t_SL _17287_ (.A(_09116_),
    .Y(_09117_));
 AO21x1_ASAP7_75t_R _17288_ (.A1(_09014_),
    .A2(_09117_),
    .B(_08924_),
    .Y(_09118_));
 AOI21x1_ASAP7_75t_SL _17289_ (.A1(_09115_),
    .A2(_09118_),
    .B(_08937_),
    .Y(_09119_));
 NOR2x1_ASAP7_75t_R _17290_ (.A(_09027_),
    .B(_08918_),
    .Y(_09120_));
 NAND2x1_ASAP7_75t_SL _17291_ (.A(_01002_),
    .B(_08919_),
    .Y(_09121_));
 NAND2x1_ASAP7_75t_R _17292_ (.A(_08924_),
    .B(_09121_),
    .Y(_09122_));
 OA21x2_ASAP7_75t_SL _17293_ (.A1(_09122_),
    .A2(_09032_),
    .B(_08929_),
    .Y(_09123_));
 OAI21x1_ASAP7_75t_SL _17294_ (.A1(_09091_),
    .A2(_09120_),
    .B(_09123_),
    .Y(_09124_));
 NAND2x1_ASAP7_75t_SL _17295_ (.A(_09119_),
    .B(_09124_),
    .Y(_09125_));
 NOR2x1_ASAP7_75t_SL _17296_ (.A(_08918_),
    .B(_00997_),
    .Y(_09126_));
 INVx2_ASAP7_75t_SL _17297_ (.A(_09126_),
    .Y(_09127_));
 AO21x1_ASAP7_75t_R _17298_ (.A1(_09127_),
    .A2(_09001_),
    .B(_08924_),
    .Y(_09128_));
 NOR2x1_ASAP7_75t_R _17299_ (.A(_09000_),
    .B(_08918_),
    .Y(_09129_));
 AO21x1_ASAP7_75t_R _17300_ (.A1(_08924_),
    .A2(_09129_),
    .B(_08929_),
    .Y(_09130_));
 NOR2x1_ASAP7_75t_R _17301_ (.A(_09069_),
    .B(_09130_),
    .Y(_09131_));
 NAND2x1_ASAP7_75t_SL _17302_ (.A(_09128_),
    .B(_09131_),
    .Y(_09132_));
 AND2x2_ASAP7_75t_L _17303_ (.A(_09011_),
    .B(_09113_),
    .Y(_09133_));
 AO21x2_ASAP7_75t_SL _17304_ (.A1(_08917_),
    .A2(_08912_),
    .B(_09009_),
    .Y(_09134_));
 INVx2_ASAP7_75t_SL _17305_ (.A(_09134_),
    .Y(_09135_));
 NAND2x1p5_ASAP7_75t_SL _17306_ (.A(_09135_),
    .B(_08925_),
    .Y(_09136_));
 NAND2x1_ASAP7_75t_SL _17307_ (.A(_09136_),
    .B(_08929_),
    .Y(_09137_));
 OA21x2_ASAP7_75t_SL _17308_ (.A1(_09137_),
    .A2(_09133_),
    .B(_08937_),
    .Y(_09138_));
 AOI21x1_ASAP7_75t_SL _17309_ (.A1(_09132_),
    .A2(_09138_),
    .B(_08941_),
    .Y(_09139_));
 AOI21x1_ASAP7_75t_SL _17310_ (.A1(_09139_),
    .A2(_09125_),
    .B(_08934_),
    .Y(_09140_));
 OAI21x1_ASAP7_75t_SL _17311_ (.A1(_09025_),
    .A2(_09111_),
    .B(_09140_),
    .Y(_09141_));
 NAND2x1_ASAP7_75t_SL _17312_ (.A(_09141_),
    .B(_09085_),
    .Y(_00008_));
 AND2x2_ASAP7_75t_SL _17313_ (.A(_09107_),
    .B(_09026_),
    .Y(_09142_));
 OAI21x1_ASAP7_75t_SL _17315_ (.A1(_08919_),
    .A2(_08907_),
    .B(_08924_),
    .Y(_09144_));
 OAI21x1_ASAP7_75t_SL _17317_ (.A1(_09129_),
    .A2(_09144_),
    .B(_08929_),
    .Y(_09146_));
 NOR2x1_ASAP7_75t_SL _17318_ (.A(_09142_),
    .B(_09146_),
    .Y(_09147_));
 NAND2x1_ASAP7_75t_SL _17319_ (.A(_09094_),
    .B(_09030_),
    .Y(_09148_));
 NOR2x1_ASAP7_75t_SL _17320_ (.A(_01002_),
    .B(_08907_),
    .Y(_09149_));
 NOR2x1_ASAP7_75t_SL _17321_ (.A(_08918_),
    .B(_08995_),
    .Y(_09150_));
 OAI21x1_ASAP7_75t_SL _17322_ (.A1(_09149_),
    .A2(_09150_),
    .B(_08925_),
    .Y(_09151_));
 AOI21x1_ASAP7_75t_SL _17323_ (.A1(_09148_),
    .A2(_09151_),
    .B(_08929_),
    .Y(_09152_));
 OAI21x1_ASAP7_75t_SL _17324_ (.A1(_09147_),
    .A2(_09152_),
    .B(_08933_),
    .Y(_09153_));
 INVx3_ASAP7_75t_SL _17325_ (.A(_09010_),
    .Y(_09154_));
 AO21x1_ASAP7_75t_R _17326_ (.A1(_08917_),
    .A2(_08912_),
    .B(_09006_),
    .Y(_09155_));
 AO21x1_ASAP7_75t_SL _17328_ (.A1(_09155_),
    .A2(_09154_),
    .B(_08924_),
    .Y(_09157_));
 INVx1_ASAP7_75t_SL _17330_ (.A(_01001_),
    .Y(_09159_));
 NAND2x1_ASAP7_75t_R _17331_ (.A(_09159_),
    .B(_08919_),
    .Y(_09160_));
 OA21x2_ASAP7_75t_SL _17332_ (.A1(_08925_),
    .A2(_09160_),
    .B(_09020_),
    .Y(_09161_));
 AOI21x1_ASAP7_75t_SL _17334_ (.A1(_09157_),
    .A2(_09161_),
    .B(_08933_),
    .Y(_09163_));
 AND2x2_ASAP7_75t_R _17335_ (.A(_09028_),
    .B(_08925_),
    .Y(_09164_));
 AOI21x1_ASAP7_75t_SL _17336_ (.A1(_09121_),
    .A2(_09164_),
    .B(_09020_),
    .Y(_09165_));
 OAI21x1_ASAP7_75t_SL _17337_ (.A1(_08925_),
    .A2(_09117_),
    .B(_09165_),
    .Y(_09166_));
 NAND2x1_ASAP7_75t_SL _17338_ (.A(_09163_),
    .B(_09166_),
    .Y(_09167_));
 AO21x1_ASAP7_75t_SL _17340_ (.A1(_09167_),
    .A2(_09153_),
    .B(_08937_),
    .Y(_09169_));
 OA21x2_ASAP7_75t_SL _17341_ (.A1(_08925_),
    .A2(_09107_),
    .B(_08929_),
    .Y(_09170_));
 NAND2x1_ASAP7_75t_R _17342_ (.A(_01008_),
    .B(_08925_),
    .Y(_09171_));
 OA21x2_ASAP7_75t_SL _17343_ (.A1(_09121_),
    .A2(_08925_),
    .B(_09171_),
    .Y(_09172_));
 AOI21x1_ASAP7_75t_SL _17345_ (.A1(_09170_),
    .A2(_09172_),
    .B(_08934_),
    .Y(_09174_));
 NAND2x1_ASAP7_75t_SL _17346_ (.A(_09027_),
    .B(_08919_),
    .Y(_09175_));
 AO21x1_ASAP7_75t_SL _17347_ (.A1(_09175_),
    .A2(_09056_),
    .B(_08924_),
    .Y(_09176_));
 NOR2x1_ASAP7_75t_SL _17348_ (.A(_09073_),
    .B(_09108_),
    .Y(_09177_));
 OA21x2_ASAP7_75t_SL _17349_ (.A1(_09177_),
    .A2(_08925_),
    .B(_09020_),
    .Y(_09178_));
 NAND2x1_ASAP7_75t_SL _17350_ (.A(_09176_),
    .B(_09178_),
    .Y(_09179_));
 NAND2x1_ASAP7_75t_SL _17351_ (.A(_09174_),
    .B(_09179_),
    .Y(_09180_));
 NAND2x1_ASAP7_75t_SL _17352_ (.A(_01001_),
    .B(_08919_),
    .Y(_09181_));
 AOI21x1_ASAP7_75t_SL _17353_ (.A1(_09181_),
    .A2(_09089_),
    .B(_09020_),
    .Y(_09182_));
 OAI21x1_ASAP7_75t_SL _17354_ (.A1(_09010_),
    .A2(_09091_),
    .B(_09182_),
    .Y(_09183_));
 AO21x1_ASAP7_75t_SL _17355_ (.A1(_08917_),
    .A2(_08912_),
    .B(_09031_),
    .Y(_09184_));
 OA21x2_ASAP7_75t_SL _17357_ (.A1(_08924_),
    .A2(_09184_),
    .B(_09020_),
    .Y(_09186_));
 NAND2x1_ASAP7_75t_R _17358_ (.A(_01002_),
    .B(_08995_),
    .Y(_09187_));
 NAND2x1_ASAP7_75t_SL _17359_ (.A(_00994_),
    .B(_08918_),
    .Y(_09188_));
 AO21x1_ASAP7_75t_SL _17360_ (.A1(_09187_),
    .A2(_09188_),
    .B(_08925_),
    .Y(_09189_));
 AOI21x1_ASAP7_75t_SL _17361_ (.A1(_09186_),
    .A2(_09189_),
    .B(_08933_),
    .Y(_09190_));
 NAND2x1_ASAP7_75t_SL _17362_ (.A(_09183_),
    .B(_09190_),
    .Y(_09191_));
 AOI21x1_ASAP7_75t_SL _17363_ (.A1(_09180_),
    .A2(_09191_),
    .B(_08938_),
    .Y(_09192_));
 NOR2x1_ASAP7_75t_SL _17364_ (.A(_09025_),
    .B(_09192_),
    .Y(_09193_));
 AO21x1_ASAP7_75t_SL _17365_ (.A1(_09160_),
    .A2(_09188_),
    .B(_08924_),
    .Y(_09194_));
 NAND2x1_ASAP7_75t_SL _17366_ (.A(_08929_),
    .B(_09194_),
    .Y(_09195_));
 INVx1_ASAP7_75t_SL _17367_ (.A(_09113_),
    .Y(_09196_));
 NOR2x1_ASAP7_75t_SL _17368_ (.A(_09196_),
    .B(_09150_),
    .Y(_09197_));
 OAI21x1_ASAP7_75t_SL _17369_ (.A1(_08925_),
    .A2(_09197_),
    .B(_08933_),
    .Y(_09198_));
 NOR2x1_ASAP7_75t_SL _17370_ (.A(_09195_),
    .B(_09198_),
    .Y(_09199_));
 AO21x1_ASAP7_75t_SL _17371_ (.A1(_09117_),
    .A2(_09184_),
    .B(_08924_),
    .Y(_09200_));
 OA21x2_ASAP7_75t_R _17372_ (.A1(_08919_),
    .A2(_01005_),
    .B(_08924_),
    .Y(_09201_));
 NAND2x1_ASAP7_75t_SL _17373_ (.A(_09030_),
    .B(_09201_),
    .Y(_09202_));
 AOI21x1_ASAP7_75t_SL _17375_ (.A1(_09200_),
    .A2(_09202_),
    .B(_09020_),
    .Y(_09204_));
 AO21x1_ASAP7_75t_SL _17377_ (.A1(_09117_),
    .A2(_09061_),
    .B(_08925_),
    .Y(_09206_));
 AND2x2_ASAP7_75t_R _17378_ (.A(_08925_),
    .B(_01014_),
    .Y(_09207_));
 OAI21x1_ASAP7_75t_SL _17379_ (.A1(_08929_),
    .A2(_09207_),
    .B(_08933_),
    .Y(_09208_));
 OAI21x1_ASAP7_75t_SL _17380_ (.A1(_08929_),
    .A2(_09206_),
    .B(_09208_),
    .Y(_09209_));
 NOR2x1_ASAP7_75t_SL _17381_ (.A(_09204_),
    .B(_09209_),
    .Y(_09210_));
 OAI21x1_ASAP7_75t_SL _17382_ (.A1(_09199_),
    .A2(_09210_),
    .B(_08937_),
    .Y(_09211_));
 INVx1_ASAP7_75t_SL _17383_ (.A(_09120_),
    .Y(_09212_));
 AOI21x1_ASAP7_75t_R _17384_ (.A1(_01006_),
    .A2(_08918_),
    .B(_08925_),
    .Y(_09213_));
 NAND2x1_ASAP7_75t_SL _17385_ (.A(_09212_),
    .B(_09213_),
    .Y(_09214_));
 NAND3x1_ASAP7_75t_SL _17386_ (.A(_09157_),
    .B(_09214_),
    .C(_08929_),
    .Y(_09215_));
 NOR2x1p5_ASAP7_75t_SL _17387_ (.A(_08929_),
    .B(_09026_),
    .Y(_09216_));
 NOR2x1_ASAP7_75t_SL _17388_ (.A(_08919_),
    .B(_08907_),
    .Y(_09217_));
 OAI21x1_ASAP7_75t_SL _17389_ (.A1(_09116_),
    .A2(_09217_),
    .B(_08924_),
    .Y(_09218_));
 AOI21x1_ASAP7_75t_SL _17390_ (.A1(_09218_),
    .A2(_09216_),
    .B(_08934_),
    .Y(_09219_));
 AOI21x1_ASAP7_75t_SL _17391_ (.A1(_09215_),
    .A2(_09219_),
    .B(_08937_),
    .Y(_09220_));
 NAND2x1_ASAP7_75t_R _17392_ (.A(_01005_),
    .B(_08919_),
    .Y(_09221_));
 AO21x1_ASAP7_75t_SL _17393_ (.A1(_09221_),
    .A2(_09056_),
    .B(_08924_),
    .Y(_09222_));
 OAI21x1_ASAP7_75t_SL _17394_ (.A1(_09048_),
    .A2(_09217_),
    .B(_08924_),
    .Y(_09223_));
 AOI21x1_ASAP7_75t_SL _17395_ (.A1(_09222_),
    .A2(_09223_),
    .B(_09020_),
    .Y(_09224_));
 INVx1_ASAP7_75t_R _17396_ (.A(_09001_),
    .Y(_09225_));
 OAI21x1_ASAP7_75t_SL _17397_ (.A1(_09225_),
    .A2(_09150_),
    .B(_08924_),
    .Y(_09226_));
 AOI21x1_ASAP7_75t_SL _17398_ (.A1(_09194_),
    .A2(_09226_),
    .B(_08929_),
    .Y(_09227_));
 OAI21x1_ASAP7_75t_SL _17399_ (.A1(_09224_),
    .A2(_09227_),
    .B(_08934_),
    .Y(_09228_));
 NAND2x1_ASAP7_75t_SL _17400_ (.A(_09228_),
    .B(_09220_),
    .Y(_09229_));
 AOI21x1_ASAP7_75t_SL _17401_ (.A1(_09211_),
    .A2(_09229_),
    .B(_08941_),
    .Y(_09230_));
 AOI21x1_ASAP7_75t_SL _17402_ (.A1(_09169_),
    .A2(_09193_),
    .B(_09230_),
    .Y(_00009_));
 AND3x1_ASAP7_75t_SL _17403_ (.A(_08924_),
    .B(_09127_),
    .C(_09113_),
    .Y(_09231_));
 AO21x1_ASAP7_75t_SL _17404_ (.A1(_08917_),
    .A2(_08912_),
    .B(_01006_),
    .Y(_09232_));
 INVx1_ASAP7_75t_R _17405_ (.A(_09232_),
    .Y(_09233_));
 NOR2x1_ASAP7_75t_R _17406_ (.A(_09233_),
    .B(_09064_),
    .Y(_09234_));
 OAI21x1_ASAP7_75t_R _17407_ (.A1(_09231_),
    .A2(_09234_),
    .B(_08929_),
    .Y(_09235_));
 AO21x1_ASAP7_75t_R _17408_ (.A1(_09006_),
    .A2(_08918_),
    .B(_08924_),
    .Y(_09236_));
 INVx1_ASAP7_75t_R _17409_ (.A(_09236_),
    .Y(_09237_));
 AOI21x1_ASAP7_75t_R _17410_ (.A1(_09212_),
    .A2(_09237_),
    .B(_09033_),
    .Y(_09238_));
 AOI21x1_ASAP7_75t_R _17411_ (.A1(_09020_),
    .A2(_09238_),
    .B(_08933_),
    .Y(_09239_));
 NAND2x1_ASAP7_75t_R _17412_ (.A(_09235_),
    .B(_09239_),
    .Y(_09240_));
 OA21x2_ASAP7_75t_R _17413_ (.A1(_08918_),
    .A2(_09159_),
    .B(_08924_),
    .Y(_09241_));
 NAND2x1_ASAP7_75t_SL _17414_ (.A(_09028_),
    .B(_09241_),
    .Y(_09242_));
 AO21x1_ASAP7_75t_R _17415_ (.A1(_09121_),
    .A2(_09184_),
    .B(_08924_),
    .Y(_09243_));
 AOI21x1_ASAP7_75t_R _17416_ (.A1(_09242_),
    .A2(_09243_),
    .B(_09020_),
    .Y(_09244_));
 AOI21x1_ASAP7_75t_R _17417_ (.A1(_08925_),
    .A2(_09177_),
    .B(_08929_),
    .Y(_09245_));
 AO21x1_ASAP7_75t_SL _17418_ (.A1(_09134_),
    .A2(_09121_),
    .B(_08925_),
    .Y(_09246_));
 AND2x2_ASAP7_75t_L _17419_ (.A(_09245_),
    .B(_09246_),
    .Y(_09247_));
 OAI21x1_ASAP7_75t_SL _17420_ (.A1(_09247_),
    .A2(_09244_),
    .B(_08933_),
    .Y(_09248_));
 AOI21x1_ASAP7_75t_SL _17421_ (.A1(_09248_),
    .A2(_09240_),
    .B(_08938_),
    .Y(_09249_));
 INVx1_ASAP7_75t_SL _17422_ (.A(_09100_),
    .Y(_09250_));
 AO21x1_ASAP7_75t_SL _17423_ (.A1(_09250_),
    .A2(_09107_),
    .B(_08925_),
    .Y(_09251_));
 AO21x1_ASAP7_75t_R _17424_ (.A1(_09055_),
    .A2(_09107_),
    .B(_08924_),
    .Y(_09252_));
 NAND3x1_ASAP7_75t_R _17425_ (.A(_09251_),
    .B(_09252_),
    .C(_09020_),
    .Y(_09253_));
 AO21x1_ASAP7_75t_R _17426_ (.A1(_09027_),
    .A2(_08918_),
    .B(_08925_),
    .Y(_09254_));
 OAI21x1_ASAP7_75t_R _17427_ (.A1(_09108_),
    .A2(_09064_),
    .B(_09254_),
    .Y(_09255_));
 AOI21x1_ASAP7_75t_R _17428_ (.A1(_09102_),
    .A2(_09255_),
    .B(_08934_),
    .Y(_09256_));
 NAND2x1_ASAP7_75t_R _17429_ (.A(_09253_),
    .B(_09256_),
    .Y(_09257_));
 NAND2x1p5_ASAP7_75t_SL _17430_ (.A(_09026_),
    .B(_09056_),
    .Y(_09258_));
 NOR2x1_ASAP7_75t_R _17431_ (.A(_08925_),
    .B(_09078_),
    .Y(_09259_));
 NAND2x1_ASAP7_75t_SL _17432_ (.A(_09030_),
    .B(_09259_),
    .Y(_09260_));
 AOI21x1_ASAP7_75t_SL _17433_ (.A1(_09260_),
    .A2(_09258_),
    .B(_08929_),
    .Y(_09261_));
 AO21x1_ASAP7_75t_R _17434_ (.A1(_09250_),
    .A2(_09113_),
    .B(_08924_),
    .Y(_09262_));
 AND2x2_ASAP7_75t_R _17435_ (.A(_08918_),
    .B(_09027_),
    .Y(_09263_));
 NOR2x1_ASAP7_75t_R _17436_ (.A(_08918_),
    .B(_08907_),
    .Y(_09264_));
 OAI21x1_ASAP7_75t_R _17437_ (.A1(_09263_),
    .A2(_09264_),
    .B(_08924_),
    .Y(_09265_));
 AOI21x1_ASAP7_75t_R _17438_ (.A1(_09262_),
    .A2(_09265_),
    .B(_09020_),
    .Y(_09266_));
 OAI21x1_ASAP7_75t_SL _17439_ (.A1(_09266_),
    .A2(_09261_),
    .B(_08934_),
    .Y(_09267_));
 AOI21x1_ASAP7_75t_SL _17440_ (.A1(_09267_),
    .A2(_09257_),
    .B(_08937_),
    .Y(_09268_));
 OAI21x1_ASAP7_75t_SL _17441_ (.A1(_09268_),
    .A2(_09249_),
    .B(_09025_),
    .Y(_09269_));
 INVx1_ASAP7_75t_R _17442_ (.A(_01010_),
    .Y(_09270_));
 OAI21x1_ASAP7_75t_SL _17444_ (.A1(_09270_),
    .A2(_09264_),
    .B(_08925_),
    .Y(_09272_));
 AOI21x1_ASAP7_75t_R _17445_ (.A1(_09246_),
    .A2(_09272_),
    .B(_09020_),
    .Y(_09273_));
 NAND2x1_ASAP7_75t_SL _17446_ (.A(_09095_),
    .B(_08924_),
    .Y(_09274_));
 AND2x4_ASAP7_75t_SL _17447_ (.A(_08925_),
    .B(_09134_),
    .Y(_09275_));
 NAND2x1_ASAP7_75t_L _17448_ (.A(_09088_),
    .B(_09275_),
    .Y(_09276_));
 AOI21x1_ASAP7_75t_SL _17449_ (.A1(_09274_),
    .A2(_09276_),
    .B(_08929_),
    .Y(_09277_));
 OA21x2_ASAP7_75t_SL _17450_ (.A1(_09277_),
    .A2(_09273_),
    .B(_08934_),
    .Y(_09278_));
 NAND2x1_ASAP7_75t_R _17451_ (.A(_01014_),
    .B(_08924_),
    .Y(_09279_));
 AO21x1_ASAP7_75t_SL _17452_ (.A1(_09187_),
    .A2(_09188_),
    .B(_08924_),
    .Y(_09280_));
 AOI21x1_ASAP7_75t_R _17453_ (.A1(_09279_),
    .A2(_09280_),
    .B(_08929_),
    .Y(_09281_));
 AND2x4_ASAP7_75t_SL _17454_ (.A(_09056_),
    .B(_08925_),
    .Y(_09282_));
 AND3x1_ASAP7_75t_R _17455_ (.A(_09055_),
    .B(_08924_),
    .C(_09001_),
    .Y(_09283_));
 AOI211x1_ASAP7_75t_SL _17456_ (.A1(_08997_),
    .A2(_09282_),
    .B(_09283_),
    .C(_09020_),
    .Y(_09284_));
 NOR2x1_ASAP7_75t_SL _17457_ (.A(_09284_),
    .B(_09281_),
    .Y(_09285_));
 OAI21x1_ASAP7_75t_SL _17458_ (.A1(_09285_),
    .A2(_08934_),
    .B(_08938_),
    .Y(_09286_));
 OA21x2_ASAP7_75t_R _17459_ (.A1(_01010_),
    .A2(_08925_),
    .B(_08929_),
    .Y(_09287_));
 AOI21x1_ASAP7_75t_R _17460_ (.A1(_09287_),
    .A2(_09243_),
    .B(_08934_),
    .Y(_09288_));
 AOI21x1_ASAP7_75t_R _17461_ (.A1(_01012_),
    .A2(_08925_),
    .B(_09033_),
    .Y(_09289_));
 NAND2x1_ASAP7_75t_R _17462_ (.A(_09020_),
    .B(_09289_),
    .Y(_09290_));
 NAND2x1_ASAP7_75t_R _17463_ (.A(_09288_),
    .B(_09290_),
    .Y(_09291_));
 NAND2x1_ASAP7_75t_R _17464_ (.A(_09018_),
    .B(_09237_),
    .Y(_09292_));
 NAND3x1_ASAP7_75t_R _17465_ (.A(_09292_),
    .B(_09206_),
    .C(_08929_),
    .Y(_09293_));
 OA21x2_ASAP7_75t_SL _17466_ (.A1(_09126_),
    .A2(_09108_),
    .B(_08925_),
    .Y(_09294_));
 OA21x2_ASAP7_75t_R _17467_ (.A1(_09294_),
    .A2(_09130_),
    .B(_08934_),
    .Y(_09295_));
 AOI21x1_ASAP7_75t_R _17468_ (.A1(_09293_),
    .A2(_09295_),
    .B(_08938_),
    .Y(_09296_));
 AOI21x1_ASAP7_75t_SL _17469_ (.A1(_09296_),
    .A2(_09291_),
    .B(_09025_),
    .Y(_09297_));
 OAI21x1_ASAP7_75t_SL _17470_ (.A1(_09278_),
    .A2(_09286_),
    .B(_09297_),
    .Y(_09298_));
 NAND2x1_ASAP7_75t_SL _17471_ (.A(_09298_),
    .B(_09269_),
    .Y(_00010_));
 AND2x2_ASAP7_75t_SL _17472_ (.A(_08924_),
    .B(_09010_),
    .Y(_09299_));
 AO21x1_ASAP7_75t_SL _17473_ (.A1(_08934_),
    .A2(_09299_),
    .B(_09071_),
    .Y(_09300_));
 AO21x1_ASAP7_75t_SL _17474_ (.A1(_09121_),
    .A2(_09061_),
    .B(_08925_),
    .Y(_09301_));
 AOI21x1_ASAP7_75t_SL _17475_ (.A1(_09136_),
    .A2(_09301_),
    .B(_08934_),
    .Y(_09302_));
 OAI21x1_ASAP7_75t_SL _17476_ (.A1(_09302_),
    .A2(_09300_),
    .B(_08929_),
    .Y(_09303_));
 AND2x2_ASAP7_75t_SL _17477_ (.A(_09100_),
    .B(_08925_),
    .Y(_09304_));
 NOR2x1_ASAP7_75t_SL _17478_ (.A(_08933_),
    .B(_09304_),
    .Y(_09305_));
 AOI21x1_ASAP7_75t_SL _17479_ (.A1(_09305_),
    .A2(_09260_),
    .B(_08929_),
    .Y(_09306_));
 INVx1_ASAP7_75t_SL _17480_ (.A(_09164_),
    .Y(_09307_));
 AOI21x1_ASAP7_75t_SL _17481_ (.A1(_09154_),
    .A2(_09039_),
    .B(_08934_),
    .Y(_09308_));
 OAI21x1_ASAP7_75t_SL _17482_ (.A1(_09264_),
    .A2(_09307_),
    .B(_09308_),
    .Y(_09309_));
 AOI21x1_ASAP7_75t_SL _17483_ (.A1(_09306_),
    .A2(_09309_),
    .B(_08938_),
    .Y(_09310_));
 AOI21x1_ASAP7_75t_SL _17484_ (.A1(_09310_),
    .A2(_09303_),
    .B(_08941_),
    .Y(_09311_));
 AO21x1_ASAP7_75t_SL _17485_ (.A1(_08917_),
    .A2(_08912_),
    .B(_01004_),
    .Y(_09312_));
 AO21x1_ASAP7_75t_R _17486_ (.A1(_09030_),
    .A2(_09312_),
    .B(_08924_),
    .Y(_09313_));
 AOI21x1_ASAP7_75t_SL _17487_ (.A1(_09206_),
    .A2(_09313_),
    .B(_08929_),
    .Y(_09314_));
 INVx1_ASAP7_75t_R _17488_ (.A(_09263_),
    .Y(_09315_));
 AND3x1_ASAP7_75t_SL _17489_ (.A(_09018_),
    .B(_08924_),
    .C(_09315_),
    .Y(_09316_));
 OAI21x1_ASAP7_75t_SL _17490_ (.A1(_09020_),
    .A2(_09316_),
    .B(_08933_),
    .Y(_09317_));
 NOR2x1_ASAP7_75t_SL _17491_ (.A(_09314_),
    .B(_09317_),
    .Y(_09318_));
 NOR2x1_ASAP7_75t_SL _17492_ (.A(_08919_),
    .B(_08995_),
    .Y(_09319_));
 OAI21x1_ASAP7_75t_SL _17493_ (.A1(_09100_),
    .A2(_09319_),
    .B(_08925_),
    .Y(_09320_));
 NAND2x1_ASAP7_75t_SL _17494_ (.A(_09028_),
    .B(_09011_),
    .Y(_09321_));
 NAND3x1_ASAP7_75t_SL _17495_ (.A(_09320_),
    .B(_09321_),
    .C(_08929_),
    .Y(_09322_));
 NAND2x1_ASAP7_75t_SL _17496_ (.A(_09189_),
    .B(_09093_),
    .Y(_09323_));
 AOI21x1_ASAP7_75t_SL _17497_ (.A1(_09323_),
    .A2(_09322_),
    .B(_08933_),
    .Y(_09324_));
 OAI21x1_ASAP7_75t_SL _17498_ (.A1(_09324_),
    .A2(_09318_),
    .B(_08938_),
    .Y(_09325_));
 NAND2x1_ASAP7_75t_SL _17499_ (.A(_09311_),
    .B(_09325_),
    .Y(_09326_));
 AOI21x1_ASAP7_75t_SL _17500_ (.A1(_09184_),
    .A2(_08997_),
    .B(_08924_),
    .Y(_09327_));
 NOR2x1_ASAP7_75t_SL _17501_ (.A(_08925_),
    .B(_09104_),
    .Y(_09328_));
 AND2x2_ASAP7_75t_SL _17502_ (.A(_09134_),
    .B(_09328_),
    .Y(_09329_));
 OAI21x1_ASAP7_75t_SL _17503_ (.A1(_09327_),
    .A2(_09329_),
    .B(_09020_),
    .Y(_09330_));
 NAND2x1_ASAP7_75t_SL _17504_ (.A(_09330_),
    .B(_08934_),
    .Y(_09331_));
 AND2x2_ASAP7_75t_SL _17505_ (.A(_09061_),
    .B(_09011_),
    .Y(_09332_));
 AOI211x1_ASAP7_75t_SL _17506_ (.A1(_09019_),
    .A2(_08925_),
    .B(_09020_),
    .C(_09332_),
    .Y(_09333_));
 NOR2x1_ASAP7_75t_SL _17507_ (.A(_09331_),
    .B(_09333_),
    .Y(_09334_));
 INVx1_ASAP7_75t_SL _17508_ (.A(_09259_),
    .Y(_09335_));
 OAI21x1_ASAP7_75t_SL _17509_ (.A1(_09126_),
    .A2(_09335_),
    .B(_09165_),
    .Y(_09336_));
 NOR2x1_ASAP7_75t_SL _17510_ (.A(_00994_),
    .B(_08995_),
    .Y(_09337_));
 OAI21x1_ASAP7_75t_SL _17511_ (.A1(_09217_),
    .A2(_09337_),
    .B(_08924_),
    .Y(_09338_));
 AO21x1_ASAP7_75t_SL _17512_ (.A1(_09031_),
    .A2(_08918_),
    .B(_08924_),
    .Y(_09339_));
 NAND3x1_ASAP7_75t_SL _17513_ (.A(_09338_),
    .B(_09020_),
    .C(_09339_),
    .Y(_09340_));
 AOI21x1_ASAP7_75t_SL _17514_ (.A1(_09336_),
    .A2(_09340_),
    .B(_08934_),
    .Y(_09341_));
 OAI21x1_ASAP7_75t_SL _17515_ (.A1(_09341_),
    .A2(_09334_),
    .B(_08938_),
    .Y(_09342_));
 AOI21x1_ASAP7_75t_SL _17516_ (.A1(_09107_),
    .A2(_09175_),
    .B(_08924_),
    .Y(_09343_));
 OA21x2_ASAP7_75t_SL _17517_ (.A1(_09343_),
    .A2(_09231_),
    .B(_09020_),
    .Y(_09344_));
 AND3x1_ASAP7_75t_SL _17518_ (.A(_09221_),
    .B(_08925_),
    .C(_09134_),
    .Y(_09345_));
 AOI211x1_ASAP7_75t_SL _17519_ (.A1(_08997_),
    .A2(_09089_),
    .B(_09345_),
    .C(_09020_),
    .Y(_09346_));
 OAI21x1_ASAP7_75t_SL _17520_ (.A1(_09346_),
    .A2(_09344_),
    .B(_08934_),
    .Y(_09347_));
 AO21x1_ASAP7_75t_SL _17521_ (.A1(_09188_),
    .A2(_09127_),
    .B(_08924_),
    .Y(_09348_));
 NAND3x1_ASAP7_75t_SL _17522_ (.A(_09338_),
    .B(_09020_),
    .C(_09348_),
    .Y(_09349_));
 NOR2x1_ASAP7_75t_SL _17523_ (.A(_09020_),
    .B(_09275_),
    .Y(_09350_));
 AO21x1_ASAP7_75t_SL _17524_ (.A1(_09018_),
    .A2(_01010_),
    .B(_08925_),
    .Y(_09351_));
 AOI21x1_ASAP7_75t_SL _17525_ (.A1(_09350_),
    .A2(_09351_),
    .B(_08934_),
    .Y(_09352_));
 AOI21x1_ASAP7_75t_SL _17526_ (.A1(_09349_),
    .A2(_09352_),
    .B(_08938_),
    .Y(_09353_));
 AOI21x1_ASAP7_75t_SL _17527_ (.A1(_09353_),
    .A2(_09347_),
    .B(_09025_),
    .Y(_09354_));
 NAND2x1_ASAP7_75t_SL _17528_ (.A(_09342_),
    .B(_09354_),
    .Y(_09355_));
 NAND2x1_ASAP7_75t_SL _17529_ (.A(_09326_),
    .B(_09355_),
    .Y(_00011_));
 AO21x1_ASAP7_75t_SL _17530_ (.A1(_09013_),
    .A2(_09113_),
    .B(_08925_),
    .Y(_09356_));
 AO21x1_ASAP7_75t_SL _17532_ (.A1(_09055_),
    .A2(_09001_),
    .B(_08924_),
    .Y(_09358_));
 AO21x1_ASAP7_75t_SL _17533_ (.A1(_09356_),
    .A2(_09358_),
    .B(_09020_),
    .Y(_09359_));
 AO21x1_ASAP7_75t_SL _17534_ (.A1(_09030_),
    .A2(_09113_),
    .B(_08925_),
    .Y(_09360_));
 AO21x1_ASAP7_75t_SL _17535_ (.A1(_09280_),
    .A2(_09360_),
    .B(_08929_),
    .Y(_09361_));
 AOI21x1_ASAP7_75t_SL _17536_ (.A1(_09359_),
    .A2(_09361_),
    .B(_08937_),
    .Y(_09362_));
 AO21x1_ASAP7_75t_SL _17537_ (.A1(_09221_),
    .A2(_09188_),
    .B(_08924_),
    .Y(_09363_));
 AO21x1_ASAP7_75t_SL _17538_ (.A1(_09178_),
    .A2(_09363_),
    .B(_08938_),
    .Y(_09364_));
 OA211x2_ASAP7_75t_SL _17539_ (.A1(_09077_),
    .A2(_09196_),
    .B(_09242_),
    .C(_08929_),
    .Y(_09365_));
 OAI21x1_ASAP7_75t_SL _17540_ (.A1(_09364_),
    .A2(_09365_),
    .B(_08941_),
    .Y(_09366_));
 NOR2x1_ASAP7_75t_SL _17541_ (.A(_09362_),
    .B(_09366_),
    .Y(_09367_));
 AO21x1_ASAP7_75t_SL _17542_ (.A1(_09221_),
    .A2(_09113_),
    .B(_08925_),
    .Y(_09368_));
 AND3x1_ASAP7_75t_SL _17543_ (.A(_09194_),
    .B(_09368_),
    .C(_08929_),
    .Y(_09369_));
 AO21x1_ASAP7_75t_SL _17544_ (.A1(_09030_),
    .A2(_09315_),
    .B(_08925_),
    .Y(_09370_));
 OA21x2_ASAP7_75t_SL _17545_ (.A1(_08919_),
    .A2(_08924_),
    .B(_09020_),
    .Y(_09371_));
 AO21x1_ASAP7_75t_SL _17546_ (.A1(_09370_),
    .A2(_09371_),
    .B(_08937_),
    .Y(_09372_));
 OAI21x1_ASAP7_75t_SL _17547_ (.A1(_09369_),
    .A2(_09372_),
    .B(_09025_),
    .Y(_09373_));
 AO21x1_ASAP7_75t_SL _17548_ (.A1(_09018_),
    .A2(_09017_),
    .B(_08924_),
    .Y(_09374_));
 AND3x1_ASAP7_75t_SL _17549_ (.A(_09374_),
    .B(_09020_),
    .C(_09051_),
    .Y(_09375_));
 AND3x1_ASAP7_75t_SL _17550_ (.A(_09013_),
    .B(_08924_),
    .C(_09113_),
    .Y(_09376_));
 NAND2x1_ASAP7_75t_SL _17551_ (.A(_08929_),
    .B(_09313_),
    .Y(_09377_));
 OAI21x1_ASAP7_75t_SL _17552_ (.A1(_09376_),
    .A2(_09377_),
    .B(_08937_),
    .Y(_09378_));
 NOR2x1_ASAP7_75t_SL _17553_ (.A(_09375_),
    .B(_09378_),
    .Y(_09379_));
 OAI21x1_ASAP7_75t_SL _17554_ (.A1(_09373_),
    .A2(_09379_),
    .B(_08933_),
    .Y(_09380_));
 AND2x2_ASAP7_75t_SL _17555_ (.A(_09241_),
    .B(_09056_),
    .Y(_09381_));
 NAND2x1_ASAP7_75t_R _17556_ (.A(_08929_),
    .B(_09236_),
    .Y(_09382_));
 OA21x2_ASAP7_75t_SL _17557_ (.A1(_09382_),
    .A2(_09213_),
    .B(_08938_),
    .Y(_09383_));
 OAI21x1_ASAP7_75t_SL _17558_ (.A1(_09105_),
    .A2(_09381_),
    .B(_09383_),
    .Y(_09384_));
 AO21x1_ASAP7_75t_R _17559_ (.A1(_09055_),
    .A2(_09312_),
    .B(_08924_),
    .Y(_09385_));
 NAND2x1_ASAP7_75t_SL _17560_ (.A(_09385_),
    .B(_09075_),
    .Y(_09386_));
 AO21x1_ASAP7_75t_SL _17561_ (.A1(_00996_),
    .A2(_08924_),
    .B(_08929_),
    .Y(_09387_));
 OA21x2_ASAP7_75t_SL _17562_ (.A1(_09387_),
    .A2(_09282_),
    .B(_08937_),
    .Y(_09388_));
 AOI21x1_ASAP7_75t_SL _17563_ (.A1(_09386_),
    .A2(_09388_),
    .B(_08941_),
    .Y(_09389_));
 AOI21x1_ASAP7_75t_SL _17564_ (.A1(_09384_),
    .A2(_09389_),
    .B(_08933_),
    .Y(_09390_));
 NOR2x1_ASAP7_75t_SL _17565_ (.A(_09020_),
    .B(_09304_),
    .Y(_09391_));
 OR3x1_ASAP7_75t_SL _17566_ (.A(_08919_),
    .B(_00997_),
    .C(_08924_),
    .Y(_09392_));
 AND3x1_ASAP7_75t_SL _17567_ (.A(_09391_),
    .B(_09251_),
    .C(_09392_),
    .Y(_09393_));
 NOR2x1_ASAP7_75t_SL _17568_ (.A(_08925_),
    .B(_09120_),
    .Y(_09394_));
 NAND2x1_ASAP7_75t_SL _17569_ (.A(_09134_),
    .B(_09394_),
    .Y(_09395_));
 AO21x1_ASAP7_75t_SL _17570_ (.A1(_09079_),
    .A2(_09395_),
    .B(_08938_),
    .Y(_09396_));
 AO21x1_ASAP7_75t_R _17571_ (.A1(_01004_),
    .A2(_08918_),
    .B(_08924_),
    .Y(_09397_));
 AND3x1_ASAP7_75t_SL _17572_ (.A(_09397_),
    .B(_08929_),
    .C(_09049_),
    .Y(_09398_));
 NOR2x1_ASAP7_75t_SL _17573_ (.A(_08937_),
    .B(_09398_),
    .Y(_09399_));
 OA21x2_ASAP7_75t_SL _17574_ (.A1(_01015_),
    .A2(_08924_),
    .B(_09020_),
    .Y(_09400_));
 NOR2x1_ASAP7_75t_SL _17575_ (.A(_08924_),
    .B(_08907_),
    .Y(_09401_));
 NAND2x1_ASAP7_75t_SL _17576_ (.A(_08919_),
    .B(_09401_),
    .Y(_09402_));
 NAND3x1_ASAP7_75t_SL _17577_ (.A(_09400_),
    .B(_09202_),
    .C(_09402_),
    .Y(_09403_));
 AOI21x1_ASAP7_75t_SL _17578_ (.A1(_09399_),
    .A2(_09403_),
    .B(_09025_),
    .Y(_09404_));
 OAI21x1_ASAP7_75t_SL _17579_ (.A1(_09393_),
    .A2(_09396_),
    .B(_09404_),
    .Y(_09405_));
 NAND2x1_ASAP7_75t_SL _17580_ (.A(_09390_),
    .B(_09405_),
    .Y(_09406_));
 OAI21x1_ASAP7_75t_SL _17581_ (.A1(_09367_),
    .A2(_09380_),
    .B(_09406_),
    .Y(_00012_));
 NOR2x1_ASAP7_75t_SL _17582_ (.A(_08924_),
    .B(_09056_),
    .Y(_09407_));
 AO21x1_ASAP7_75t_SL _17583_ (.A1(_09213_),
    .A2(_09055_),
    .B(_09407_),
    .Y(_09408_));
 AOI21x1_ASAP7_75t_SL _17584_ (.A1(_08929_),
    .A2(_09408_),
    .B(_08934_),
    .Y(_09409_));
 AO221x1_ASAP7_75t_SL _17585_ (.A1(_08924_),
    .A2(_09315_),
    .B1(_09026_),
    .B2(_09001_),
    .C(_08929_),
    .Y(_09410_));
 NAND2x1_ASAP7_75t_SL _17586_ (.A(_09409_),
    .B(_09410_),
    .Y(_09411_));
 AND3x1_ASAP7_75t_SL _17587_ (.A(_09117_),
    .B(_08925_),
    .C(_09061_),
    .Y(_09412_));
 NAND2x1_ASAP7_75t_SL _17588_ (.A(_00994_),
    .B(_08995_),
    .Y(_09413_));
 AO21x1_ASAP7_75t_SL _17589_ (.A1(_09039_),
    .A2(_09413_),
    .B(_09020_),
    .Y(_09414_));
 NAND2x1_ASAP7_75t_SL _17590_ (.A(_08924_),
    .B(_08995_),
    .Y(_09415_));
 AO21x1_ASAP7_75t_SL _17591_ (.A1(_09415_),
    .A2(_00994_),
    .B(_09114_),
    .Y(_09416_));
 AOI21x1_ASAP7_75t_SL _17592_ (.A1(_09020_),
    .A2(_09416_),
    .B(_08933_),
    .Y(_09417_));
 OAI21x1_ASAP7_75t_SL _17593_ (.A1(_09412_),
    .A2(_09414_),
    .B(_09417_),
    .Y(_09418_));
 AOI21x1_ASAP7_75t_SL _17594_ (.A1(_09411_),
    .A2(_09418_),
    .B(_09025_),
    .Y(_09419_));
 AO21x1_ASAP7_75t_SL _17595_ (.A1(_09315_),
    .A2(_09154_),
    .B(_08925_),
    .Y(_09420_));
 NOR2x1_ASAP7_75t_SL _17596_ (.A(_09126_),
    .B(_09062_),
    .Y(_09421_));
 OA21x2_ASAP7_75t_SL _17597_ (.A1(_09421_),
    .A2(_08924_),
    .B(_08929_),
    .Y(_09422_));
 AO21x1_ASAP7_75t_SL _17598_ (.A1(_01003_),
    .A2(_08925_),
    .B(_08929_),
    .Y(_09423_));
 OAI21x1_ASAP7_75t_SL _17599_ (.A1(_09328_),
    .A2(_09423_),
    .B(_08933_),
    .Y(_09424_));
 AOI21x1_ASAP7_75t_SL _17600_ (.A1(_09420_),
    .A2(_09422_),
    .B(_09424_),
    .Y(_09425_));
 AO21x1_ASAP7_75t_SL _17601_ (.A1(_09170_),
    .A2(_09307_),
    .B(_08933_),
    .Y(_09426_));
 AO21x1_ASAP7_75t_SL _17602_ (.A1(_09117_),
    .A2(_09184_),
    .B(_08925_),
    .Y(_09427_));
 AND3x1_ASAP7_75t_SL _17603_ (.A(_09427_),
    .B(_09020_),
    .C(_09064_),
    .Y(_09428_));
 OAI21x1_ASAP7_75t_SL _17604_ (.A1(_09426_),
    .A2(_09428_),
    .B(_09025_),
    .Y(_09429_));
 OAI21x1_ASAP7_75t_SL _17605_ (.A1(_09425_),
    .A2(_09429_),
    .B(_08937_),
    .Y(_09430_));
 OAI21x1_ASAP7_75t_SL _17606_ (.A1(_09401_),
    .A2(_09015_),
    .B(_09020_),
    .Y(_09431_));
 AO21x1_ASAP7_75t_SL _17607_ (.A1(_09184_),
    .A2(_09127_),
    .B(_08924_),
    .Y(_09432_));
 AO21x1_ASAP7_75t_SL _17608_ (.A1(_09055_),
    .A2(_09312_),
    .B(_08925_),
    .Y(_09433_));
 AO21x1_ASAP7_75t_SL _17609_ (.A1(_09432_),
    .A2(_09433_),
    .B(_09020_),
    .Y(_09434_));
 AOI21x1_ASAP7_75t_SL _17610_ (.A1(_09431_),
    .A2(_09434_),
    .B(_08933_),
    .Y(_09435_));
 OA21x2_ASAP7_75t_SL _17611_ (.A1(_08924_),
    .A2(_09061_),
    .B(_08929_),
    .Y(_09436_));
 NAND2x1_ASAP7_75t_SL _17612_ (.A(_09028_),
    .B(_09328_),
    .Y(_09437_));
 AO21x1_ASAP7_75t_SL _17613_ (.A1(_09436_),
    .A2(_09437_),
    .B(_08934_),
    .Y(_09438_));
 OA21x2_ASAP7_75t_SL _17614_ (.A1(_09264_),
    .A2(_09108_),
    .B(_08924_),
    .Y(_09439_));
 NOR2x1_ASAP7_75t_SL _17615_ (.A(_09105_),
    .B(_09439_),
    .Y(_09440_));
 OAI21x1_ASAP7_75t_SL _17616_ (.A1(_09438_),
    .A2(_09440_),
    .B(_09025_),
    .Y(_09441_));
 OAI21x1_ASAP7_75t_SL _17617_ (.A1(_09435_),
    .A2(_09441_),
    .B(_08938_),
    .Y(_09442_));
 NAND2x1_ASAP7_75t_SL _17618_ (.A(_09181_),
    .B(_09164_),
    .Y(_09443_));
 AO21x1_ASAP7_75t_SL _17619_ (.A1(_09115_),
    .A2(_09443_),
    .B(_08933_),
    .Y(_09444_));
 OA21x2_ASAP7_75t_SL _17620_ (.A1(_08919_),
    .A2(_09159_),
    .B(_08925_),
    .Y(_09445_));
 AOI221x1_ASAP7_75t_SL _17621_ (.A1(_09088_),
    .A2(_09259_),
    .B1(_09018_),
    .B2(_09445_),
    .C(_09020_),
    .Y(_09446_));
 NAND2x1_ASAP7_75t_SL _17622_ (.A(_09184_),
    .B(_08929_),
    .Y(_09447_));
 OA21x2_ASAP7_75t_SL _17623_ (.A1(_09447_),
    .A2(_09241_),
    .B(_08933_),
    .Y(_09448_));
 NOR2x1p5_ASAP7_75t_SL _17624_ (.A(_09011_),
    .B(_08929_),
    .Y(_09449_));
 NAND2x1p5_ASAP7_75t_SL _17625_ (.A(_09449_),
    .B(_09320_),
    .Y(_09450_));
 AOI21x1_ASAP7_75t_SL _17626_ (.A1(_09448_),
    .A2(_09450_),
    .B(_09025_),
    .Y(_09451_));
 OA21x2_ASAP7_75t_SL _17627_ (.A1(_09444_),
    .A2(_09446_),
    .B(_09451_),
    .Y(_09452_));
 OAI22x1_ASAP7_75t_SL _17628_ (.A1(_09419_),
    .A2(_09430_),
    .B1(_09442_),
    .B2(_09452_),
    .Y(_00013_));
 NAND2x1_ASAP7_75t_R _17629_ (.A(_09127_),
    .B(_09213_),
    .Y(_09453_));
 AO21x1_ASAP7_75t_R _17630_ (.A1(_09055_),
    .A2(_09184_),
    .B(_08924_),
    .Y(_09454_));
 AOI21x1_ASAP7_75t_R _17631_ (.A1(_09453_),
    .A2(_09454_),
    .B(_08929_),
    .Y(_09455_));
 AO21x1_ASAP7_75t_SL _17632_ (.A1(_09010_),
    .A2(_08924_),
    .B(_09020_),
    .Y(_09456_));
 NOR2x1_ASAP7_75t_L _17633_ (.A(_09456_),
    .B(_09289_),
    .Y(_09457_));
 OAI21x1_ASAP7_75t_SL _17634_ (.A1(_09457_),
    .A2(_09455_),
    .B(_08934_),
    .Y(_09458_));
 OAI21x1_ASAP7_75t_SL _17635_ (.A1(_09150_),
    .A2(_09135_),
    .B(_08924_),
    .Y(_09459_));
 OAI21x1_ASAP7_75t_SL _17636_ (.A1(_09217_),
    .A2(_09077_),
    .B(_09459_),
    .Y(_09460_));
 NOR2x1_ASAP7_75t_R _17637_ (.A(_09020_),
    .B(_09069_),
    .Y(_09461_));
 AO21x1_ASAP7_75t_R _17638_ (.A1(_09074_),
    .A2(_09113_),
    .B(_08924_),
    .Y(_09462_));
 AOI21x1_ASAP7_75t_R _17639_ (.A1(_09461_),
    .A2(_09462_),
    .B(_08934_),
    .Y(_09463_));
 OAI21x1_ASAP7_75t_SL _17640_ (.A1(_09460_),
    .A2(_08929_),
    .B(_09463_),
    .Y(_09464_));
 AOI21x1_ASAP7_75t_SL _17641_ (.A1(_09464_),
    .A2(_09458_),
    .B(_08938_),
    .Y(_09465_));
 NAND2x1_ASAP7_75t_R _17642_ (.A(_08924_),
    .B(_09129_),
    .Y(_09466_));
 OA21x2_ASAP7_75t_R _17643_ (.A1(_08924_),
    .A2(_09232_),
    .B(_09466_),
    .Y(_09467_));
 AOI21x1_ASAP7_75t_R _17644_ (.A1(_09391_),
    .A2(_09467_),
    .B(_08933_),
    .Y(_09468_));
 OA21x2_ASAP7_75t_R _17645_ (.A1(_00994_),
    .A2(_08925_),
    .B(_09020_),
    .Y(_09469_));
 AO21x1_ASAP7_75t_SL _17646_ (.A1(_09413_),
    .A2(_09121_),
    .B(_08924_),
    .Y(_09470_));
 NAND2x1_ASAP7_75t_R _17647_ (.A(_09469_),
    .B(_09470_),
    .Y(_09471_));
 NAND2x1_ASAP7_75t_R _17648_ (.A(_09468_),
    .B(_09471_),
    .Y(_09472_));
 AO21x1_ASAP7_75t_R _17649_ (.A1(_09175_),
    .A2(_09312_),
    .B(_08925_),
    .Y(_09473_));
 AO21x1_ASAP7_75t_R _17650_ (.A1(_09049_),
    .A2(_09155_),
    .B(_08924_),
    .Y(_09474_));
 AOI21x1_ASAP7_75t_R _17651_ (.A1(_09473_),
    .A2(_09474_),
    .B(_08929_),
    .Y(_09475_));
 AOI21x1_ASAP7_75t_SL _17652_ (.A1(_09320_),
    .A2(_09459_),
    .B(_09020_),
    .Y(_09476_));
 OAI21x1_ASAP7_75t_SL _17653_ (.A1(_09476_),
    .A2(_09475_),
    .B(_08933_),
    .Y(_09477_));
 AOI21x1_ASAP7_75t_SL _17654_ (.A1(_09477_),
    .A2(_09472_),
    .B(_08937_),
    .Y(_09478_));
 OAI21x1_ASAP7_75t_SL _17655_ (.A1(_09478_),
    .A2(_09465_),
    .B(_08941_),
    .Y(_09479_));
 AO21x1_ASAP7_75t_R _17656_ (.A1(_09217_),
    .A2(_08924_),
    .B(_09020_),
    .Y(_09480_));
 AND3x1_ASAP7_75t_L _17657_ (.A(_09028_),
    .B(_08925_),
    .C(_09127_),
    .Y(_09481_));
 AOI21x1_ASAP7_75t_R _17658_ (.A1(_01009_),
    .A2(_08925_),
    .B(_08929_),
    .Y(_09482_));
 AOI21x1_ASAP7_75t_R _17659_ (.A1(_09482_),
    .A2(_09433_),
    .B(_08933_),
    .Y(_09483_));
 OAI21x1_ASAP7_75t_R _17660_ (.A1(_09480_),
    .A2(_09481_),
    .B(_09483_),
    .Y(_09484_));
 AO21x1_ASAP7_75t_R _17661_ (.A1(_09060_),
    .A2(_08918_),
    .B(_08925_),
    .Y(_09485_));
 AOI21x1_ASAP7_75t_R _17662_ (.A1(_09485_),
    .A2(_09385_),
    .B(_09020_),
    .Y(_09486_));
 OAI21x1_ASAP7_75t_R _17663_ (.A1(_09245_),
    .A2(_09486_),
    .B(_08933_),
    .Y(_09487_));
 AOI21x1_ASAP7_75t_R _17664_ (.A1(_09484_),
    .A2(_09487_),
    .B(_08938_),
    .Y(_09488_));
 AOI21x1_ASAP7_75t_R _17665_ (.A1(_09171_),
    .A2(_09034_),
    .B(_09020_),
    .Y(_09489_));
 NAND2x1_ASAP7_75t_SL _17666_ (.A(_08924_),
    .B(_09126_),
    .Y(_09490_));
 AOI21x1_ASAP7_75t_R _17667_ (.A1(_09490_),
    .A2(_09320_),
    .B(_08929_),
    .Y(_09491_));
 OAI21x1_ASAP7_75t_R _17668_ (.A1(_09489_),
    .A2(_09491_),
    .B(_08933_),
    .Y(_09492_));
 NAND2x1_ASAP7_75t_R _17669_ (.A(_09394_),
    .B(_09014_),
    .Y(_09493_));
 NOR2x1_ASAP7_75t_R _17670_ (.A(_01002_),
    .B(_08995_),
    .Y(_09494_));
 OAI21x1_ASAP7_75t_R _17671_ (.A1(_09264_),
    .A2(_09494_),
    .B(_08925_),
    .Y(_09495_));
 AOI21x1_ASAP7_75t_R _17672_ (.A1(_09493_),
    .A2(_09495_),
    .B(_09020_),
    .Y(_09496_));
 AO21x1_ASAP7_75t_R _17673_ (.A1(_09121_),
    .A2(_09184_),
    .B(_08925_),
    .Y(_09497_));
 OAI21x1_ASAP7_75t_R _17674_ (.A1(_09217_),
    .A2(_09337_),
    .B(_08925_),
    .Y(_09498_));
 AOI21x1_ASAP7_75t_R _17675_ (.A1(_09497_),
    .A2(_09498_),
    .B(_08929_),
    .Y(_09499_));
 OAI21x1_ASAP7_75t_R _17676_ (.A1(_09496_),
    .A2(_09499_),
    .B(_08934_),
    .Y(_09500_));
 AOI21x1_ASAP7_75t_R _17677_ (.A1(_09492_),
    .A2(_09500_),
    .B(_08937_),
    .Y(_09501_));
 OAI21x1_ASAP7_75t_R _17678_ (.A1(_09488_),
    .A2(_09501_),
    .B(_09025_),
    .Y(_09502_));
 NAND2x1_ASAP7_75t_SL _17679_ (.A(_09479_),
    .B(_09502_),
    .Y(_00014_));
 NOR2x1_ASAP7_75t_SL _17680_ (.A(_09092_),
    .B(_08929_),
    .Y(_09503_));
 AO21x1_ASAP7_75t_SL _17681_ (.A1(_08925_),
    .A2(_09188_),
    .B(_09213_),
    .Y(_09504_));
 AOI21x1_ASAP7_75t_SL _17682_ (.A1(_09503_),
    .A2(_09504_),
    .B(_08934_),
    .Y(_09505_));
 NAND2x1_ASAP7_75t_SL _17683_ (.A(_09159_),
    .B(_08924_),
    .Y(_09506_));
 AO21x1_ASAP7_75t_SL _17684_ (.A1(_09470_),
    .A2(_09506_),
    .B(_09020_),
    .Y(_09507_));
 NAND2x1_ASAP7_75t_SL _17685_ (.A(_09505_),
    .B(_09507_),
    .Y(_09508_));
 AO21x1_ASAP7_75t_SL _17686_ (.A1(_09154_),
    .A2(_09061_),
    .B(_08924_),
    .Y(_09509_));
 AO21x1_ASAP7_75t_SL _17687_ (.A1(_09221_),
    .A2(_09155_),
    .B(_08925_),
    .Y(_09510_));
 AND3x1_ASAP7_75t_SL _17688_ (.A(_09509_),
    .B(_09510_),
    .C(_09020_),
    .Y(_09511_));
 AND3x1_ASAP7_75t_SL _17689_ (.A(_09008_),
    .B(_08924_),
    .C(_09055_),
    .Y(_09512_));
 NOR2x1_ASAP7_75t_SL _17690_ (.A(_09512_),
    .B(_09377_),
    .Y(_09513_));
 OAI21x1_ASAP7_75t_SL _17691_ (.A1(_09511_),
    .A2(_09513_),
    .B(_08934_),
    .Y(_09514_));
 AOI21x1_ASAP7_75t_SL _17692_ (.A1(_09514_),
    .A2(_09508_),
    .B(_08937_),
    .Y(_09515_));
 NOR2x1_ASAP7_75t_SL _17693_ (.A(_00996_),
    .B(_08924_),
    .Y(_09516_));
 AO21x1_ASAP7_75t_SL _17694_ (.A1(_08924_),
    .A2(_09232_),
    .B(_09516_),
    .Y(_09517_));
 AO21x1_ASAP7_75t_SL _17695_ (.A1(_09517_),
    .A2(_09020_),
    .B(_08933_),
    .Y(_09518_));
 INVx1_ASAP7_75t_SL _17696_ (.A(_09114_),
    .Y(_09519_));
 AND3x1_ASAP7_75t_SL _17697_ (.A(_09075_),
    .B(_09519_),
    .C(_09194_),
    .Y(_09520_));
 NOR2x1_ASAP7_75t_SL _17698_ (.A(_09518_),
    .B(_09520_),
    .Y(_09521_));
 NOR2x1_ASAP7_75t_SL _17699_ (.A(_08925_),
    .B(_09134_),
    .Y(_09522_));
 NAND2x1_ASAP7_75t_SL _17700_ (.A(_09101_),
    .B(_09400_),
    .Y(_09523_));
 OAI21x1_ASAP7_75t_SL _17701_ (.A1(_09522_),
    .A2(_09523_),
    .B(_08933_),
    .Y(_09524_));
 NAND2x1_ASAP7_75t_SL _17702_ (.A(_08924_),
    .B(_09217_),
    .Y(_09525_));
 AO21x1_ASAP7_75t_SL _17703_ (.A1(_09154_),
    .A2(_09056_),
    .B(_08924_),
    .Y(_09526_));
 AND4x1_ASAP7_75t_SL _17704_ (.A(_09525_),
    .B(_09526_),
    .C(_08929_),
    .D(_09274_),
    .Y(_09527_));
 OAI21x1_ASAP7_75t_SL _17705_ (.A1(_09527_),
    .A2(_09524_),
    .B(_08937_),
    .Y(_09528_));
 OAI21x1_ASAP7_75t_SL _17706_ (.A1(_09528_),
    .A2(_09521_),
    .B(_08941_),
    .Y(_09529_));
 OA21x2_ASAP7_75t_SL _17707_ (.A1(_08925_),
    .A2(_09007_),
    .B(_09077_),
    .Y(_09530_));
 NAND2x1_ASAP7_75t_SL _17708_ (.A(_08929_),
    .B(_09490_),
    .Y(_09531_));
 OAI21x1_ASAP7_75t_SL _17709_ (.A1(_08924_),
    .A2(_09116_),
    .B(_09449_),
    .Y(_09532_));
 OAI21x1_ASAP7_75t_SL _17710_ (.A1(_09530_),
    .A2(_09531_),
    .B(_09532_),
    .Y(_09533_));
 AOI21x1_ASAP7_75t_SL _17711_ (.A1(_08933_),
    .A2(_09533_),
    .B(_08938_),
    .Y(_09534_));
 AO21x1_ASAP7_75t_SL _17712_ (.A1(_09055_),
    .A2(_09155_),
    .B(_08925_),
    .Y(_09535_));
 NAND2x1_ASAP7_75t_SL _17713_ (.A(_09535_),
    .B(_09280_),
    .Y(_09536_));
 NOR2x1_ASAP7_75t_SL _17714_ (.A(_09196_),
    .B(_09064_),
    .Y(_09537_));
 NAND2x1_ASAP7_75t_SL _17715_ (.A(_08929_),
    .B(_09415_),
    .Y(_09538_));
 OA21x2_ASAP7_75t_SL _17716_ (.A1(_09537_),
    .A2(_09538_),
    .B(_08934_),
    .Y(_09539_));
 OAI21x1_ASAP7_75t_SL _17717_ (.A1(_08929_),
    .A2(_09536_),
    .B(_09539_),
    .Y(_09540_));
 NAND2x1_ASAP7_75t_SL _17718_ (.A(_09540_),
    .B(_09534_),
    .Y(_09541_));
 NOR2x1_ASAP7_75t_SL _17719_ (.A(_08929_),
    .B(_09394_),
    .Y(_09542_));
 AOI21x1_ASAP7_75t_SL _17720_ (.A1(_09542_),
    .A2(_09385_),
    .B(_08933_),
    .Y(_09543_));
 OAI21x1_ASAP7_75t_SL _17721_ (.A1(_09092_),
    .A2(_09236_),
    .B(_08929_),
    .Y(_09544_));
 AO21x1_ASAP7_75t_SL _17722_ (.A1(_09039_),
    .A2(_09088_),
    .B(_09544_),
    .Y(_09545_));
 AOI21x1_ASAP7_75t_SL _17723_ (.A1(_09543_),
    .A2(_09545_),
    .B(_08937_),
    .Y(_09546_));
 AO22x2_ASAP7_75t_SL _17724_ (.A1(_09039_),
    .A2(_09154_),
    .B1(_09212_),
    .B2(_09275_),
    .Y(_09547_));
 AOI21x1_ASAP7_75t_SL _17725_ (.A1(_09212_),
    .A2(_09259_),
    .B(_08929_),
    .Y(_09548_));
 AOI21x1_ASAP7_75t_SL _17726_ (.A1(_09272_),
    .A2(_09548_),
    .B(_08934_),
    .Y(_09549_));
 OAI21x1_ASAP7_75t_SL _17727_ (.A1(_09547_),
    .A2(_09020_),
    .B(_09549_),
    .Y(_09550_));
 AOI21x1_ASAP7_75t_SL _17728_ (.A1(_09550_),
    .A2(_09546_),
    .B(_08941_),
    .Y(_09551_));
 NAND2x1_ASAP7_75t_SL _17729_ (.A(_09551_),
    .B(_09541_),
    .Y(_09552_));
 OAI21x1_ASAP7_75t_SL _17730_ (.A1(_09515_),
    .A2(_09529_),
    .B(_09552_),
    .Y(_00015_));
 XOR2x2_ASAP7_75t_SL _17731_ (.A(_00945_),
    .B(_08787_),
    .Y(_09553_));
 AOI21x1_ASAP7_75t_SL _17732_ (.A1(_08005_),
    .A2(_09553_),
    .B(_08869_),
    .Y(_09554_));
 XOR2x2_ASAP7_75t_SL _17736_ (.A(_00934_),
    .B(_08785_),
    .Y(_09556_));
 AOI21x1_ASAP7_75t_SL _17737_ (.A1(_09556_),
    .A2(_08005_),
    .B(_08864_),
    .Y(_09557_));
 INVx1_ASAP7_75t_SL _17739_ (.A(_01019_),
    .Y(_09558_));
 NOR2x1p5_ASAP7_75t_SL _17740_ (.A(_09558_),
    .B(_08878_),
    .Y(_09559_));
 INVx2_ASAP7_75t_SL _17741_ (.A(_09559_),
    .Y(_09560_));
 AO21x2_ASAP7_75t_R _17743_ (.A1(_08877_),
    .A2(_08872_),
    .B(_01018_),
    .Y(_09562_));
 AND3x1_ASAP7_75t_SL _17744_ (.A(_09560_),
    .B(_08884_),
    .C(_09562_),
    .Y(_09563_));
 INVx1_ASAP7_75t_SL _17745_ (.A(_01025_),
    .Y(_09564_));
 NAND2x1_ASAP7_75t_R _17747_ (.A(_09564_),
    .B(_08879_),
    .Y(_09566_));
 AO21x1_ASAP7_75t_R _17751_ (.A1(_08877_),
    .A2(_08872_),
    .B(_01027_),
    .Y(_09570_));
 AND3x1_ASAP7_75t_R _17752_ (.A(_09566_),
    .B(_08885_),
    .C(_09570_),
    .Y(_09571_));
 INVx2_ASAP7_75t_SL _17753_ (.A(_08890_),
    .Y(_09572_));
 OA21x2_ASAP7_75t_R _17755_ (.A1(_09563_),
    .A2(_09571_),
    .B(_09572_),
    .Y(_09574_));
 NAND2x1_ASAP7_75t_SL _17756_ (.A(_08866_),
    .B(_08871_),
    .Y(_09575_));
 AOI21x1_ASAP7_75t_R _17757_ (.A1(_08879_),
    .A2(_09557_),
    .B(_08885_),
    .Y(_09576_));
 NAND2x1_ASAP7_75t_SL _17758_ (.A(_09575_),
    .B(_09576_),
    .Y(_09577_));
 NAND2x1_ASAP7_75t_SL _17759_ (.A(_08879_),
    .B(_09557_),
    .Y(_09578_));
 AO21x1_ASAP7_75t_R _17762_ (.A1(_09575_),
    .A2(_09578_),
    .B(_08884_),
    .Y(_09581_));
 AOI21x1_ASAP7_75t_R _17763_ (.A1(_09577_),
    .A2(_09581_),
    .B(_09572_),
    .Y(_09582_));
 OAI21x1_ASAP7_75t_R _17764_ (.A1(_09574_),
    .A2(_09582_),
    .B(_08894_),
    .Y(_09583_));
 INVx1_ASAP7_75t_SL _17765_ (.A(_08894_),
    .Y(_09584_));
 NOR2x1_ASAP7_75t_SL _17769_ (.A(_08878_),
    .B(_01019_),
    .Y(_09588_));
 AO21x1_ASAP7_75t_R _17770_ (.A1(_09554_),
    .A2(_08878_),
    .B(_09588_),
    .Y(_09589_));
 AO21x2_ASAP7_75t_SL _17771_ (.A1(_08877_),
    .A2(_08872_),
    .B(_09558_),
    .Y(_09590_));
 NAND2x1p5_ASAP7_75t_SL _17772_ (.A(_09590_),
    .B(_08885_),
    .Y(_09591_));
 AND2x4_ASAP7_75t_SL _17773_ (.A(_09591_),
    .B(_08890_),
    .Y(_09592_));
 OAI21x1_ASAP7_75t_SL _17774_ (.A1(_08885_),
    .A2(_09589_),
    .B(_09592_),
    .Y(_09593_));
 AO21x1_ASAP7_75t_R _17775_ (.A1(_08877_),
    .A2(_08872_),
    .B(_09564_),
    .Y(_09594_));
 NAND2x1_ASAP7_75t_SL _17777_ (.A(_01027_),
    .B(_08879_),
    .Y(_09596_));
 AOI21x1_ASAP7_75t_R _17778_ (.A1(_09594_),
    .A2(_09596_),
    .B(_08885_),
    .Y(_09597_));
 NOR2x2_ASAP7_75t_SL _17779_ (.A(_09559_),
    .B(_08884_),
    .Y(_09598_));
 AND2x2_ASAP7_75t_SL _17780_ (.A(_09570_),
    .B(_09598_),
    .Y(_09599_));
 OAI21x1_ASAP7_75t_SL _17781_ (.A1(_09599_),
    .A2(_09597_),
    .B(_09572_),
    .Y(_09600_));
 NAND2x1_ASAP7_75t_SL _17782_ (.A(_09600_),
    .B(_09593_),
    .Y(_09601_));
 AOI21x1_ASAP7_75t_SL _17783_ (.A1(_09584_),
    .A2(_09601_),
    .B(_08902_),
    .Y(_09602_));
 NAND2x1_ASAP7_75t_SL _17784_ (.A(_09602_),
    .B(_09583_),
    .Y(_09603_));
 NOR2x1_ASAP7_75t_SL _17785_ (.A(_08879_),
    .B(_09557_),
    .Y(_09604_));
 INVx1_ASAP7_75t_SL _17786_ (.A(_01022_),
    .Y(_09605_));
 NOR2x1_ASAP7_75t_L _17787_ (.A(_09605_),
    .B(_08878_),
    .Y(_09606_));
 OA21x2_ASAP7_75t_R _17789_ (.A1(_09604_),
    .A2(_09606_),
    .B(_08884_),
    .Y(_09608_));
 NOR2x1_ASAP7_75t_L _17790_ (.A(_01027_),
    .B(_08878_),
    .Y(_09609_));
 INVx1_ASAP7_75t_R _17791_ (.A(_09609_),
    .Y(_09610_));
 AOI21x1_ASAP7_75t_R _17792_ (.A1(_08878_),
    .A2(_08866_),
    .B(_08884_),
    .Y(_09611_));
 AOI21x1_ASAP7_75t_R _17794_ (.A1(_09610_),
    .A2(_09611_),
    .B(_08890_),
    .Y(_09613_));
 INVx1_ASAP7_75t_R _17795_ (.A(_09613_),
    .Y(_09614_));
 AO21x2_ASAP7_75t_SL _17798_ (.A1(_08877_),
    .A2(_08872_),
    .B(_01019_),
    .Y(_09617_));
 AND2x4_ASAP7_75t_L _17799_ (.A(_09617_),
    .B(_08884_),
    .Y(_09618_));
 AO21x1_ASAP7_75t_R _17800_ (.A1(_01035_),
    .A2(_08885_),
    .B(_09618_),
    .Y(_09619_));
 AOI21x1_ASAP7_75t_R _17802_ (.A1(_08890_),
    .A2(_09619_),
    .B(_08894_),
    .Y(_09621_));
 OAI21x1_ASAP7_75t_SL _17803_ (.A1(_09608_),
    .A2(_09614_),
    .B(_09621_),
    .Y(_09622_));
 INVx1_ASAP7_75t_R _17804_ (.A(_09606_),
    .Y(_09623_));
 AO21x1_ASAP7_75t_R _17805_ (.A1(_09623_),
    .A2(_09594_),
    .B(_08885_),
    .Y(_09624_));
 NOR2x1_ASAP7_75t_R _17806_ (.A(_01028_),
    .B(_08878_),
    .Y(_09625_));
 INVx1_ASAP7_75t_R _17807_ (.A(_09625_),
    .Y(_09626_));
 OA21x2_ASAP7_75t_R _17809_ (.A1(_09626_),
    .A2(_08884_),
    .B(_08890_),
    .Y(_09628_));
 AOI21x1_ASAP7_75t_R _17810_ (.A1(_09624_),
    .A2(_09628_),
    .B(_09584_),
    .Y(_09629_));
 NAND2x1_ASAP7_75t_R _17811_ (.A(_08884_),
    .B(_09625_),
    .Y(_09630_));
 AO21x1_ASAP7_75t_R _17812_ (.A1(_08877_),
    .A2(_08872_),
    .B(_01026_),
    .Y(_09631_));
 AO21x1_ASAP7_75t_R _17813_ (.A1(_09623_),
    .A2(_09631_),
    .B(_08884_),
    .Y(_09632_));
 AND2x2_ASAP7_75t_R _17814_ (.A(_09632_),
    .B(_09572_),
    .Y(_09633_));
 NAND2x1_ASAP7_75t_R _17815_ (.A(_09630_),
    .B(_09633_),
    .Y(_09634_));
 INVx2_ASAP7_75t_SL _17816_ (.A(_08902_),
    .Y(_09635_));
 AOI21x1_ASAP7_75t_R _17817_ (.A1(_09629_),
    .A2(_09634_),
    .B(_09635_),
    .Y(_09636_));
 AOI21x1_ASAP7_75t_R _17818_ (.A1(_09622_),
    .A2(_09636_),
    .B(_08899_),
    .Y(_09637_));
 NAND2x1_ASAP7_75t_SL _17819_ (.A(_09603_),
    .B(_09637_),
    .Y(_09638_));
 NAND2x1_ASAP7_75t_SL _17820_ (.A(_08879_),
    .B(_08871_),
    .Y(_09639_));
 AND2x2_ASAP7_75t_L _17822_ (.A(_08878_),
    .B(_09605_),
    .Y(_09641_));
 NOR2x1p5_ASAP7_75t_SL _17823_ (.A(_08885_),
    .B(_09641_),
    .Y(_09642_));
 NAND2x1_ASAP7_75t_SL _17824_ (.A(_01020_),
    .B(_08879_),
    .Y(_09643_));
 AND2x2_ASAP7_75t_R _17825_ (.A(_09611_),
    .B(_09643_),
    .Y(_09644_));
 AOI21x1_ASAP7_75t_R _17826_ (.A1(_09639_),
    .A2(_09642_),
    .B(_09644_),
    .Y(_09645_));
 INVx1_ASAP7_75t_SL _17827_ (.A(_01018_),
    .Y(_09646_));
 NAND2x1_ASAP7_75t_SL _17828_ (.A(_09646_),
    .B(_08879_),
    .Y(_09647_));
 AOI21x1_ASAP7_75t_SL _17829_ (.A1(_09647_),
    .A2(_09611_),
    .B(_08890_),
    .Y(_09648_));
 NOR2x1_ASAP7_75t_R _17830_ (.A(_08879_),
    .B(_09554_),
    .Y(_09649_));
 OAI21x1_ASAP7_75t_R _17831_ (.A1(_09625_),
    .A2(_09649_),
    .B(_08884_),
    .Y(_09650_));
 AO21x1_ASAP7_75t_R _17833_ (.A1(_09648_),
    .A2(_09650_),
    .B(_08894_),
    .Y(_09652_));
 AOI21x1_ASAP7_75t_R _17834_ (.A1(_08890_),
    .A2(_09645_),
    .B(_09652_),
    .Y(_09653_));
 INVx1_ASAP7_75t_R _17835_ (.A(_01020_),
    .Y(_09654_));
 AO21x2_ASAP7_75t_R _17836_ (.A1(_08877_),
    .A2(_08872_),
    .B(_09654_),
    .Y(_09655_));
 AND2x2_ASAP7_75t_L _17837_ (.A(_09655_),
    .B(_08885_),
    .Y(_09656_));
 NAND2x1_ASAP7_75t_R _17838_ (.A(_08879_),
    .B(_08866_),
    .Y(_09657_));
 AO21x1_ASAP7_75t_SL _17841_ (.A1(_09642_),
    .A2(_09657_),
    .B(_09572_),
    .Y(_09660_));
 AO21x1_ASAP7_75t_R _17842_ (.A1(_09560_),
    .A2(_09656_),
    .B(_09660_),
    .Y(_09661_));
 AO21x1_ASAP7_75t_R _17844_ (.A1(_08879_),
    .A2(_01023_),
    .B(_08884_),
    .Y(_09663_));
 OAI21x1_ASAP7_75t_R _17845_ (.A1(_08879_),
    .A2(_09557_),
    .B(_08884_),
    .Y(_09664_));
 OA21x2_ASAP7_75t_R _17846_ (.A1(_09641_),
    .A2(_09663_),
    .B(_09664_),
    .Y(_09665_));
 AOI21x1_ASAP7_75t_R _17848_ (.A1(_09572_),
    .A2(_09665_),
    .B(_09584_),
    .Y(_09667_));
 AO21x1_ASAP7_75t_R _17849_ (.A1(_09661_),
    .A2(_09667_),
    .B(_08902_),
    .Y(_09668_));
 AOI21x1_ASAP7_75t_SL _17851_ (.A1(_09639_),
    .A2(_09590_),
    .B(_08885_),
    .Y(_09670_));
 OA21x2_ASAP7_75t_R _17852_ (.A1(_08879_),
    .A2(_01025_),
    .B(_08885_),
    .Y(_09671_));
 AO21x1_ASAP7_75t_R _17854_ (.A1(_09671_),
    .A2(_09657_),
    .B(_08890_),
    .Y(_09673_));
 INVx1_ASAP7_75t_R _17855_ (.A(_01027_),
    .Y(_09674_));
 AO21x1_ASAP7_75t_R _17856_ (.A1(_08877_),
    .A2(_08872_),
    .B(_09674_),
    .Y(_09675_));
 AO21x1_ASAP7_75t_R _17857_ (.A1(_09626_),
    .A2(_09675_),
    .B(_08885_),
    .Y(_09676_));
 AND2x2_ASAP7_75t_L _17858_ (.A(_09663_),
    .B(_08890_),
    .Y(_09677_));
 AOI21x1_ASAP7_75t_R _17859_ (.A1(_09676_),
    .A2(_09677_),
    .B(_09584_),
    .Y(_09678_));
 OAI21x1_ASAP7_75t_R _17860_ (.A1(_09670_),
    .A2(_09673_),
    .B(_09678_),
    .Y(_09679_));
 NOR2x1_ASAP7_75t_L _17861_ (.A(_09572_),
    .B(_09598_),
    .Y(_09680_));
 NOR2x1_ASAP7_75t_SL _17862_ (.A(_01026_),
    .B(_08878_),
    .Y(_09681_));
 INVx1_ASAP7_75t_R _17863_ (.A(_09681_),
    .Y(_09682_));
 AO21x1_ASAP7_75t_L _17864_ (.A1(_08877_),
    .A2(_08872_),
    .B(_01023_),
    .Y(_09683_));
 AO21x1_ASAP7_75t_L _17865_ (.A1(_09682_),
    .A2(_09683_),
    .B(_08885_),
    .Y(_09684_));
 AOI21x1_ASAP7_75t_R _17866_ (.A1(_09680_),
    .A2(_09684_),
    .B(_08894_),
    .Y(_09685_));
 OAI21x1_ASAP7_75t_R _17867_ (.A1(_08885_),
    .A2(_09683_),
    .B(_09648_),
    .Y(_09686_));
 AOI21x1_ASAP7_75t_R _17868_ (.A1(_09685_),
    .A2(_09686_),
    .B(_09635_),
    .Y(_09687_));
 AOI21x1_ASAP7_75t_SL _17871_ (.A1(_09687_),
    .A2(_09679_),
    .B(_08898_),
    .Y(_09690_));
 OAI21x1_ASAP7_75t_SL _17872_ (.A1(_09653_),
    .A2(_09668_),
    .B(_09690_),
    .Y(_09691_));
 NAND2x1_ASAP7_75t_SL _17873_ (.A(_09691_),
    .B(_09638_),
    .Y(_00016_));
 INVx1_ASAP7_75t_SL _17874_ (.A(_09663_),
    .Y(_09692_));
 NAND2x1_ASAP7_75t_R _17875_ (.A(_08878_),
    .B(_08871_),
    .Y(_09693_));
 AO21x1_ASAP7_75t_R _17876_ (.A1(_09692_),
    .A2(_09693_),
    .B(_09572_),
    .Y(_09694_));
 NAND2x1_ASAP7_75t_R _17877_ (.A(_08878_),
    .B(_09554_),
    .Y(_09695_));
 AND2x2_ASAP7_75t_R _17878_ (.A(_09576_),
    .B(_09695_),
    .Y(_09696_));
 NOR3x1_ASAP7_75t_R _17879_ (.A(_09694_),
    .B(_09696_),
    .C(_08894_),
    .Y(_09697_));
 AO21x1_ASAP7_75t_R _17881_ (.A1(_01036_),
    .A2(_08885_),
    .B(_08890_),
    .Y(_09699_));
 NOR2x1_ASAP7_75t_R _17882_ (.A(_09646_),
    .B(_08878_),
    .Y(_09700_));
 INVx1_ASAP7_75t_SL _17883_ (.A(_09700_),
    .Y(_09701_));
 AO21x1_ASAP7_75t_R _17884_ (.A1(_08877_),
    .A2(_08872_),
    .B(_09605_),
    .Y(_09702_));
 AO21x1_ASAP7_75t_R _17885_ (.A1(_09701_),
    .A2(_09702_),
    .B(_08884_),
    .Y(_09703_));
 AND2x2_ASAP7_75t_R _17886_ (.A(_09570_),
    .B(_08884_),
    .Y(_09704_));
 NAND2x1_ASAP7_75t_R _17887_ (.A(_09704_),
    .B(_09657_),
    .Y(_09705_));
 AOI21x1_ASAP7_75t_R _17888_ (.A1(_09703_),
    .A2(_09705_),
    .B(_09572_),
    .Y(_09706_));
 AO21x2_ASAP7_75t_R _17889_ (.A1(_09701_),
    .A2(_09594_),
    .B(_08885_),
    .Y(_09707_));
 NOR2x1_ASAP7_75t_R _17890_ (.A(_08890_),
    .B(_09707_),
    .Y(_09708_));
 AOI211x1_ASAP7_75t_R _17891_ (.A1(_09584_),
    .A2(_09699_),
    .B(_09706_),
    .C(_09708_),
    .Y(_09709_));
 OAI21x1_ASAP7_75t_R _17892_ (.A1(_09697_),
    .A2(_09709_),
    .B(_08898_),
    .Y(_09710_));
 NOR2x1_ASAP7_75t_R _17893_ (.A(_09609_),
    .B(_09591_),
    .Y(_09711_));
 NAND2x1_ASAP7_75t_SL _17894_ (.A(_08878_),
    .B(_09557_),
    .Y(_09712_));
 OA21x2_ASAP7_75t_SL _17895_ (.A1(_09712_),
    .A2(_08885_),
    .B(_08890_),
    .Y(_09713_));
 NAND2x1_ASAP7_75t_R _17896_ (.A(_09630_),
    .B(_09713_),
    .Y(_09714_));
 NAND2x1_ASAP7_75t_R _17897_ (.A(_09693_),
    .B(_09692_),
    .Y(_09715_));
 AOI21x1_ASAP7_75t_R _17898_ (.A1(_09570_),
    .A2(_09576_),
    .B(_08890_),
    .Y(_09716_));
 AOI21x1_ASAP7_75t_R _17899_ (.A1(_09715_),
    .A2(_09716_),
    .B(_09584_),
    .Y(_09717_));
 OAI21x1_ASAP7_75t_R _17900_ (.A1(_09711_),
    .A2(_09714_),
    .B(_09717_),
    .Y(_09718_));
 INVx1_ASAP7_75t_R _17901_ (.A(_01028_),
    .Y(_09719_));
 OA21x2_ASAP7_75t_R _17902_ (.A1(_08879_),
    .A2(_09719_),
    .B(_08884_),
    .Y(_09720_));
 NAND2x1_ASAP7_75t_R _17903_ (.A(_09643_),
    .B(_09720_),
    .Y(_09721_));
 INVx2_ASAP7_75t_SL _17904_ (.A(_09588_),
    .Y(_09722_));
 NAND2x1_ASAP7_75t_R _17905_ (.A(_08885_),
    .B(_09562_),
    .Y(_09723_));
 INVx2_ASAP7_75t_R _17906_ (.A(_09723_),
    .Y(_09724_));
 NAND2x1_ASAP7_75t_R _17907_ (.A(_09722_),
    .B(_09724_),
    .Y(_09725_));
 NAND3x1_ASAP7_75t_R _17908_ (.A(_09721_),
    .B(_09725_),
    .C(_08890_),
    .Y(_09726_));
 NOR2x1_ASAP7_75t_R _17909_ (.A(_08890_),
    .B(_09598_),
    .Y(_09727_));
 AO21x1_ASAP7_75t_R _17910_ (.A1(_09712_),
    .A2(_09701_),
    .B(_08885_),
    .Y(_09728_));
 AOI21x1_ASAP7_75t_R _17911_ (.A1(_09727_),
    .A2(_09728_),
    .B(_08894_),
    .Y(_09729_));
 AOI21x1_ASAP7_75t_R _17912_ (.A1(_09726_),
    .A2(_09729_),
    .B(_08898_),
    .Y(_09730_));
 AOI21x1_ASAP7_75t_R _17913_ (.A1(_09718_),
    .A2(_09730_),
    .B(_08902_),
    .Y(_09731_));
 NAND2x1_ASAP7_75t_SL _17914_ (.A(_09710_),
    .B(_09731_),
    .Y(_09732_));
 NAND2x1_ASAP7_75t_R _17915_ (.A(_09557_),
    .B(_09554_),
    .Y(_09733_));
 AO21x1_ASAP7_75t_R _17917_ (.A1(_09733_),
    .A2(_09657_),
    .B(_08884_),
    .Y(_09735_));
 NAND2x1_ASAP7_75t_R _17919_ (.A(_09618_),
    .B(_09657_),
    .Y(_09737_));
 AND3x1_ASAP7_75t_R _17920_ (.A(_09735_),
    .B(_09572_),
    .C(_09737_),
    .Y(_09738_));
 NOR2x1_ASAP7_75t_SL _17921_ (.A(_08879_),
    .B(_08866_),
    .Y(_09739_));
 NOR2x1_ASAP7_75t_R _17922_ (.A(_08885_),
    .B(_09739_),
    .Y(_09740_));
 AOI22x1_ASAP7_75t_R _17923_ (.A1(_09598_),
    .A2(_09683_),
    .B1(_09740_),
    .B2(_09596_),
    .Y(_09741_));
 OAI21x1_ASAP7_75t_R _17924_ (.A1(_09572_),
    .A2(_09741_),
    .B(_09584_),
    .Y(_09742_));
 INVx1_ASAP7_75t_SL _17925_ (.A(_01023_),
    .Y(_09743_));
 NAND2x1_ASAP7_75t_R _17926_ (.A(_09743_),
    .B(_08879_),
    .Y(_09744_));
 OA21x2_ASAP7_75t_R _17927_ (.A1(_08885_),
    .A2(_09744_),
    .B(_09572_),
    .Y(_09745_));
 AOI21x1_ASAP7_75t_R _17928_ (.A1(_09725_),
    .A2(_09745_),
    .B(_09584_),
    .Y(_09746_));
 AOI21x1_ASAP7_75t_R _17929_ (.A1(_09656_),
    .A2(_09639_),
    .B(_09572_),
    .Y(_09747_));
 OAI21x1_ASAP7_75t_R _17930_ (.A1(_08885_),
    .A2(_09701_),
    .B(_09747_),
    .Y(_09748_));
 AOI21x1_ASAP7_75t_R _17931_ (.A1(_09746_),
    .A2(_09748_),
    .B(_08898_),
    .Y(_09749_));
 OAI21x1_ASAP7_75t_R _17932_ (.A1(_09738_),
    .A2(_09742_),
    .B(_09749_),
    .Y(_09750_));
 NAND2x1_ASAP7_75t_R _17933_ (.A(_09654_),
    .B(_08879_),
    .Y(_09751_));
 AO21x1_ASAP7_75t_R _17934_ (.A1(_09751_),
    .A2(_09617_),
    .B(_08884_),
    .Y(_09752_));
 INVx1_ASAP7_75t_R _17935_ (.A(_09752_),
    .Y(_09753_));
 AND2x2_ASAP7_75t_R _17936_ (.A(_09606_),
    .B(_08884_),
    .Y(_09754_));
 NOR2x1_ASAP7_75t_R _17937_ (.A(_08885_),
    .B(_09683_),
    .Y(_09755_));
 OR3x1_ASAP7_75t_R _17938_ (.A(_09754_),
    .B(_09755_),
    .C(_08890_),
    .Y(_09756_));
 AOI21x1_ASAP7_75t_SL _17939_ (.A1(_01030_),
    .A2(_08885_),
    .B(_09572_),
    .Y(_09757_));
 AO21x1_ASAP7_75t_R _17940_ (.A1(_09639_),
    .A2(_09683_),
    .B(_08885_),
    .Y(_09758_));
 AOI21x1_ASAP7_75t_R _17941_ (.A1(_09757_),
    .A2(_09758_),
    .B(_08894_),
    .Y(_09759_));
 OAI21x1_ASAP7_75t_R _17942_ (.A1(_09753_),
    .A2(_09756_),
    .B(_09759_),
    .Y(_09760_));
 NAND2x1_ASAP7_75t_R _17943_ (.A(_08878_),
    .B(_08866_),
    .Y(_09761_));
 OA21x2_ASAP7_75t_SL _17944_ (.A1(_08878_),
    .A2(_09743_),
    .B(_08884_),
    .Y(_09762_));
 AOI22x1_ASAP7_75t_R _17945_ (.A1(_09761_),
    .A2(_09598_),
    .B1(_09712_),
    .B2(_09762_),
    .Y(_09763_));
 NAND2x1_ASAP7_75t_R _17946_ (.A(_08890_),
    .B(_09763_),
    .Y(_09764_));
 OA21x2_ASAP7_75t_R _17947_ (.A1(_08884_),
    .A2(_09702_),
    .B(_09572_),
    .Y(_09765_));
 NAND2x1_ASAP7_75t_SL _17948_ (.A(_08879_),
    .B(_09554_),
    .Y(_09766_));
 NAND3x1_ASAP7_75t_R _17949_ (.A(_09575_),
    .B(_09766_),
    .C(_08884_),
    .Y(_09767_));
 AOI21x1_ASAP7_75t_R _17950_ (.A1(_09765_),
    .A2(_09767_),
    .B(_09584_),
    .Y(_09768_));
 AOI21x1_ASAP7_75t_R _17951_ (.A1(_09764_),
    .A2(_09768_),
    .B(_08899_),
    .Y(_09769_));
 AOI21x1_ASAP7_75t_R _17952_ (.A1(_09760_),
    .A2(_09769_),
    .B(_09635_),
    .Y(_09770_));
 NAND2x1_ASAP7_75t_SL _17953_ (.A(_09750_),
    .B(_09770_),
    .Y(_09771_));
 NAND2x1_ASAP7_75t_SL _17954_ (.A(_09732_),
    .B(_09771_),
    .Y(_00017_));
 NAND2x1_ASAP7_75t_SL _17955_ (.A(_08885_),
    .B(_09683_),
    .Y(_09772_));
 OAI21x1_ASAP7_75t_R _17956_ (.A1(_09606_),
    .A2(_09772_),
    .B(_09572_),
    .Y(_09773_));
 NOR2x1_ASAP7_75t_L _17957_ (.A(_09773_),
    .B(_09670_),
    .Y(_09774_));
 NAND2x1_ASAP7_75t_R _17958_ (.A(_09655_),
    .B(_09762_),
    .Y(_09775_));
 NOR2x1_ASAP7_75t_L _17959_ (.A(_08884_),
    .B(_09641_),
    .Y(_09776_));
 NAND2x1_ASAP7_75t_R _17960_ (.A(_09766_),
    .B(_09776_),
    .Y(_09777_));
 AOI21x1_ASAP7_75t_R _17961_ (.A1(_09775_),
    .A2(_09777_),
    .B(_09572_),
    .Y(_09778_));
 OAI21x1_ASAP7_75t_R _17962_ (.A1(_09774_),
    .A2(_09778_),
    .B(_09584_),
    .Y(_09779_));
 NOR2x1p5_ASAP7_75t_SL _17963_ (.A(_09588_),
    .B(_08885_),
    .Y(_09780_));
 AND2x2_ASAP7_75t_SL _17964_ (.A(_09780_),
    .B(_09693_),
    .Y(_09781_));
 AND2x2_ASAP7_75t_R _17965_ (.A(_08878_),
    .B(_09719_),
    .Y(_09782_));
 AOI211x1_ASAP7_75t_R _17966_ (.A1(_09557_),
    .A2(_08879_),
    .B(_08884_),
    .C(_09782_),
    .Y(_09783_));
 OAI21x1_ASAP7_75t_R _17967_ (.A1(_09781_),
    .A2(_09783_),
    .B(_08890_),
    .Y(_09784_));
 AOI21x1_ASAP7_75t_R _17968_ (.A1(_09643_),
    .A2(_09724_),
    .B(_09642_),
    .Y(_09785_));
 AOI21x1_ASAP7_75t_R _17969_ (.A1(_09572_),
    .A2(_09785_),
    .B(_09584_),
    .Y(_09786_));
 NAND2x1_ASAP7_75t_L _17970_ (.A(_09784_),
    .B(_09786_),
    .Y(_09787_));
 AOI21x1_ASAP7_75t_R _17971_ (.A1(_09787_),
    .A2(_09779_),
    .B(_08899_),
    .Y(_09788_));
 AO21x1_ASAP7_75t_R _17972_ (.A1(_08877_),
    .A2(_08872_),
    .B(_01020_),
    .Y(_09789_));
 NAND2x1_ASAP7_75t_SL _17973_ (.A(_08884_),
    .B(_09789_),
    .Y(_09790_));
 OAI21x1_ASAP7_75t_R _17974_ (.A1(_09681_),
    .A2(_09790_),
    .B(_08890_),
    .Y(_09791_));
 AOI21x1_ASAP7_75t_R _17975_ (.A1(_09557_),
    .A2(_08879_),
    .B(_09772_),
    .Y(_09792_));
 NOR2x1_ASAP7_75t_R _17976_ (.A(_09791_),
    .B(_09792_),
    .Y(_09793_));
 AO21x2_ASAP7_75t_SL _17977_ (.A1(_08877_),
    .A2(_08872_),
    .B(_09743_),
    .Y(_09794_));
 AND2x2_ASAP7_75t_R _17978_ (.A(_09794_),
    .B(_08885_),
    .Y(_09795_));
 NAND2x1_ASAP7_75t_R _17979_ (.A(_09795_),
    .B(_09639_),
    .Y(_09796_));
 AOI21x1_ASAP7_75t_R _17980_ (.A1(_09684_),
    .A2(_09796_),
    .B(_08890_),
    .Y(_09797_));
 OAI21x1_ASAP7_75t_R _17981_ (.A1(_09793_),
    .A2(_09797_),
    .B(_09584_),
    .Y(_09798_));
 AO21x1_ASAP7_75t_SL _17982_ (.A1(_09590_),
    .A2(_09722_),
    .B(_08884_),
    .Y(_09799_));
 AOI21x1_ASAP7_75t_R _17983_ (.A1(_01026_),
    .A2(_08878_),
    .B(_08885_),
    .Y(_09800_));
 NAND2x1_ASAP7_75t_R _17984_ (.A(_09800_),
    .B(_09657_),
    .Y(_09801_));
 AOI21x1_ASAP7_75t_R _17985_ (.A1(_09799_),
    .A2(_09801_),
    .B(_08890_),
    .Y(_09802_));
 OAI21x1_ASAP7_75t_R _17987_ (.A1(_08878_),
    .A2(_08866_),
    .B(_09789_),
    .Y(_09804_));
 NAND2x1_ASAP7_75t_R _17988_ (.A(_08884_),
    .B(_09804_),
    .Y(_09805_));
 OAI21x1_ASAP7_75t_R _17989_ (.A1(_09681_),
    .A2(_09649_),
    .B(_08885_),
    .Y(_09806_));
 AOI21x1_ASAP7_75t_R _17990_ (.A1(_09805_),
    .A2(_09806_),
    .B(_09572_),
    .Y(_09807_));
 OAI21x1_ASAP7_75t_SL _17991_ (.A1(_09807_),
    .A2(_09802_),
    .B(_08894_),
    .Y(_09808_));
 AOI21x1_ASAP7_75t_SL _17992_ (.A1(_09808_),
    .A2(_09798_),
    .B(_08898_),
    .Y(_09809_));
 OAI21x1_ASAP7_75t_R _17993_ (.A1(_09788_),
    .A2(_09809_),
    .B(_09635_),
    .Y(_09810_));
 NAND2x1_ASAP7_75t_R _17994_ (.A(_01034_),
    .B(_08885_),
    .Y(_09811_));
 OAI21x1_ASAP7_75t_R _17995_ (.A1(_08885_),
    .A2(_09641_),
    .B(_09811_),
    .Y(_09812_));
 OA21x2_ASAP7_75t_R _17996_ (.A1(_01032_),
    .A2(_08885_),
    .B(_08890_),
    .Y(_09813_));
 AOI21x1_ASAP7_75t_R _17997_ (.A1(_09813_),
    .A2(_09777_),
    .B(_08894_),
    .Y(_09814_));
 OAI21x1_ASAP7_75t_R _17998_ (.A1(_08890_),
    .A2(_09812_),
    .B(_09814_),
    .Y(_09815_));
 NAND2x1p5_ASAP7_75t_L _17999_ (.A(_09794_),
    .B(_09598_),
    .Y(_09816_));
 OR3x1_ASAP7_75t_R _18000_ (.A(_08885_),
    .B(_09674_),
    .C(_08878_),
    .Y(_09817_));
 AOI21x1_ASAP7_75t_SL _18001_ (.A1(_09817_),
    .A2(_09816_),
    .B(_08890_),
    .Y(_09818_));
 NAND2x1_ASAP7_75t_R _18002_ (.A(_09724_),
    .B(_09578_),
    .Y(_09819_));
 AOI21x1_ASAP7_75t_R _18003_ (.A1(_09707_),
    .A2(_09819_),
    .B(_09572_),
    .Y(_09820_));
 OAI21x1_ASAP7_75t_R _18004_ (.A1(_09818_),
    .A2(_09820_),
    .B(_08894_),
    .Y(_09821_));
 AOI21x1_ASAP7_75t_SL _18005_ (.A1(_09821_),
    .A2(_09815_),
    .B(_08899_),
    .Y(_09822_));
 NOR2x1_ASAP7_75t_R _18006_ (.A(_01022_),
    .B(_08878_),
    .Y(_09823_));
 OR2x2_ASAP7_75t_SL _18007_ (.A(_08885_),
    .B(_01035_),
    .Y(_09824_));
 OA21x2_ASAP7_75t_SL _18008_ (.A1(_09823_),
    .A2(_09591_),
    .B(_09824_),
    .Y(_09825_));
 NOR2x1p5_ASAP7_75t_L _18009_ (.A(_08890_),
    .B(_09825_),
    .Y(_09826_));
 OAI21x1_ASAP7_75t_R _18010_ (.A1(_08878_),
    .A2(_08866_),
    .B(_01032_),
    .Y(_09827_));
 NAND2x1_ASAP7_75t_R _18011_ (.A(_08885_),
    .B(_09827_),
    .Y(_09828_));
 INVx2_ASAP7_75t_SL _18012_ (.A(_09590_),
    .Y(_09829_));
 NOR2x1_ASAP7_75t_SL _18013_ (.A(_08878_),
    .B(_09554_),
    .Y(_09830_));
 OAI21x1_ASAP7_75t_R _18014_ (.A1(_09829_),
    .A2(_09830_),
    .B(_08884_),
    .Y(_09831_));
 AOI21x1_ASAP7_75t_R _18015_ (.A1(_09828_),
    .A2(_09831_),
    .B(_09572_),
    .Y(_09832_));
 OAI21x1_ASAP7_75t_SL _18016_ (.A1(_09832_),
    .A2(_09826_),
    .B(_08894_),
    .Y(_09833_));
 NAND2x1_ASAP7_75t_R _18017_ (.A(_01025_),
    .B(_08879_),
    .Y(_09834_));
 AO21x1_ASAP7_75t_R _18018_ (.A1(_09834_),
    .A2(_09617_),
    .B(_08884_),
    .Y(_09835_));
 OAI21x1_ASAP7_75t_R _18019_ (.A1(_08878_),
    .A2(_08871_),
    .B(_09675_),
    .Y(_09836_));
 AOI21x1_ASAP7_75t_R _18020_ (.A1(_08884_),
    .A2(_09836_),
    .B(_09572_),
    .Y(_09837_));
 AOI21x1_ASAP7_75t_R _18021_ (.A1(_09835_),
    .A2(_09837_),
    .B(_08894_),
    .Y(_09838_));
 NAND2x1_ASAP7_75t_R _18022_ (.A(_01036_),
    .B(_08884_),
    .Y(_09839_));
 OA21x2_ASAP7_75t_R _18023_ (.A1(_08871_),
    .A2(_08878_),
    .B(_08885_),
    .Y(_09840_));
 AOI21x1_ASAP7_75t_R _18024_ (.A1(_09575_),
    .A2(_09840_),
    .B(_08890_),
    .Y(_09841_));
 NAND2x1_ASAP7_75t_R _18025_ (.A(_09839_),
    .B(_09841_),
    .Y(_09842_));
 NAND2x1_ASAP7_75t_R _18026_ (.A(_09838_),
    .B(_09842_),
    .Y(_09843_));
 AOI21x1_ASAP7_75t_SL _18027_ (.A1(_09843_),
    .A2(_09833_),
    .B(_08898_),
    .Y(_09844_));
 OAI21x1_ASAP7_75t_SL _18028_ (.A1(_09844_),
    .A2(_09822_),
    .B(_08902_),
    .Y(_09845_));
 NAND2x1_ASAP7_75t_SL _18029_ (.A(_09810_),
    .B(_09845_),
    .Y(_00018_));
 AND3x1_ASAP7_75t_R _18030_ (.A(_09643_),
    .B(_08885_),
    .C(_09794_),
    .Y(_09846_));
 AO21x1_ASAP7_75t_R _18031_ (.A1(_09693_),
    .A2(_09780_),
    .B(_08890_),
    .Y(_09847_));
 NAND2x1_ASAP7_75t_R _18032_ (.A(_09596_),
    .B(_08890_),
    .Y(_09848_));
 OAI21x1_ASAP7_75t_R _18033_ (.A1(_09591_),
    .A2(_09848_),
    .B(_08894_),
    .Y(_09849_));
 NAND2x1_ASAP7_75t_R _18034_ (.A(_08884_),
    .B(_08890_),
    .Y(_09850_));
 AOI21x1_ASAP7_75t_R _18035_ (.A1(_09761_),
    .A2(_09566_),
    .B(_09850_),
    .Y(_09851_));
 NOR2x1_ASAP7_75t_SL _18036_ (.A(_09849_),
    .B(_09851_),
    .Y(_09852_));
 OAI21x1_ASAP7_75t_SL _18037_ (.A1(_09846_),
    .A2(_09847_),
    .B(_09852_),
    .Y(_09853_));
 AO21x1_ASAP7_75t_R _18038_ (.A1(_08871_),
    .A2(_08878_),
    .B(_08884_),
    .Y(_09854_));
 NOR2x1_ASAP7_75t_R _18039_ (.A(_09557_),
    .B(_09554_),
    .Y(_09855_));
 OAI21x1_ASAP7_75t_R _18040_ (.A1(_09739_),
    .A2(_09855_),
    .B(_08884_),
    .Y(_09856_));
 OAI21x1_ASAP7_75t_R _18041_ (.A1(_09559_),
    .A2(_09854_),
    .B(_09856_),
    .Y(_09857_));
 NAND2x1_ASAP7_75t_R _18042_ (.A(_08884_),
    .B(_09827_),
    .Y(_09858_));
 AOI21x1_ASAP7_75t_SL _18043_ (.A1(_09858_),
    .A2(_09592_),
    .B(_08894_),
    .Y(_09859_));
 OAI21x1_ASAP7_75t_SL _18044_ (.A1(_08890_),
    .A2(_09857_),
    .B(_09859_),
    .Y(_09860_));
 AOI21x1_ASAP7_75t_SL _18045_ (.A1(_09860_),
    .A2(_09853_),
    .B(_08899_),
    .Y(_09861_));
 INVx1_ASAP7_75t_SL _18046_ (.A(_09776_),
    .Y(_09862_));
 NAND2x1_ASAP7_75t_R _18047_ (.A(_09862_),
    .B(_09856_),
    .Y(_09863_));
 NAND2x1_ASAP7_75t_L _18048_ (.A(_09722_),
    .B(_09800_),
    .Y(_09864_));
 AOI21x1_ASAP7_75t_R _18049_ (.A1(_09864_),
    .A2(_09747_),
    .B(_08894_),
    .Y(_09865_));
 OAI21x1_ASAP7_75t_R _18050_ (.A1(_08890_),
    .A2(_09863_),
    .B(_09865_),
    .Y(_09866_));
 OA21x2_ASAP7_75t_SL _18051_ (.A1(_08878_),
    .A2(_01018_),
    .B(_08884_),
    .Y(_09867_));
 NAND2x1_ASAP7_75t_R _18052_ (.A(_09590_),
    .B(_09867_),
    .Y(_09868_));
 AO21x1_ASAP7_75t_R _18053_ (.A1(_09834_),
    .A2(_09702_),
    .B(_08884_),
    .Y(_09869_));
 AOI21x1_ASAP7_75t_R _18054_ (.A1(_09868_),
    .A2(_09869_),
    .B(_08890_),
    .Y(_09870_));
 AO21x1_ASAP7_75t_SL _18055_ (.A1(_09594_),
    .A2(_09560_),
    .B(_08885_),
    .Y(_09871_));
 NOR2x1_ASAP7_75t_R _18056_ (.A(_08871_),
    .B(_09557_),
    .Y(_09872_));
 OAI21x1_ASAP7_75t_R _18057_ (.A1(_09739_),
    .A2(_09872_),
    .B(_08885_),
    .Y(_09873_));
 AOI21x1_ASAP7_75t_R _18058_ (.A1(_09871_),
    .A2(_09873_),
    .B(_09572_),
    .Y(_09874_));
 OAI21x1_ASAP7_75t_R _18059_ (.A1(_09870_),
    .A2(_09874_),
    .B(_08894_),
    .Y(_09875_));
 AOI21x1_ASAP7_75t_R _18060_ (.A1(_09866_),
    .A2(_09875_),
    .B(_08898_),
    .Y(_09876_));
 OAI21x1_ASAP7_75t_SL _18061_ (.A1(_09861_),
    .A2(_09876_),
    .B(_08902_),
    .Y(_09877_));
 NAND2x1_ASAP7_75t_R _18062_ (.A(_09656_),
    .B(_09578_),
    .Y(_09878_));
 AO21x1_ASAP7_75t_SL _18063_ (.A1(_09722_),
    .A2(_09712_),
    .B(_08885_),
    .Y(_09879_));
 AOI21x1_ASAP7_75t_SL _18064_ (.A1(_09878_),
    .A2(_09879_),
    .B(_08894_),
    .Y(_09880_));
 AOI22x1_ASAP7_75t_R _18065_ (.A1(_08885_),
    .A2(_09681_),
    .B1(_09657_),
    .B2(_09800_),
    .Y(_09881_));
 OAI21x1_ASAP7_75t_R _18066_ (.A1(_09584_),
    .A2(_09881_),
    .B(_09572_),
    .Y(_09882_));
 NOR2x1_ASAP7_75t_L _18067_ (.A(_09880_),
    .B(_09882_),
    .Y(_09883_));
 AND2x2_ASAP7_75t_SL _18068_ (.A(_08884_),
    .B(_09559_),
    .Y(_09884_));
 INVx1_ASAP7_75t_R _18069_ (.A(_09884_),
    .Y(_09885_));
 OAI21x1_ASAP7_75t_R _18070_ (.A1(_09584_),
    .A2(_09885_),
    .B(_09628_),
    .Y(_09886_));
 NAND2x1_ASAP7_75t_R _18071_ (.A(_08885_),
    .B(_09829_),
    .Y(_09887_));
 AO21x1_ASAP7_75t_R _18072_ (.A1(_09639_),
    .A2(_09594_),
    .B(_08885_),
    .Y(_09888_));
 AOI21x1_ASAP7_75t_R _18073_ (.A1(_09887_),
    .A2(_09888_),
    .B(_08894_),
    .Y(_09889_));
 OAI21x1_ASAP7_75t_R _18074_ (.A1(_09889_),
    .A2(_09886_),
    .B(_08898_),
    .Y(_09890_));
 NOR2x1_ASAP7_75t_SL _18075_ (.A(_09883_),
    .B(_09890_),
    .Y(_09891_));
 NAND2x1_ASAP7_75t_SL _18076_ (.A(_09613_),
    .B(_09767_),
    .Y(_09892_));
 OAI21x1_ASAP7_75t_SL _18077_ (.A1(_09681_),
    .A2(_09604_),
    .B(_08885_),
    .Y(_09893_));
 AO21x1_ASAP7_75t_SL _18078_ (.A1(_09789_),
    .A2(_09722_),
    .B(_08885_),
    .Y(_09894_));
 NAND3x1_ASAP7_75t_L _18079_ (.A(_09893_),
    .B(_08890_),
    .C(_09894_),
    .Y(_09895_));
 AOI21x1_ASAP7_75t_R _18080_ (.A1(_09892_),
    .A2(_09895_),
    .B(_09584_),
    .Y(_09896_));
 AO21x1_ASAP7_75t_R _18081_ (.A1(_09657_),
    .A2(_09631_),
    .B(_08884_),
    .Y(_09897_));
 AOI21x1_ASAP7_75t_R _18082_ (.A1(_09707_),
    .A2(_09897_),
    .B(_08890_),
    .Y(_09898_));
 AO21x1_ASAP7_75t_R _18083_ (.A1(_09576_),
    .A2(_09789_),
    .B(_09572_),
    .Y(_09899_));
 NAND2x1_ASAP7_75t_R _18084_ (.A(_09584_),
    .B(_09899_),
    .Y(_09900_));
 OAI21x1_ASAP7_75t_R _18085_ (.A1(_09898_),
    .A2(_09900_),
    .B(_08899_),
    .Y(_09901_));
 NOR2x1_ASAP7_75t_SL _18086_ (.A(_09896_),
    .B(_09901_),
    .Y(_09902_));
 OAI21x1_ASAP7_75t_SL _18087_ (.A1(_09891_),
    .A2(_09902_),
    .B(_09635_),
    .Y(_09903_));
 NAND2x1_ASAP7_75t_SL _18088_ (.A(_09903_),
    .B(_09877_),
    .Y(_00019_));
 NOR2x1_ASAP7_75t_R _18089_ (.A(_09609_),
    .B(_09854_),
    .Y(_09904_));
 OAI21x1_ASAP7_75t_R _18090_ (.A1(_09904_),
    .A2(_09756_),
    .B(_08898_),
    .Y(_09905_));
 AO21x1_ASAP7_75t_R _18091_ (.A1(_08879_),
    .A2(_09605_),
    .B(_08884_),
    .Y(_09906_));
 OA211x2_ASAP7_75t_R _18092_ (.A1(_09649_),
    .A2(_09906_),
    .B(_09775_),
    .C(_08890_),
    .Y(_09907_));
 OAI21x1_ASAP7_75t_R _18093_ (.A1(_09905_),
    .A2(_09907_),
    .B(_08902_),
    .Y(_09908_));
 AND3x1_ASAP7_75t_SL _18094_ (.A(_09575_),
    .B(_08885_),
    .C(_09766_),
    .Y(_09909_));
 OAI21x1_ASAP7_75t_R _18095_ (.A1(_09696_),
    .A2(_09909_),
    .B(_09572_),
    .Y(_09910_));
 AO21x1_ASAP7_75t_R _18096_ (.A1(_09639_),
    .A2(_09570_),
    .B(_08884_),
    .Y(_09911_));
 NOR2x1_ASAP7_75t_R _18097_ (.A(_08866_),
    .B(_08871_),
    .Y(_09912_));
 OA21x2_ASAP7_75t_R _18098_ (.A1(_09912_),
    .A2(_09830_),
    .B(_08884_),
    .Y(_09913_));
 NOR2x1_ASAP7_75t_R _18099_ (.A(_09572_),
    .B(_09913_),
    .Y(_09914_));
 NAND2x1_ASAP7_75t_R _18100_ (.A(_09911_),
    .B(_09914_),
    .Y(_09915_));
 AOI21x1_ASAP7_75t_R _18101_ (.A1(_09910_),
    .A2(_09915_),
    .B(_08898_),
    .Y(_09916_));
 NOR2x1_ASAP7_75t_R _18102_ (.A(_09908_),
    .B(_09916_),
    .Y(_09917_));
 AND3x1_ASAP7_75t_R _18103_ (.A(_09695_),
    .B(_08884_),
    .C(_09610_),
    .Y(_09918_));
 NOR2x1_ASAP7_75t_R _18104_ (.A(_09918_),
    .B(_09694_),
    .Y(_09919_));
 AO21x1_ASAP7_75t_R _18105_ (.A1(_08878_),
    .A2(_08885_),
    .B(_08890_),
    .Y(_09920_));
 AO21x1_ASAP7_75t_R _18106_ (.A1(_09655_),
    .A2(_09576_),
    .B(_09920_),
    .Y(_09921_));
 NAND2x1_ASAP7_75t_R _18107_ (.A(_08899_),
    .B(_09921_),
    .Y(_09922_));
 OAI21x1_ASAP7_75t_R _18108_ (.A1(_09919_),
    .A2(_09922_),
    .B(_09635_),
    .Y(_09923_));
 AND3x1_ASAP7_75t_R _18109_ (.A(_09581_),
    .B(_09572_),
    .C(_09676_),
    .Y(_09924_));
 NAND2x1_ASAP7_75t_R _18110_ (.A(_08890_),
    .B(_09897_),
    .Y(_09925_));
 OAI21x1_ASAP7_75t_R _18111_ (.A1(_09913_),
    .A2(_09925_),
    .B(_08898_),
    .Y(_09926_));
 NOR2x1_ASAP7_75t_R _18112_ (.A(_09924_),
    .B(_09926_),
    .Y(_09927_));
 OAI21x1_ASAP7_75t_R _18113_ (.A1(_09923_),
    .A2(_09927_),
    .B(_09584_),
    .Y(_09928_));
 AO21x1_ASAP7_75t_SL _18114_ (.A1(_01026_),
    .A2(_08878_),
    .B(_08884_),
    .Y(_09929_));
 AND3x1_ASAP7_75t_SL _18115_ (.A(_09929_),
    .B(_08890_),
    .C(_09626_),
    .Y(_09930_));
 NOR2x1_ASAP7_75t_R _18116_ (.A(_08898_),
    .B(_09930_),
    .Y(_09931_));
 OR3x1_ASAP7_75t_R _18117_ (.A(_08866_),
    .B(_08878_),
    .C(_08884_),
    .Y(_09932_));
 OA21x2_ASAP7_75t_R _18118_ (.A1(_01037_),
    .A2(_08884_),
    .B(_09572_),
    .Y(_09933_));
 NAND3x1_ASAP7_75t_R _18119_ (.A(_09932_),
    .B(_09933_),
    .C(_09705_),
    .Y(_09934_));
 AOI21x1_ASAP7_75t_R _18120_ (.A1(_09931_),
    .A2(_09934_),
    .B(_09635_),
    .Y(_09935_));
 OA21x2_ASAP7_75t_R _18121_ (.A1(_09682_),
    .A2(_08884_),
    .B(_08890_),
    .Y(_09936_));
 OR2x2_ASAP7_75t_SL _18122_ (.A(_09617_),
    .B(_08884_),
    .Y(_09937_));
 NAND3x1_ASAP7_75t_R _18123_ (.A(_09936_),
    .B(_09684_),
    .C(_09937_),
    .Y(_09938_));
 AO21x1_ASAP7_75t_R _18124_ (.A1(_09751_),
    .A2(_09617_),
    .B(_08885_),
    .Y(_09939_));
 AOI21x1_ASAP7_75t_R _18125_ (.A1(_09939_),
    .A2(_09633_),
    .B(_08899_),
    .Y(_09940_));
 NAND2x1_ASAP7_75t_SL _18126_ (.A(_09938_),
    .B(_09940_),
    .Y(_09941_));
 NAND2x1_ASAP7_75t_R _18127_ (.A(_09935_),
    .B(_09941_),
    .Y(_09942_));
 NAND2x1_ASAP7_75t_R _18128_ (.A(_09617_),
    .B(_09762_),
    .Y(_09943_));
 NAND2x1_ASAP7_75t_R _18129_ (.A(_08890_),
    .B(_09723_),
    .Y(_09944_));
 OAI21x1_ASAP7_75t_R _18130_ (.A1(_09720_),
    .A2(_09944_),
    .B(_08899_),
    .Y(_09945_));
 AO21x1_ASAP7_75t_R _18131_ (.A1(_09648_),
    .A2(_09943_),
    .B(_09945_),
    .Y(_09946_));
 OAI21x1_ASAP7_75t_R _18132_ (.A1(_01018_),
    .A2(_08885_),
    .B(_09937_),
    .Y(_09947_));
 AOI21x1_ASAP7_75t_R _18133_ (.A1(_09572_),
    .A2(_09947_),
    .B(_08899_),
    .Y(_09948_));
 INVx1_ASAP7_75t_R _18134_ (.A(_09754_),
    .Y(_09949_));
 OA21x2_ASAP7_75t_SL _18135_ (.A1(_09830_),
    .A2(_09929_),
    .B(_08890_),
    .Y(_09950_));
 NAND2x1_ASAP7_75t_R _18136_ (.A(_09949_),
    .B(_09950_),
    .Y(_09951_));
 AOI21x1_ASAP7_75t_R _18137_ (.A1(_09948_),
    .A2(_09951_),
    .B(_08902_),
    .Y(_09952_));
 AOI21x1_ASAP7_75t_R _18138_ (.A1(_09946_),
    .A2(_09952_),
    .B(_09584_),
    .Y(_09953_));
 NAND2x1_ASAP7_75t_L _18139_ (.A(_09942_),
    .B(_09953_),
    .Y(_09954_));
 OAI21x1_ASAP7_75t_SL _18140_ (.A1(_09917_),
    .A2(_09928_),
    .B(_09954_),
    .Y(_00020_));
 AO21x1_ASAP7_75t_SL _18141_ (.A1(_01022_),
    .A2(_08878_),
    .B(_09762_),
    .Y(_09955_));
 OA21x2_ASAP7_75t_R _18142_ (.A1(_08885_),
    .A2(_09559_),
    .B(_09572_),
    .Y(_09956_));
 AOI21x1_ASAP7_75t_SL _18143_ (.A1(_09956_),
    .A2(_09893_),
    .B(_08894_),
    .Y(_09957_));
 OAI21x1_ASAP7_75t_SL _18144_ (.A1(_09572_),
    .A2(_09955_),
    .B(_09957_),
    .Y(_09958_));
 AO21x1_ASAP7_75t_R _18145_ (.A1(_09623_),
    .A2(_09631_),
    .B(_08885_),
    .Y(_09959_));
 NAND2x1_ASAP7_75t_R _18146_ (.A(_09795_),
    .B(_09578_),
    .Y(_09960_));
 AOI21x1_ASAP7_75t_SL _18147_ (.A1(_09959_),
    .A2(_09960_),
    .B(_09572_),
    .Y(_09961_));
 AO21x1_ASAP7_75t_R _18148_ (.A1(_09744_),
    .A2(_09789_),
    .B(_08884_),
    .Y(_09962_));
 AOI21x1_ASAP7_75t_SL _18149_ (.A1(_09962_),
    .A2(_09650_),
    .B(_08890_),
    .Y(_09963_));
 OAI21x1_ASAP7_75t_SL _18150_ (.A1(_09961_),
    .A2(_09963_),
    .B(_08894_),
    .Y(_09964_));
 AOI21x1_ASAP7_75t_SL _18151_ (.A1(_09958_),
    .A2(_09964_),
    .B(_08898_),
    .Y(_09965_));
 AO21x1_ASAP7_75t_R _18152_ (.A1(_09557_),
    .A2(_08884_),
    .B(_08871_),
    .Y(_09966_));
 NAND2x1_ASAP7_75t_R _18153_ (.A(_08884_),
    .B(_09649_),
    .Y(_09967_));
 AOI21x1_ASAP7_75t_SL _18154_ (.A1(_09966_),
    .A2(_09967_),
    .B(_08890_),
    .Y(_09968_));
 AND3x1_ASAP7_75t_SL _18155_ (.A(_09701_),
    .B(_08885_),
    .C(_09594_),
    .Y(_09969_));
 OAI21x1_ASAP7_75t_SL _18156_ (.A1(_09912_),
    .A2(_09664_),
    .B(_08890_),
    .Y(_09970_));
 NOR2x1_ASAP7_75t_SL _18157_ (.A(_09969_),
    .B(_09970_),
    .Y(_09971_));
 OAI21x1_ASAP7_75t_SL _18158_ (.A1(_09968_),
    .A2(_09971_),
    .B(_08894_),
    .Y(_09972_));
 NAND2x1_ASAP7_75t_SL _18159_ (.A(_09766_),
    .B(_09720_),
    .Y(_09973_));
 AOI21x1_ASAP7_75t_SL _18160_ (.A1(_09937_),
    .A2(_09973_),
    .B(_09572_),
    .Y(_09974_));
 NAND2x1_ASAP7_75t_SL _18161_ (.A(_09675_),
    .B(_09598_),
    .Y(_09975_));
 AND3x1_ASAP7_75t_SL _18162_ (.A(_09975_),
    .B(_09572_),
    .C(_09790_),
    .Y(_09976_));
 OAI21x1_ASAP7_75t_SL _18163_ (.A1(_09974_),
    .A2(_09976_),
    .B(_09584_),
    .Y(_09977_));
 AOI21x1_ASAP7_75t_SL _18164_ (.A1(_09972_),
    .A2(_09977_),
    .B(_08899_),
    .Y(_09978_));
 NOR2x1_ASAP7_75t_SL _18165_ (.A(_09965_),
    .B(_09978_),
    .Y(_09979_));
 AND3x1_ASAP7_75t_SL _18166_ (.A(_09657_),
    .B(_08884_),
    .C(_09794_),
    .Y(_09980_));
 INVx1_ASAP7_75t_SL _18167_ (.A(_09648_),
    .Y(_09981_));
 NAND2x1_ASAP7_75t_SL _18168_ (.A(_09655_),
    .B(_09867_),
    .Y(_09982_));
 OA21x2_ASAP7_75t_SL _18169_ (.A1(_08884_),
    .A2(_09594_),
    .B(_08890_),
    .Y(_09983_));
 AOI21x1_ASAP7_75t_SL _18170_ (.A1(_09982_),
    .A2(_09983_),
    .B(_08894_),
    .Y(_09984_));
 OAI21x1_ASAP7_75t_SL _18171_ (.A1(_09980_),
    .A2(_09981_),
    .B(_09984_),
    .Y(_09985_));
 AOI21x1_ASAP7_75t_SL _18172_ (.A1(_09800_),
    .A2(_09639_),
    .B(_09572_),
    .Y(_09986_));
 OAI21x1_ASAP7_75t_SL _18173_ (.A1(_09559_),
    .A2(_09862_),
    .B(_09986_),
    .Y(_09987_));
 OA21x2_ASAP7_75t_SL _18174_ (.A1(_08866_),
    .A2(_08884_),
    .B(_09572_),
    .Y(_09988_));
 AOI21x1_ASAP7_75t_SL _18175_ (.A1(_09988_),
    .A2(_09577_),
    .B(_09584_),
    .Y(_09989_));
 NAND2x1_ASAP7_75t_SL _18176_ (.A(_09987_),
    .B(_09989_),
    .Y(_09990_));
 AOI21x1_ASAP7_75t_SL _18177_ (.A1(_09985_),
    .A2(_09990_),
    .B(_08898_),
    .Y(_09991_));
 OAI21x1_ASAP7_75t_SL _18178_ (.A1(_09755_),
    .A2(_09656_),
    .B(_08894_),
    .Y(_09992_));
 NAND2x1_ASAP7_75t_SL _18179_ (.A(_08890_),
    .B(_09992_),
    .Y(_09993_));
 NAND2x1_ASAP7_75t_SL _18180_ (.A(_09655_),
    .B(_09780_),
    .Y(_09994_));
 AO21x1_ASAP7_75t_SL _18181_ (.A1(_09722_),
    .A2(_09594_),
    .B(_08884_),
    .Y(_09995_));
 AOI21x1_ASAP7_75t_SL _18182_ (.A1(_09994_),
    .A2(_09995_),
    .B(_08894_),
    .Y(_09996_));
 OAI21x1_ASAP7_75t_SL _18183_ (.A1(_09993_),
    .A2(_09996_),
    .B(_08898_),
    .Y(_09997_));
 AO21x1_ASAP7_75t_SL _18184_ (.A1(_01025_),
    .A2(_08885_),
    .B(_09867_),
    .Y(_09998_));
 AND3x1_ASAP7_75t_SL _18185_ (.A(_09578_),
    .B(_08885_),
    .C(_08894_),
    .Y(_09999_));
 AO21x1_ASAP7_75t_SL _18186_ (.A1(_09642_),
    .A2(_09647_),
    .B(_08890_),
    .Y(_10000_));
 AOI211x1_ASAP7_75t_SL _18187_ (.A1(_09584_),
    .A2(_09998_),
    .B(_09999_),
    .C(_10000_),
    .Y(_10001_));
 NOR2x1_ASAP7_75t_SL _18188_ (.A(_09997_),
    .B(_10001_),
    .Y(_10002_));
 OAI21x1_ASAP7_75t_SL _18189_ (.A1(_09991_),
    .A2(_10002_),
    .B(_09635_),
    .Y(_10003_));
 OAI21x1_ASAP7_75t_SL _18190_ (.A1(_09635_),
    .A2(_09979_),
    .B(_10003_),
    .Y(_00021_));
 OA21x2_ASAP7_75t_R _18191_ (.A1(_09554_),
    .A2(_08885_),
    .B(_09572_),
    .Y(_10004_));
 AO21x1_ASAP7_75t_R _18192_ (.A1(_09733_),
    .A2(_09639_),
    .B(_08884_),
    .Y(_10005_));
 AOI21x1_ASAP7_75t_SL _18193_ (.A1(_10004_),
    .A2(_10005_),
    .B(_09584_),
    .Y(_10006_));
 INVx1_ASAP7_75t_R _18194_ (.A(_09782_),
    .Y(_10007_));
 OA21x2_ASAP7_75t_R _18195_ (.A1(_08884_),
    .A2(_10007_),
    .B(_09817_),
    .Y(_10008_));
 NAND2x1_ASAP7_75t_SL _18196_ (.A(_09936_),
    .B(_10008_),
    .Y(_10009_));
 AOI21x1_ASAP7_75t_SL _18197_ (.A1(_10006_),
    .A2(_10009_),
    .B(_08898_),
    .Y(_10010_));
 NAND2x1_ASAP7_75t_R _18198_ (.A(_09618_),
    .B(_09578_),
    .Y(_10011_));
 NAND3x1_ASAP7_75t_SL _18199_ (.A(_09893_),
    .B(_08890_),
    .C(_10011_),
    .Y(_10012_));
 AO21x1_ASAP7_75t_R _18200_ (.A1(_08877_),
    .A2(_08872_),
    .B(_09646_),
    .Y(_10013_));
 AO21x1_ASAP7_75t_R _18201_ (.A1(_09626_),
    .A2(_10013_),
    .B(_08884_),
    .Y(_10014_));
 AOI21x1_ASAP7_75t_R _18202_ (.A1(_09643_),
    .A2(_09800_),
    .B(_08890_),
    .Y(_10015_));
 NAND2x1_ASAP7_75t_SL _18203_ (.A(_10014_),
    .B(_10015_),
    .Y(_10016_));
 NAND3x1_ASAP7_75t_SL _18204_ (.A(_10012_),
    .B(_09584_),
    .C(_10016_),
    .Y(_10017_));
 NAND2x1_ASAP7_75t_SL _18205_ (.A(_10010_),
    .B(_10017_),
    .Y(_10018_));
 NAND2x1_ASAP7_75t_R _18206_ (.A(_09722_),
    .B(_09720_),
    .Y(_10019_));
 NAND2x1_ASAP7_75t_R _18207_ (.A(_09639_),
    .B(_09776_),
    .Y(_10020_));
 AOI21x1_ASAP7_75t_SL _18208_ (.A1(_10019_),
    .A2(_10020_),
    .B(_08890_),
    .Y(_10021_));
 AND3x1_ASAP7_75t_SL _18209_ (.A(_09812_),
    .B(_08890_),
    .C(_09885_),
    .Y(_10022_));
 OAI21x1_ASAP7_75t_SL _18210_ (.A1(_10021_),
    .A2(_10022_),
    .B(_08894_),
    .Y(_10023_));
 AOI21x1_ASAP7_75t_R _18211_ (.A1(_09618_),
    .A2(_09578_),
    .B(_08890_),
    .Y(_10024_));
 OAI21x1_ASAP7_75t_SL _18212_ (.A1(_09739_),
    .A2(_09906_),
    .B(_10024_),
    .Y(_10025_));
 OA21x2_ASAP7_75t_SL _18213_ (.A1(_08885_),
    .A2(_09594_),
    .B(_08890_),
    .Y(_10026_));
 AO21x1_ASAP7_75t_SL _18214_ (.A1(_09554_),
    .A2(_08878_),
    .B(_09906_),
    .Y(_10027_));
 AOI21x1_ASAP7_75t_SL _18215_ (.A1(_10026_),
    .A2(_10027_),
    .B(_08894_),
    .Y(_10028_));
 AOI21x1_ASAP7_75t_SL _18216_ (.A1(_10025_),
    .A2(_10028_),
    .B(_08899_),
    .Y(_10029_));
 AOI21x1_ASAP7_75t_SL _18217_ (.A1(_10023_),
    .A2(_10029_),
    .B(_09635_),
    .Y(_10030_));
 NAND2x1_ASAP7_75t_SL _18218_ (.A(_10018_),
    .B(_10030_),
    .Y(_10031_));
 AND2x2_ASAP7_75t_SL _18219_ (.A(_09643_),
    .B(_08884_),
    .Y(_10032_));
 AND3x1_ASAP7_75t_SL _18220_ (.A(_09575_),
    .B(_08885_),
    .C(_09712_),
    .Y(_10033_));
 AOI211x1_ASAP7_75t_SL _18221_ (.A1(_09712_),
    .A2(_10032_),
    .B(_10033_),
    .C(_09572_),
    .Y(_10034_));
 AND3x1_ASAP7_75t_SL _18222_ (.A(_09639_),
    .B(_08884_),
    .C(_09702_),
    .Y(_10035_));
 OAI21x1_ASAP7_75t_SL _18223_ (.A1(_10035_),
    .A2(_10033_),
    .B(_09572_),
    .Y(_10036_));
 NAND2x1_ASAP7_75t_SL _18224_ (.A(_08894_),
    .B(_10036_),
    .Y(_10037_));
 NOR2x1_ASAP7_75t_SL _18225_ (.A(_10034_),
    .B(_10037_),
    .Y(_10038_));
 NAND2x1_ASAP7_75t_SL _18226_ (.A(_08884_),
    .B(_09588_),
    .Y(_10039_));
 NAND3x1_ASAP7_75t_SL _18227_ (.A(_09893_),
    .B(_09572_),
    .C(_10039_),
    .Y(_10040_));
 NAND2x1_ASAP7_75t_SL _18228_ (.A(_09657_),
    .B(_09642_),
    .Y(_10041_));
 AOI21x1_ASAP7_75t_SL _18229_ (.A1(_09757_),
    .A2(_10041_),
    .B(_08894_),
    .Y(_10042_));
 AO21x1_ASAP7_75t_SL _18230_ (.A1(_10040_),
    .A2(_10042_),
    .B(_08898_),
    .Y(_10043_));
 AO21x1_ASAP7_75t_SL _18231_ (.A1(_09564_),
    .A2(_08878_),
    .B(_08885_),
    .Y(_10044_));
 NOR2x1_ASAP7_75t_SL _18232_ (.A(_09606_),
    .B(_09772_),
    .Y(_10045_));
 AO21x1_ASAP7_75t_SL _18233_ (.A1(_10045_),
    .A2(_09572_),
    .B(_08894_),
    .Y(_10046_));
 AO21x1_ASAP7_75t_SL _18234_ (.A1(_10044_),
    .A2(_09950_),
    .B(_10046_),
    .Y(_10047_));
 AOI21x1_ASAP7_75t_SL _18235_ (.A1(_01031_),
    .A2(_08885_),
    .B(_08890_),
    .Y(_10048_));
 NAND2x1_ASAP7_75t_SL _18236_ (.A(_09800_),
    .B(_09639_),
    .Y(_10049_));
 AOI21x1_ASAP7_75t_SL _18237_ (.A1(_10048_),
    .A2(_10049_),
    .B(_09584_),
    .Y(_10050_));
 NAND2x1_ASAP7_75t_SL _18238_ (.A(_09722_),
    .B(_09656_),
    .Y(_10051_));
 NAND2x1_ASAP7_75t_SL _18239_ (.A(_10051_),
    .B(_09713_),
    .Y(_10052_));
 AOI21x1_ASAP7_75t_SL _18240_ (.A1(_10050_),
    .A2(_10052_),
    .B(_08899_),
    .Y(_10053_));
 AOI21x1_ASAP7_75t_SL _18241_ (.A1(_10047_),
    .A2(_10053_),
    .B(_08902_),
    .Y(_10054_));
 OAI21x1_ASAP7_75t_SL _18242_ (.A1(_10038_),
    .A2(_10043_),
    .B(_10054_),
    .Y(_10055_));
 NAND2x1_ASAP7_75t_SL _18243_ (.A(_10031_),
    .B(_10055_),
    .Y(_00022_));
 AND3x1_ASAP7_75t_R _18244_ (.A(_09967_),
    .B(_08890_),
    .C(_09949_),
    .Y(_10056_));
 AO21x1_ASAP7_75t_R _18245_ (.A1(_01018_),
    .A2(_08885_),
    .B(_08890_),
    .Y(_10057_));
 AO21x1_ASAP7_75t_R _18246_ (.A1(_08884_),
    .A2(_09782_),
    .B(_10057_),
    .Y(_10058_));
 NAND2x1_ASAP7_75t_R _18247_ (.A(_08894_),
    .B(_10058_),
    .Y(_10059_));
 AOI21x1_ASAP7_75t_R _18248_ (.A1(_09715_),
    .A2(_10056_),
    .B(_10059_),
    .Y(_10060_));
 AO21x1_ASAP7_75t_R _18249_ (.A1(_09682_),
    .A2(_09590_),
    .B(_08885_),
    .Y(_10061_));
 OAI21x1_ASAP7_75t_R _18250_ (.A1(_01037_),
    .A2(_08884_),
    .B(_10061_),
    .Y(_10062_));
 OAI21x1_ASAP7_75t_R _18251_ (.A1(_08890_),
    .A2(_10062_),
    .B(_09584_),
    .Y(_10063_));
 AO21x1_ASAP7_75t_R _18252_ (.A1(_09560_),
    .A2(_09617_),
    .B(_08884_),
    .Y(_10064_));
 AND3x1_ASAP7_75t_R _18253_ (.A(_09713_),
    .B(_09824_),
    .C(_10064_),
    .Y(_10065_));
 OAI21x1_ASAP7_75t_R _18254_ (.A1(_10063_),
    .A2(_10065_),
    .B(_08898_),
    .Y(_10066_));
 NOR2x1_ASAP7_75t_R _18255_ (.A(_10060_),
    .B(_10066_),
    .Y(_10067_));
 AND3x1_ASAP7_75t_R _18256_ (.A(_09610_),
    .B(_08884_),
    .C(_09562_),
    .Y(_10068_));
 AO21x1_ASAP7_75t_R _18257_ (.A1(_09671_),
    .A2(_09722_),
    .B(_08890_),
    .Y(_10069_));
 OAI21x1_ASAP7_75t_R _18258_ (.A1(_10068_),
    .A2(_10069_),
    .B(_08894_),
    .Y(_10070_));
 AND3x1_ASAP7_75t_R _18259_ (.A(_09766_),
    .B(_08884_),
    .C(_09562_),
    .Y(_10071_));
 NOR2x1_ASAP7_75t_R _18260_ (.A(_10071_),
    .B(_09925_),
    .Y(_10072_));
 NOR2x1_ASAP7_75t_SL _18261_ (.A(_10070_),
    .B(_10072_),
    .Y(_10073_));
 AO21x1_ASAP7_75t_R _18262_ (.A1(_09695_),
    .A2(_08885_),
    .B(_09720_),
    .Y(_10074_));
 AOI21x1_ASAP7_75t_R _18263_ (.A1(_09610_),
    .A2(_10074_),
    .B(_08890_),
    .Y(_10075_));
 OA21x2_ASAP7_75t_R _18264_ (.A1(_01023_),
    .A2(_08885_),
    .B(_08890_),
    .Y(_10076_));
 AO21x1_ASAP7_75t_R _18265_ (.A1(_10005_),
    .A2(_10076_),
    .B(_08894_),
    .Y(_10077_));
 OAI21x1_ASAP7_75t_R _18266_ (.A1(_10075_),
    .A2(_10077_),
    .B(_08899_),
    .Y(_10078_));
 OAI21x1_ASAP7_75t_R _18267_ (.A1(_10073_),
    .A2(_10078_),
    .B(_08902_),
    .Y(_10079_));
 NAND2x1_ASAP7_75t_R _18268_ (.A(_09752_),
    .B(_09879_),
    .Y(_10080_));
 AOI21x1_ASAP7_75t_R _18269_ (.A1(_10015_),
    .A2(_09828_),
    .B(_08894_),
    .Y(_10081_));
 OAI21x1_ASAP7_75t_R _18270_ (.A1(_09572_),
    .A2(_10080_),
    .B(_10081_),
    .Y(_10082_));
 OA21x2_ASAP7_75t_R _18271_ (.A1(_09723_),
    .A2(_09609_),
    .B(_08890_),
    .Y(_10083_));
 OAI21x1_ASAP7_75t_R _18272_ (.A1(_09664_),
    .A2(_09823_),
    .B(_10083_),
    .Y(_10084_));
 NOR2x1_ASAP7_75t_R _18273_ (.A(_09929_),
    .B(_09830_),
    .Y(_10085_));
 AO21x1_ASAP7_75t_SL _18274_ (.A1(_09643_),
    .A2(_08884_),
    .B(_08890_),
    .Y(_10086_));
 OA21x2_ASAP7_75t_R _18275_ (.A1(_10085_),
    .A2(_10086_),
    .B(_08894_),
    .Y(_10087_));
 AOI21x1_ASAP7_75t_R _18276_ (.A1(_10084_),
    .A2(_10087_),
    .B(_08898_),
    .Y(_10088_));
 AOI21x1_ASAP7_75t_R _18277_ (.A1(_10082_),
    .A2(_10088_),
    .B(_08902_),
    .Y(_10089_));
 AO21x1_ASAP7_75t_R _18278_ (.A1(_09560_),
    .A2(_10013_),
    .B(_08885_),
    .Y(_10090_));
 AO21x1_ASAP7_75t_R _18279_ (.A1(_10090_),
    .A2(_09906_),
    .B(_09572_),
    .Y(_10091_));
 OAI21x1_ASAP7_75t_R _18280_ (.A1(_08884_),
    .A2(_09700_),
    .B(_09956_),
    .Y(_10092_));
 AO21x1_ASAP7_75t_R _18281_ (.A1(_10091_),
    .A2(_10092_),
    .B(_08894_),
    .Y(_10093_));
 OA21x2_ASAP7_75t_R _18282_ (.A1(_08866_),
    .A2(_08885_),
    .B(_08890_),
    .Y(_10094_));
 AO21x1_ASAP7_75t_R _18283_ (.A1(_09695_),
    .A2(_09657_),
    .B(_08884_),
    .Y(_10095_));
 AOI21x1_ASAP7_75t_R _18284_ (.A1(_10094_),
    .A2(_10095_),
    .B(_09584_),
    .Y(_10096_));
 AO21x1_ASAP7_75t_R _18285_ (.A1(_09766_),
    .A2(_10013_),
    .B(_08885_),
    .Y(_10097_));
 NAND2x1_ASAP7_75t_R _18286_ (.A(_10097_),
    .B(_09841_),
    .Y(_10098_));
 AOI21x1_ASAP7_75t_R _18287_ (.A1(_10096_),
    .A2(_10098_),
    .B(_08899_),
    .Y(_10099_));
 NAND2x1_ASAP7_75t_R _18288_ (.A(_10093_),
    .B(_10099_),
    .Y(_10100_));
 NAND2x1_ASAP7_75t_SL _18289_ (.A(_10089_),
    .B(_10100_),
    .Y(_10101_));
 OAI21x1_ASAP7_75t_SL _18290_ (.A1(_10067_),
    .A2(_10079_),
    .B(_10101_),
    .Y(_00023_));
 XNOR2x2_ASAP7_75t_SL _18291_ (.A(_08769_),
    .B(_08947_),
    .Y(_10102_));
 AOI21x1_ASAP7_75t_SL _18292_ (.A1(_08005_),
    .A2(_10102_),
    .B(_08949_),
    .Y(_10103_));
 INVx3_ASAP7_75t_SL _18294_ (.A(_08958_),
    .Y(_10104_));
 INVx1_ASAP7_75t_R _18296_ (.A(_08942_),
    .Y(_10105_));
 INVx1_ASAP7_75t_R _18297_ (.A(_00886_),
    .Y(_10106_));
 XOR2x2_ASAP7_75t_R _18298_ (.A(_08684_),
    .B(_10106_),
    .Y(_10107_));
 OAI21x1_ASAP7_75t_R _18299_ (.A1(_10105_),
    .A2(_10107_),
    .B(_08005_),
    .Y(_10108_));
 INVx1_ASAP7_75t_R _18300_ (.A(_08946_),
    .Y(_10109_));
 OAI21x1_ASAP7_75t_R _18301_ (.A1(_08944_),
    .A2(_10108_),
    .B(_10109_),
    .Y(_10110_));
 NOR2x2_ASAP7_75t_SL _18305_ (.A(_01050_),
    .B(_08958_),
    .Y(_10113_));
 AOI21x1_ASAP7_75t_R _18306_ (.A1(_08960_),
    .A2(_08773_),
    .B(ld),
    .Y(_10114_));
 INVx1_ASAP7_75t_R _18307_ (.A(_08961_),
    .Y(_10115_));
 AOI21x1_ASAP7_75t_R _18308_ (.A1(_10114_),
    .A2(_10115_),
    .B(_08966_),
    .Y(_10116_));
 AND2x2_ASAP7_75t_SL _18311_ (.A(_10113_),
    .B(_10116_),
    .Y(_10119_));
 NAND2x2_ASAP7_75t_SL _18312_ (.A(_08958_),
    .B(_01048_),
    .Y(_10120_));
 INVx2_ASAP7_75t_R _18313_ (.A(_10120_),
    .Y(_10121_));
 OAI21x1_ASAP7_75t_SL _18315_ (.A1(_01044_),
    .A2(_08958_),
    .B(_08968_),
    .Y(_10123_));
 OAI21x1_ASAP7_75t_SL _18318_ (.A1(_10121_),
    .A2(_10123_),
    .B(_08975_),
    .Y(_10126_));
 OAI21x1_ASAP7_75t_SL _18319_ (.A1(_10119_),
    .A2(_10126_),
    .B(_08982_),
    .Y(_10127_));
 INVx2_ASAP7_75t_R _18320_ (.A(_01044_),
    .Y(_10128_));
 NOR2x2_ASAP7_75t_SL _18321_ (.A(_10128_),
    .B(_08958_),
    .Y(_10129_));
 AND2x2_ASAP7_75t_SL _18323_ (.A(_10129_),
    .B(_10116_),
    .Y(_10131_));
 NAND2x2_ASAP7_75t_SL _18325_ (.A(_01047_),
    .B(_08958_),
    .Y(_10133_));
 OAI21x1_ASAP7_75t_R _18326_ (.A1(_08968_),
    .A2(_10133_),
    .B(_08976_),
    .Y(_10134_));
 AOI211x1_ASAP7_75t_R _18327_ (.A1(_08968_),
    .A2(_10113_),
    .B(_10131_),
    .C(_10134_),
    .Y(_10135_));
 OAI21x1_ASAP7_75t_R _18330_ (.A1(_10127_),
    .A2(_10135_),
    .B(_08987_),
    .Y(_10138_));
 NAND2x2_ASAP7_75t_SL _18331_ (.A(_10110_),
    .B(_08958_),
    .Y(_10139_));
 OA21x2_ASAP7_75t_SL _18332_ (.A1(_08958_),
    .A2(_01044_),
    .B(_10116_),
    .Y(_10140_));
 NAND2x1_ASAP7_75t_R _18333_ (.A(_10139_),
    .B(_10140_),
    .Y(_10141_));
 INVx2_ASAP7_75t_SL _18335_ (.A(_01049_),
    .Y(_10143_));
 NOR2x2_ASAP7_75t_SL _18336_ (.A(_10143_),
    .B(_08958_),
    .Y(_10144_));
 INVx2_ASAP7_75t_SL _18337_ (.A(_10139_),
    .Y(_10145_));
 OAI21x1_ASAP7_75t_R _18339_ (.A1(_10144_),
    .A2(_10145_),
    .B(_08968_),
    .Y(_10147_));
 AND3x1_ASAP7_75t_SL _18340_ (.A(_10141_),
    .B(_08975_),
    .C(_10147_),
    .Y(_10148_));
 INVx1_ASAP7_75t_R _18341_ (.A(_08982_),
    .Y(_10149_));
 INVx2_ASAP7_75t_SL _18344_ (.A(_01041_),
    .Y(_10152_));
 NAND2x2_ASAP7_75t_SL _18345_ (.A(_08958_),
    .B(_10152_),
    .Y(_10153_));
 INVx3_ASAP7_75t_SL _18346_ (.A(_10153_),
    .Y(_10154_));
 INVx1_ASAP7_75t_R _18347_ (.A(_01054_),
    .Y(_10155_));
 AO21x1_ASAP7_75t_R _18348_ (.A1(_10155_),
    .A2(_08968_),
    .B(_08975_),
    .Y(_10156_));
 AO21x1_ASAP7_75t_SL _18349_ (.A1(_10154_),
    .A2(_10116_),
    .B(_10156_),
    .Y(_10157_));
 NAND2x1_ASAP7_75t_L _18350_ (.A(_10149_),
    .B(_10157_),
    .Y(_10158_));
 NOR2x1_ASAP7_75t_SL _18351_ (.A(_10148_),
    .B(_10158_),
    .Y(_10159_));
 OAI21x1_ASAP7_75t_SL _18352_ (.A1(_10159_),
    .A2(_10138_),
    .B(_08992_),
    .Y(_10160_));
 NOR2x2_ASAP7_75t_SL _18353_ (.A(_10152_),
    .B(_08958_),
    .Y(_10161_));
 NOR2x2_ASAP7_75t_SL _18354_ (.A(_10161_),
    .B(_10116_),
    .Y(_10162_));
 NOR2x1_ASAP7_75t_R _18355_ (.A(key[26]),
    .B(_08005_),
    .Y(_10163_));
 INVx1_ASAP7_75t_R _18356_ (.A(_10163_),
    .Y(_10164_));
 NOR2x1_ASAP7_75t_R _18357_ (.A(_08951_),
    .B(_08771_),
    .Y(_10165_));
 NOR2x1_ASAP7_75t_R _18358_ (.A(_08952_),
    .B(_08954_),
    .Y(_10166_));
 OAI21x1_ASAP7_75t_R _18359_ (.A1(_10165_),
    .A2(_10166_),
    .B(_08005_),
    .Y(_10167_));
 AOI21x1_ASAP7_75t_R _18361_ (.A1(_10164_),
    .A2(_10167_),
    .B(_01045_),
    .Y(_10169_));
 NOR2x2_ASAP7_75t_SL _18362_ (.A(_01048_),
    .B(_08958_),
    .Y(_10170_));
 OA21x2_ASAP7_75t_R _18363_ (.A1(_10169_),
    .A2(_10170_),
    .B(_10116_),
    .Y(_10171_));
 OAI21x1_ASAP7_75t_SL _18364_ (.A1(_10171_),
    .A2(_10162_),
    .B(_08976_),
    .Y(_10172_));
 INVx1_ASAP7_75t_R _18365_ (.A(_01045_),
    .Y(_10173_));
 NAND2x2_ASAP7_75t_SL _18366_ (.A(_10173_),
    .B(_08958_),
    .Y(_10174_));
 NOR2x1_ASAP7_75t_L _18367_ (.A(_08968_),
    .B(_10174_),
    .Y(_10175_));
 INVx1_ASAP7_75t_R _18368_ (.A(_01040_),
    .Y(_10176_));
 NOR2x2_ASAP7_75t_SL _18369_ (.A(_10176_),
    .B(_08958_),
    .Y(_10177_));
 OA21x2_ASAP7_75t_R _18370_ (.A1(_10145_),
    .A2(_10177_),
    .B(_08968_),
    .Y(_10178_));
 OAI21x1_ASAP7_75t_R _18372_ (.A1(_10175_),
    .A2(_10178_),
    .B(_08975_),
    .Y(_10180_));
 AOI21x1_ASAP7_75t_R _18373_ (.A1(_10172_),
    .A2(_10180_),
    .B(_08982_),
    .Y(_10181_));
 AOI21x1_ASAP7_75t_SL _18374_ (.A1(_10104_),
    .A2(_10103_),
    .B(_08968_),
    .Y(_10182_));
 NAND2x1p5_ASAP7_75t_L _18375_ (.A(_10153_),
    .B(_10182_),
    .Y(_10183_));
 INVx2_ASAP7_75t_R _18376_ (.A(_10183_),
    .Y(_10184_));
 INVx1_ASAP7_75t_R _18377_ (.A(_01047_),
    .Y(_10185_));
 AND2x2_ASAP7_75t_R _18378_ (.A(_08958_),
    .B(_10185_),
    .Y(_10186_));
 OA21x2_ASAP7_75t_R _18379_ (.A1(_08958_),
    .A2(_10110_),
    .B(_08968_),
    .Y(_10187_));
 INVx1_ASAP7_75t_SL _18380_ (.A(_10187_),
    .Y(_10188_));
 OAI21x1_ASAP7_75t_R _18381_ (.A1(_10186_),
    .A2(_10188_),
    .B(_08975_),
    .Y(_10189_));
 NOR2x1_ASAP7_75t_SL _18382_ (.A(_10184_),
    .B(_10189_),
    .Y(_10190_));
 NOR2x1_ASAP7_75t_SL _18384_ (.A(_10173_),
    .B(_08958_),
    .Y(_10192_));
 NOR2x1_ASAP7_75t_SL _18385_ (.A(_10116_),
    .B(_10192_),
    .Y(_10193_));
 NOR2x1_ASAP7_75t_R _18386_ (.A(_08975_),
    .B(_10193_),
    .Y(_10194_));
 AND2x2_ASAP7_75t_SL _18388_ (.A(_08958_),
    .B(_01049_),
    .Y(_10196_));
 OAI21x1_ASAP7_75t_SL _18389_ (.A1(_10113_),
    .A2(_10196_),
    .B(_10116_),
    .Y(_10197_));
 AO21x1_ASAP7_75t_SL _18390_ (.A1(_10194_),
    .A2(_10197_),
    .B(_10149_),
    .Y(_10198_));
 OAI21x1_ASAP7_75t_R _18391_ (.A1(_10190_),
    .A2(_10198_),
    .B(_08988_),
    .Y(_10199_));
 NOR2x1_ASAP7_75t_SL _18392_ (.A(_10181_),
    .B(_10199_),
    .Y(_10200_));
 NAND2x2_ASAP7_75t_SL _18393_ (.A(_10176_),
    .B(_08958_),
    .Y(_10201_));
 NOR2x2_ASAP7_75t_SL _18394_ (.A(_10161_),
    .B(_08968_),
    .Y(_10202_));
 NOR2x1_ASAP7_75t_SL _18395_ (.A(_10185_),
    .B(_08958_),
    .Y(_10203_));
 OA21x2_ASAP7_75t_SL _18396_ (.A1(_10196_),
    .A2(_10203_),
    .B(_08968_),
    .Y(_10204_));
 AOI21x1_ASAP7_75t_SL _18397_ (.A1(_10202_),
    .A2(_10201_),
    .B(_10204_),
    .Y(_10205_));
 AOI21x1_ASAP7_75t_SL _18398_ (.A1(_10110_),
    .A2(_10104_),
    .B(_08968_),
    .Y(_10206_));
 NAND2x1_ASAP7_75t_R _18399_ (.A(_01043_),
    .B(_01046_),
    .Y(_10207_));
 AND2x2_ASAP7_75t_SL _18400_ (.A(_10206_),
    .B(_10207_),
    .Y(_10208_));
 NOR2x1_ASAP7_75t_R _18401_ (.A(_10110_),
    .B(_01046_),
    .Y(_10209_));
 AO21x1_ASAP7_75t_SL _18402_ (.A1(_08958_),
    .A2(_10110_),
    .B(_10116_),
    .Y(_10210_));
 OAI21x1_ASAP7_75t_R _18404_ (.A1(_10209_),
    .A2(_10210_),
    .B(_08976_),
    .Y(_10212_));
 OAI21x1_ASAP7_75t_R _18405_ (.A1(_10208_),
    .A2(_10212_),
    .B(_08982_),
    .Y(_10213_));
 AOI21x1_ASAP7_75t_SL _18406_ (.A1(_08975_),
    .A2(_10205_),
    .B(_10213_),
    .Y(_10214_));
 AOI21x1_ASAP7_75t_SL _18407_ (.A1(_01041_),
    .A2(_08958_),
    .B(_10116_),
    .Y(_10215_));
 INVx1_ASAP7_75t_SL _18408_ (.A(_10215_),
    .Y(_10216_));
 NAND2x1_ASAP7_75t_L _18409_ (.A(_08958_),
    .B(_10103_),
    .Y(_10217_));
 OA21x2_ASAP7_75t_SL _18410_ (.A1(_08958_),
    .A2(_01041_),
    .B(_10116_),
    .Y(_10218_));
 NAND2x1_ASAP7_75t_R _18411_ (.A(_10217_),
    .B(_10218_),
    .Y(_10219_));
 AOI21x1_ASAP7_75t_R _18412_ (.A1(_10216_),
    .A2(_10219_),
    .B(_08975_),
    .Y(_10220_));
 AO21x1_ASAP7_75t_R _18414_ (.A1(_10144_),
    .A2(_10116_),
    .B(_08976_),
    .Y(_10222_));
 AO21x1_ASAP7_75t_SL _18415_ (.A1(_08958_),
    .A2(_10143_),
    .B(_10116_),
    .Y(_10223_));
 INVx1_ASAP7_75t_SL _18416_ (.A(_10133_),
    .Y(_10224_));
 NAND2x1_ASAP7_75t_R _18417_ (.A(_10116_),
    .B(_10224_),
    .Y(_10225_));
 OAI21x1_ASAP7_75t_SL _18418_ (.A1(_10223_),
    .A2(_10161_),
    .B(_10225_),
    .Y(_10226_));
 OAI21x1_ASAP7_75t_R _18421_ (.A1(_10222_),
    .A2(_10226_),
    .B(_10149_),
    .Y(_10229_));
 OAI21x1_ASAP7_75t_R _18422_ (.A1(_10220_),
    .A2(_10229_),
    .B(_08987_),
    .Y(_10230_));
 NOR2x1_ASAP7_75t_L _18423_ (.A(_10214_),
    .B(_10230_),
    .Y(_10231_));
 AND2x2_ASAP7_75t_SL _18424_ (.A(_08958_),
    .B(_08968_),
    .Y(_10232_));
 NAND2x1_ASAP7_75t_R _18425_ (.A(_10110_),
    .B(_10232_),
    .Y(_10233_));
 AOI21x1_ASAP7_75t_SL _18426_ (.A1(_08968_),
    .A2(_10177_),
    .B(_08976_),
    .Y(_10234_));
 NAND2x1_ASAP7_75t_SL _18427_ (.A(_10233_),
    .B(_10234_),
    .Y(_10235_));
 NOR2x1_ASAP7_75t_SL _18428_ (.A(_10104_),
    .B(_10103_),
    .Y(_10236_));
 OA21x2_ASAP7_75t_SL _18429_ (.A1(_10236_),
    .A2(_10113_),
    .B(_10116_),
    .Y(_10237_));
 NOR2x1_ASAP7_75t_R _18430_ (.A(_10235_),
    .B(_10237_),
    .Y(_10238_));
 NOR2x1_ASAP7_75t_SL _18431_ (.A(_08958_),
    .B(_10103_),
    .Y(_10239_));
 AO21x1_ASAP7_75t_SL _18432_ (.A1(_08958_),
    .A2(_10128_),
    .B(_08968_),
    .Y(_10240_));
 NOR2x1_ASAP7_75t_R _18433_ (.A(_10239_),
    .B(_10240_),
    .Y(_10241_));
 INVx1_ASAP7_75t_R _18434_ (.A(_01042_),
    .Y(_10242_));
 NOR2x2_ASAP7_75t_SL _18435_ (.A(_10242_),
    .B(_08958_),
    .Y(_10243_));
 AO21x1_ASAP7_75t_L _18436_ (.A1(_01043_),
    .A2(_08958_),
    .B(_10116_),
    .Y(_10244_));
 OAI21x1_ASAP7_75t_R _18437_ (.A1(_10243_),
    .A2(_10244_),
    .B(_08976_),
    .Y(_10245_));
 OAI21x1_ASAP7_75t_R _18438_ (.A1(_10241_),
    .A2(_10245_),
    .B(_10149_),
    .Y(_10246_));
 NOR2x1_ASAP7_75t_SL _18439_ (.A(_10238_),
    .B(_10246_),
    .Y(_10247_));
 AO21x1_ASAP7_75t_SL _18440_ (.A1(_08958_),
    .A2(_01042_),
    .B(_10116_),
    .Y(_10248_));
 NOR2x1_ASAP7_75t_L _18441_ (.A(_10161_),
    .B(_10248_),
    .Y(_10249_));
 NOR2x1_ASAP7_75t_SL _18442_ (.A(_10110_),
    .B(_08958_),
    .Y(_10250_));
 OAI21x1_ASAP7_75t_R _18443_ (.A1(_10250_),
    .A2(_10240_),
    .B(_08976_),
    .Y(_10251_));
 NOR2x1_ASAP7_75t_SL _18444_ (.A(_10249_),
    .B(_10251_),
    .Y(_10252_));
 AO21x1_ASAP7_75t_SL _18445_ (.A1(_08958_),
    .A2(_10128_),
    .B(_10116_),
    .Y(_10253_));
 NOR2x1_ASAP7_75t_R _18446_ (.A(_10192_),
    .B(_10253_),
    .Y(_10254_));
 NAND2x1_ASAP7_75t_SL _18447_ (.A(_08958_),
    .B(_01043_),
    .Y(_10255_));
 AO21x1_ASAP7_75t_R _18449_ (.A1(_10255_),
    .A2(_10116_),
    .B(_08976_),
    .Y(_10257_));
 OAI21x1_ASAP7_75t_R _18450_ (.A1(_10254_),
    .A2(_10257_),
    .B(_08982_),
    .Y(_10258_));
 OAI21x1_ASAP7_75t_R _18451_ (.A1(_10252_),
    .A2(_10258_),
    .B(_08988_),
    .Y(_10259_));
 INVx2_ASAP7_75t_SL _18452_ (.A(_08992_),
    .Y(_10260_));
 OAI21x1_ASAP7_75t_R _18453_ (.A1(_10247_),
    .A2(_10259_),
    .B(_10260_),
    .Y(_10261_));
 OAI22x1_ASAP7_75t_SL _18454_ (.A1(_10160_),
    .A2(_10200_),
    .B1(_10231_),
    .B2(_10261_),
    .Y(_00024_));
 NOR2x1_ASAP7_75t_SL _18455_ (.A(_01045_),
    .B(_08958_),
    .Y(_10262_));
 AOI21x1_ASAP7_75t_SL _18456_ (.A1(_10176_),
    .A2(_08958_),
    .B(_10116_),
    .Y(_10263_));
 NAND2x2_ASAP7_75t_SL _18457_ (.A(_10104_),
    .B(_10152_),
    .Y(_10264_));
 AOI22x1_ASAP7_75t_SL _18458_ (.A1(_10116_),
    .A2(_10262_),
    .B1(_10263_),
    .B2(_10264_),
    .Y(_10265_));
 AOI21x1_ASAP7_75t_R _18459_ (.A1(_08975_),
    .A2(_10265_),
    .B(_10149_),
    .Y(_10266_));
 INVx1_ASAP7_75t_SL _18460_ (.A(_10177_),
    .Y(_10267_));
 NAND2x1_ASAP7_75t_SL _18461_ (.A(_10104_),
    .B(_01046_),
    .Y(_10268_));
 INVx1_ASAP7_75t_SL _18462_ (.A(_10248_),
    .Y(_10269_));
 AOI21x1_ASAP7_75t_R _18463_ (.A1(_10268_),
    .A2(_10269_),
    .B(_08975_),
    .Y(_10270_));
 OAI21x1_ASAP7_75t_R _18464_ (.A1(_08968_),
    .A2(_10267_),
    .B(_10270_),
    .Y(_10271_));
 AND2x2_ASAP7_75t_R _18465_ (.A(_10266_),
    .B(_10271_),
    .Y(_10272_));
 OA21x2_ASAP7_75t_SL _18466_ (.A1(_10139_),
    .A2(_08968_),
    .B(_08976_),
    .Y(_10273_));
 AND2x2_ASAP7_75t_SL _18467_ (.A(_10144_),
    .B(_10116_),
    .Y(_10274_));
 INVx2_ASAP7_75t_SL _18468_ (.A(_10161_),
    .Y(_10275_));
 AOI21x1_ASAP7_75t_SL _18470_ (.A1(_10174_),
    .A2(_10275_),
    .B(_10116_),
    .Y(_10277_));
 NOR2x1_ASAP7_75t_L _18471_ (.A(_10274_),
    .B(_10277_),
    .Y(_10278_));
 AOI21x1_ASAP7_75t_R _18473_ (.A1(_10273_),
    .A2(_10278_),
    .B(_08982_),
    .Y(_10280_));
 AOI21x1_ASAP7_75t_SL _18474_ (.A1(_01043_),
    .A2(_10104_),
    .B(_08968_),
    .Y(_10281_));
 AOI21x1_ASAP7_75t_R _18475_ (.A1(_10153_),
    .A2(_10281_),
    .B(_08976_),
    .Y(_10282_));
 NAND2x1_ASAP7_75t_R _18476_ (.A(_10110_),
    .B(_10103_),
    .Y(_10283_));
 INVx1_ASAP7_75t_R _18477_ (.A(_10250_),
    .Y(_10284_));
 AO21x1_ASAP7_75t_R _18478_ (.A1(_10283_),
    .A2(_10284_),
    .B(_10116_),
    .Y(_10285_));
 NAND2x1_ASAP7_75t_R _18479_ (.A(_10282_),
    .B(_10285_),
    .Y(_10286_));
 AO21x1_ASAP7_75t_SL _18480_ (.A1(_10286_),
    .A2(_10280_),
    .B(_08987_),
    .Y(_10287_));
 AO21x1_ASAP7_75t_R _18481_ (.A1(_10104_),
    .A2(_01045_),
    .B(_08968_),
    .Y(_10288_));
 OAI22x1_ASAP7_75t_R _18482_ (.A1(_10288_),
    .A2(_10145_),
    .B1(_10161_),
    .B2(_10244_),
    .Y(_10289_));
 NAND2x1_ASAP7_75t_L _18483_ (.A(_10207_),
    .B(_10182_),
    .Y(_10290_));
 NAND2x2_ASAP7_75t_SL _18484_ (.A(_01044_),
    .B(_08958_),
    .Y(_10291_));
 OA21x2_ASAP7_75t_R _18486_ (.A1(_10291_),
    .A2(_10116_),
    .B(_08975_),
    .Y(_10293_));
 AOI21x1_ASAP7_75t_R _18487_ (.A1(_10290_),
    .A2(_10293_),
    .B(_10149_),
    .Y(_10294_));
 OAI21x1_ASAP7_75t_SL _18488_ (.A1(_08975_),
    .A2(_10289_),
    .B(_10294_),
    .Y(_10295_));
 AOI21x1_ASAP7_75t_R _18490_ (.A1(_01056_),
    .A2(_08968_),
    .B(_08975_),
    .Y(_10297_));
 NAND2x1_ASAP7_75t_SL _18491_ (.A(_01045_),
    .B(_08958_),
    .Y(_10298_));
 NAND2x1_ASAP7_75t_L _18492_ (.A(_10298_),
    .B(_10182_),
    .Y(_10299_));
 NAND2x1_ASAP7_75t_R _18493_ (.A(_10297_),
    .B(_10299_),
    .Y(_10300_));
 NAND2x1_ASAP7_75t_SL _18494_ (.A(_10298_),
    .B(_10140_),
    .Y(_10301_));
 INVx1_ASAP7_75t_R _18495_ (.A(_10243_),
    .Y(_10302_));
 AOI21x1_ASAP7_75t_SL _18496_ (.A1(_10302_),
    .A2(_10215_),
    .B(_08976_),
    .Y(_10303_));
 AOI21x1_ASAP7_75t_SL _18497_ (.A1(_10301_),
    .A2(_10303_),
    .B(_08982_),
    .Y(_10304_));
 AOI21x1_ASAP7_75t_R _18498_ (.A1(_10300_),
    .A2(_10304_),
    .B(_08988_),
    .Y(_10305_));
 AOI21x1_ASAP7_75t_R _18499_ (.A1(_10295_),
    .A2(_10305_),
    .B(_10260_),
    .Y(_10306_));
 OAI21x1_ASAP7_75t_SL _18500_ (.A1(_10272_),
    .A2(_10287_),
    .B(_10306_),
    .Y(_10307_));
 NAND2x1_ASAP7_75t_SL _18501_ (.A(_10143_),
    .B(_08958_),
    .Y(_10308_));
 NAND2x1_ASAP7_75t_SL _18502_ (.A(_10308_),
    .B(_10281_),
    .Y(_10309_));
 INVx1_ASAP7_75t_R _18503_ (.A(_10291_),
    .Y(_10310_));
 OAI21x1_ASAP7_75t_R _18504_ (.A1(_10177_),
    .A2(_10310_),
    .B(_08968_),
    .Y(_10311_));
 NAND3x1_ASAP7_75t_SL _18505_ (.A(_10309_),
    .B(_10311_),
    .C(_08982_),
    .Y(_10312_));
 NAND2x1_ASAP7_75t_L _18506_ (.A(_08958_),
    .B(_01046_),
    .Y(_10313_));
 NAND2x1_ASAP7_75t_SL _18507_ (.A(_10313_),
    .B(_10193_),
    .Y(_10314_));
 NAND2x1_ASAP7_75t_SL _18508_ (.A(_10217_),
    .B(_10206_),
    .Y(_10315_));
 NAND3x1_ASAP7_75t_R _18509_ (.A(_10314_),
    .B(_10315_),
    .C(_10149_),
    .Y(_10316_));
 NAND2x1_ASAP7_75t_SL _18510_ (.A(_10312_),
    .B(_10316_),
    .Y(_10317_));
 AND3x1_ASAP7_75t_R _18511_ (.A(_10149_),
    .B(_01058_),
    .C(_08968_),
    .Y(_10318_));
 OAI21x1_ASAP7_75t_SL _18512_ (.A1(_10177_),
    .A2(_10224_),
    .B(_10116_),
    .Y(_10319_));
 NAND2x1_ASAP7_75t_R _18513_ (.A(_08975_),
    .B(_10319_),
    .Y(_10320_));
 OAI21x1_ASAP7_75t_R _18514_ (.A1(_10318_),
    .A2(_10320_),
    .B(_08987_),
    .Y(_10321_));
 AOI21x1_ASAP7_75t_R _18515_ (.A1(_08976_),
    .A2(_10317_),
    .B(_10321_),
    .Y(_10322_));
 AOI21x1_ASAP7_75t_R _18517_ (.A1(_01050_),
    .A2(_08958_),
    .B(_08968_),
    .Y(_10324_));
 AOI22x1_ASAP7_75t_R _18518_ (.A1(_10324_),
    .A2(_10302_),
    .B1(_10263_),
    .B2(_10264_),
    .Y(_10325_));
 NAND2x1_ASAP7_75t_SL _18519_ (.A(_08976_),
    .B(_10325_),
    .Y(_10326_));
 NOR2x1p5_ASAP7_75t_L _18520_ (.A(_10145_),
    .B(_10162_),
    .Y(_10327_));
 OA21x2_ASAP7_75t_SL _18521_ (.A1(_10267_),
    .A2(_08968_),
    .B(_08975_),
    .Y(_10328_));
 AOI21x1_ASAP7_75t_SL _18522_ (.A1(_10328_),
    .A2(_10327_),
    .B(_08982_),
    .Y(_10329_));
 NAND2x1_ASAP7_75t_SL _18523_ (.A(_10326_),
    .B(_10329_),
    .Y(_10330_));
 OAI21x1_ASAP7_75t_R _18524_ (.A1(_10144_),
    .A2(_10154_),
    .B(_08968_),
    .Y(_10331_));
 OAI21x1_ASAP7_75t_R _18525_ (.A1(_10113_),
    .A2(_10145_),
    .B(_10116_),
    .Y(_10332_));
 AOI21x1_ASAP7_75t_R _18526_ (.A1(_10332_),
    .A2(_10331_),
    .B(_08975_),
    .Y(_10333_));
 NAND2x1_ASAP7_75t_SL _18527_ (.A(_10308_),
    .B(_10206_),
    .Y(_10334_));
 AOI21x1_ASAP7_75t_R _18528_ (.A1(_10334_),
    .A2(_10314_),
    .B(_08976_),
    .Y(_10335_));
 OAI21x1_ASAP7_75t_SL _18529_ (.A1(_10333_),
    .A2(_10335_),
    .B(_08982_),
    .Y(_10336_));
 AOI21x1_ASAP7_75t_SL _18530_ (.A1(_10336_),
    .A2(_10330_),
    .B(_08987_),
    .Y(_10337_));
 OAI21x1_ASAP7_75t_SL _18531_ (.A1(_10322_),
    .A2(_10337_),
    .B(_10260_),
    .Y(_10338_));
 NAND2x1_ASAP7_75t_SL _18532_ (.A(_10307_),
    .B(_10338_),
    .Y(_00025_));
 NOR2x1_ASAP7_75t_R _18533_ (.A(_10116_),
    .B(_10129_),
    .Y(_10339_));
 AOI21x1_ASAP7_75t_R _18534_ (.A1(_10174_),
    .A2(_10339_),
    .B(_08976_),
    .Y(_10340_));
 AOI21x1_ASAP7_75t_R _18535_ (.A1(_10183_),
    .A2(_10340_),
    .B(_08982_),
    .Y(_10341_));
 AO21x1_ASAP7_75t_R _18536_ (.A1(_10268_),
    .A2(_10291_),
    .B(_10116_),
    .Y(_10342_));
 AOI21x1_ASAP7_75t_R _18537_ (.A1(_10164_),
    .A2(_10167_),
    .B(_01042_),
    .Y(_10343_));
 OAI21x1_ASAP7_75t_R _18538_ (.A1(_10262_),
    .A2(_10343_),
    .B(_10116_),
    .Y(_10344_));
 AO21x1_ASAP7_75t_R _18539_ (.A1(_10342_),
    .A2(_10344_),
    .B(_08975_),
    .Y(_10345_));
 NAND2x1_ASAP7_75t_R _18540_ (.A(_10341_),
    .B(_10345_),
    .Y(_10346_));
 NAND2x1_ASAP7_75t_R _18541_ (.A(_10302_),
    .B(_10263_),
    .Y(_10347_));
 AO21x1_ASAP7_75t_R _18542_ (.A1(_10347_),
    .A2(_10240_),
    .B(_08976_),
    .Y(_10348_));
 AO21x1_ASAP7_75t_R _18543_ (.A1(_10167_),
    .A2(_10164_),
    .B(_01050_),
    .Y(_10349_));
 NOR2x2_ASAP7_75t_SL _18544_ (.A(_08958_),
    .B(_01043_),
    .Y(_10350_));
 INVx2_ASAP7_75t_L _18545_ (.A(_10350_),
    .Y(_10351_));
 NAND3x1_ASAP7_75t_R _18546_ (.A(_10349_),
    .B(_10351_),
    .C(_08968_),
    .Y(_10352_));
 NAND2x1_ASAP7_75t_SL _18547_ (.A(_10313_),
    .B(_10218_),
    .Y(_10353_));
 AND2x2_ASAP7_75t_SL _18548_ (.A(_10353_),
    .B(_08976_),
    .Y(_10354_));
 AOI21x1_ASAP7_75t_R _18549_ (.A1(_10352_),
    .A2(_10354_),
    .B(_10149_),
    .Y(_10355_));
 NAND2x1_ASAP7_75t_SL _18550_ (.A(_10348_),
    .B(_10355_),
    .Y(_10356_));
 AOI21x1_ASAP7_75t_SL _18551_ (.A1(_10346_),
    .A2(_10356_),
    .B(_08988_),
    .Y(_10357_));
 INVx1_ASAP7_75t_R _18552_ (.A(_10343_),
    .Y(_10358_));
 AOI21x1_ASAP7_75t_R _18553_ (.A1(_10358_),
    .A2(_10206_),
    .B(_08975_),
    .Y(_10359_));
 OR3x1_ASAP7_75t_R _18554_ (.A(_10236_),
    .B(_10116_),
    .C(_10170_),
    .Y(_10360_));
 NAND2x1_ASAP7_75t_R _18555_ (.A(_10359_),
    .B(_10360_),
    .Y(_10361_));
 INVx3_ASAP7_75t_SL _18556_ (.A(_10162_),
    .Y(_10362_));
 NAND2x1_ASAP7_75t_SL _18557_ (.A(_10120_),
    .B(_10281_),
    .Y(_10363_));
 OAI21x1_ASAP7_75t_SL _18558_ (.A1(_10154_),
    .A2(_10362_),
    .B(_10363_),
    .Y(_10364_));
 AOI21x1_ASAP7_75t_SL _18559_ (.A1(_08975_),
    .A2(_10364_),
    .B(_10149_),
    .Y(_10365_));
 NOR2x1_ASAP7_75t_R _18560_ (.A(_10350_),
    .B(_10169_),
    .Y(_10366_));
 AOI21x1_ASAP7_75t_R _18561_ (.A1(_10116_),
    .A2(_10343_),
    .B(_08975_),
    .Y(_10367_));
 OAI21x1_ASAP7_75t_R _18562_ (.A1(_10116_),
    .A2(_10366_),
    .B(_10367_),
    .Y(_10368_));
 AO21x1_ASAP7_75t_R _18563_ (.A1(_08958_),
    .A2(_01045_),
    .B(_10116_),
    .Y(_10369_));
 AOI21x1_ASAP7_75t_R _18564_ (.A1(_10116_),
    .A2(_10169_),
    .B(_08976_),
    .Y(_10370_));
 OAI21x1_ASAP7_75t_R _18565_ (.A1(_10239_),
    .A2(_10369_),
    .B(_10370_),
    .Y(_10371_));
 AO21x1_ASAP7_75t_R _18567_ (.A1(_10116_),
    .A2(_10170_),
    .B(_08982_),
    .Y(_10373_));
 AOI21x1_ASAP7_75t_R _18568_ (.A1(_10368_),
    .A2(_10371_),
    .B(_10373_),
    .Y(_10374_));
 AOI21x1_ASAP7_75t_SL _18569_ (.A1(_10365_),
    .A2(_10361_),
    .B(_10374_),
    .Y(_10375_));
 OAI21x1_ASAP7_75t_SL _18570_ (.A1(_10375_),
    .A2(_08987_),
    .B(_10260_),
    .Y(_10376_));
 NAND2x1_ASAP7_75t_SL _18571_ (.A(_10351_),
    .B(_10263_),
    .Y(_10377_));
 NAND3x1_ASAP7_75t_SL _18572_ (.A(_10319_),
    .B(_10377_),
    .C(_08976_),
    .Y(_10378_));
 NAND2x1p5_ASAP7_75t_SL _18573_ (.A(_10162_),
    .B(_10298_),
    .Y(_10379_));
 INVx1_ASAP7_75t_R _18574_ (.A(_10222_),
    .Y(_10380_));
 AOI21x1_ASAP7_75t_SL _18575_ (.A1(_10380_),
    .A2(_10379_),
    .B(_10149_),
    .Y(_10381_));
 NAND2x1_ASAP7_75t_SL _18576_ (.A(_10381_),
    .B(_10378_),
    .Y(_10382_));
 INVx1_ASAP7_75t_R _18577_ (.A(_01052_),
    .Y(_10383_));
 OA21x2_ASAP7_75t_R _18578_ (.A1(_10383_),
    .A2(_10116_),
    .B(_08975_),
    .Y(_10384_));
 AOI21x1_ASAP7_75t_R _18579_ (.A1(_10240_),
    .A2(_10384_),
    .B(_08982_),
    .Y(_10385_));
 OA21x2_ASAP7_75t_R _18580_ (.A1(_01057_),
    .A2(_08968_),
    .B(_08976_),
    .Y(_10386_));
 NAND2x1_ASAP7_75t_SL _18581_ (.A(_10386_),
    .B(_10342_),
    .Y(_10387_));
 AOI21x1_ASAP7_75t_R _18582_ (.A1(_10385_),
    .A2(_10387_),
    .B(_08988_),
    .Y(_10388_));
 AOI21x1_ASAP7_75t_SL _18583_ (.A1(_10388_),
    .A2(_10382_),
    .B(_10260_),
    .Y(_10389_));
 INVx1_ASAP7_75t_R _18584_ (.A(_01058_),
    .Y(_10390_));
 AOI21x1_ASAP7_75t_R _18585_ (.A1(_10104_),
    .A2(_10103_),
    .B(_10116_),
    .Y(_10391_));
 AOI21x1_ASAP7_75t_R _18586_ (.A1(_10207_),
    .A2(_10391_),
    .B(_08976_),
    .Y(_10392_));
 OA21x2_ASAP7_75t_R _18587_ (.A1(_10390_),
    .A2(_08968_),
    .B(_10392_),
    .Y(_10393_));
 AND3x1_ASAP7_75t_R _18588_ (.A(_10268_),
    .B(_10116_),
    .C(_10308_),
    .Y(_10394_));
 OAI21x1_ASAP7_75t_SL _18589_ (.A1(_10153_),
    .A2(_10116_),
    .B(_08976_),
    .Y(_10395_));
 AO21x1_ASAP7_75t_SL _18590_ (.A1(_08968_),
    .A2(_10203_),
    .B(_10395_),
    .Y(_10396_));
 OAI21x1_ASAP7_75t_R _18591_ (.A1(_10394_),
    .A2(_10396_),
    .B(_10149_),
    .Y(_10397_));
 AOI21x1_ASAP7_75t_R _18592_ (.A1(_10313_),
    .A2(_10187_),
    .B(_08975_),
    .Y(_10398_));
 NAND2x1_ASAP7_75t_R _18593_ (.A(_10183_),
    .B(_10398_),
    .Y(_10399_));
 NAND2x1_ASAP7_75t_SL _18594_ (.A(_01041_),
    .B(_08958_),
    .Y(_10400_));
 INVx2_ASAP7_75t_SL _18595_ (.A(_10400_),
    .Y(_10401_));
 NOR2x1_ASAP7_75t_R _18596_ (.A(_10401_),
    .B(_10123_),
    .Y(_10402_));
 NAND2x1_ASAP7_75t_R _18597_ (.A(_10155_),
    .B(_10116_),
    .Y(_10403_));
 NAND2x1_ASAP7_75t_R _18598_ (.A(_08975_),
    .B(_10403_),
    .Y(_10404_));
 OA21x2_ASAP7_75t_SL _18599_ (.A1(_10402_),
    .A2(_10404_),
    .B(_08982_),
    .Y(_10405_));
 AOI21x1_ASAP7_75t_SL _18600_ (.A1(_10399_),
    .A2(_10405_),
    .B(_08987_),
    .Y(_10406_));
 OAI21x1_ASAP7_75t_SL _18601_ (.A1(_10393_),
    .A2(_10397_),
    .B(_10406_),
    .Y(_10407_));
 NAND2x1_ASAP7_75t_SL _18602_ (.A(_10407_),
    .B(_10389_),
    .Y(_10408_));
 OAI21x1_ASAP7_75t_SL _18603_ (.A1(_10357_),
    .A2(_10376_),
    .B(_10408_),
    .Y(_00026_));
 OAI21x1_ASAP7_75t_R _18604_ (.A1(_10144_),
    .A2(_10401_),
    .B(_08968_),
    .Y(_10409_));
 OAI21x1_ASAP7_75t_R _18605_ (.A1(_10203_),
    .A2(_10145_),
    .B(_10116_),
    .Y(_10410_));
 AOI21x1_ASAP7_75t_R _18606_ (.A1(_10409_),
    .A2(_10410_),
    .B(_08975_),
    .Y(_10411_));
 NOR2x1_ASAP7_75t_R _18607_ (.A(_01042_),
    .B(_08958_),
    .Y(_10412_));
 OAI21x1_ASAP7_75t_R _18608_ (.A1(_10412_),
    .A2(_10169_),
    .B(_08968_),
    .Y(_10413_));
 AOI21x1_ASAP7_75t_R _18609_ (.A1(_10413_),
    .A2(_10353_),
    .B(_08976_),
    .Y(_10414_));
 OAI21x1_ASAP7_75t_R _18610_ (.A1(_10411_),
    .A2(_10414_),
    .B(_08982_),
    .Y(_10415_));
 NOR2x1_ASAP7_75t_SL _18611_ (.A(_08975_),
    .B(_10215_),
    .Y(_10416_));
 NAND2x1_ASAP7_75t_SL _18612_ (.A(_10313_),
    .B(_10281_),
    .Y(_10417_));
 AOI21x1_ASAP7_75t_R _18613_ (.A1(_10416_),
    .A2(_10417_),
    .B(_08982_),
    .Y(_10418_));
 NAND2x1_ASAP7_75t_R _18614_ (.A(_01043_),
    .B(_10103_),
    .Y(_10419_));
 AOI21x1_ASAP7_75t_R _18615_ (.A1(_10419_),
    .A2(_10206_),
    .B(_08976_),
    .Y(_10420_));
 OAI21x1_ASAP7_75t_SL _18616_ (.A1(_10236_),
    .A2(_10362_),
    .B(_10420_),
    .Y(_10421_));
 NAND2x1_ASAP7_75t_L _18617_ (.A(_10421_),
    .B(_10418_),
    .Y(_10422_));
 NAND3x1_ASAP7_75t_SL _18618_ (.A(_10422_),
    .B(_10415_),
    .C(_08987_),
    .Y(_10423_));
 AOI21x1_ASAP7_75t_SL _18619_ (.A1(_10253_),
    .A2(_10420_),
    .B(_08982_),
    .Y(_10424_));
 NAND2x1_ASAP7_75t_SL _18620_ (.A(_10120_),
    .B(_10218_),
    .Y(_10425_));
 NAND2x1_ASAP7_75t_SL _18621_ (.A(_10425_),
    .B(_10270_),
    .Y(_10426_));
 AOI21x1_ASAP7_75t_R _18622_ (.A1(_10424_),
    .A2(_10426_),
    .B(_08987_),
    .Y(_10427_));
 OAI21x1_ASAP7_75t_R _18623_ (.A1(_10203_),
    .A2(_10310_),
    .B(_08968_),
    .Y(_10428_));
 AO21x1_ASAP7_75t_R _18624_ (.A1(_10267_),
    .A2(_10153_),
    .B(_08968_),
    .Y(_10429_));
 AOI21x1_ASAP7_75t_R _18625_ (.A1(_10428_),
    .A2(_10429_),
    .B(_08976_),
    .Y(_10430_));
 AOI21x1_ASAP7_75t_R _18626_ (.A1(_10202_),
    .A2(_10133_),
    .B(_10212_),
    .Y(_10431_));
 OAI21x1_ASAP7_75t_SL _18627_ (.A1(_10430_),
    .A2(_10431_),
    .B(_08982_),
    .Y(_10432_));
 AOI21x1_ASAP7_75t_R _18628_ (.A1(_10427_),
    .A2(_10432_),
    .B(_10260_),
    .Y(_10433_));
 NAND2x1_ASAP7_75t_L _18629_ (.A(_10423_),
    .B(_10433_),
    .Y(_10434_));
 NAND2x1p5_ASAP7_75t_L _18630_ (.A(_10116_),
    .B(_10161_),
    .Y(_10435_));
 AOI21x1_ASAP7_75t_SL _18631_ (.A1(_08968_),
    .A2(_10113_),
    .B(_08975_),
    .Y(_10436_));
 OAI21x1_ASAP7_75t_R _18632_ (.A1(_10149_),
    .A2(_10435_),
    .B(_10436_),
    .Y(_10437_));
 NAND2x1_ASAP7_75t_L _18633_ (.A(_08968_),
    .B(_10401_),
    .Y(_10438_));
 OAI21x1_ASAP7_75t_R _18634_ (.A1(_10224_),
    .A2(_10239_),
    .B(_10116_),
    .Y(_10439_));
 AOI21x1_ASAP7_75t_R _18635_ (.A1(_10438_),
    .A2(_10439_),
    .B(_08982_),
    .Y(_10440_));
 OAI21x1_ASAP7_75t_SL _18636_ (.A1(_10437_),
    .A2(_10440_),
    .B(_08987_),
    .Y(_10441_));
 INVx1_ASAP7_75t_R _18637_ (.A(_10170_),
    .Y(_10442_));
 OA21x2_ASAP7_75t_SL _18638_ (.A1(_10442_),
    .A2(_10116_),
    .B(_08982_),
    .Y(_10443_));
 NAND2x1_ASAP7_75t_SL _18639_ (.A(_10363_),
    .B(_10443_),
    .Y(_10444_));
 AOI21x1_ASAP7_75t_SL _18640_ (.A1(_10202_),
    .A2(_10255_),
    .B(_08982_),
    .Y(_10445_));
 OAI21x1_ASAP7_75t_SL _18641_ (.A1(_10350_),
    .A2(_10248_),
    .B(_10445_),
    .Y(_10446_));
 AOI21x1_ASAP7_75t_SL _18642_ (.A1(_10444_),
    .A2(_10446_),
    .B(_08976_),
    .Y(_10447_));
 NOR2x1_ASAP7_75t_SL _18643_ (.A(_10441_),
    .B(_10447_),
    .Y(_10448_));
 NOR2x1_ASAP7_75t_R _18644_ (.A(_01048_),
    .B(_10104_),
    .Y(_10449_));
 OAI21x1_ASAP7_75t_R _18645_ (.A1(_10250_),
    .A2(_10449_),
    .B(_08968_),
    .Y(_10450_));
 AOI21x1_ASAP7_75t_R _18646_ (.A1(_10319_),
    .A2(_10450_),
    .B(_08976_),
    .Y(_10451_));
 OAI21x1_ASAP7_75t_R _18647_ (.A1(_10359_),
    .A2(_10451_),
    .B(_10149_),
    .Y(_10452_));
 AOI21x1_ASAP7_75t_R _18648_ (.A1(_10147_),
    .A2(_10290_),
    .B(_08976_),
    .Y(_10453_));
 INVx1_ASAP7_75t_SL _18649_ (.A(_10255_),
    .Y(_10454_));
 OAI21x1_ASAP7_75t_SL _18650_ (.A1(_10170_),
    .A2(_10454_),
    .B(_08968_),
    .Y(_10455_));
 NAND2x1_ASAP7_75t_SL _18651_ (.A(_01042_),
    .B(_08958_),
    .Y(_10456_));
 NAND2x1p5_ASAP7_75t_SL _18652_ (.A(_10202_),
    .B(_10456_),
    .Y(_10457_));
 AOI21x1_ASAP7_75t_SL _18653_ (.A1(_10455_),
    .A2(_10457_),
    .B(_08975_),
    .Y(_10458_));
 OAI21x1_ASAP7_75t_SL _18654_ (.A1(_10458_),
    .A2(_10453_),
    .B(_08982_),
    .Y(_10459_));
 AOI21x1_ASAP7_75t_SL _18655_ (.A1(_10459_),
    .A2(_10452_),
    .B(_08987_),
    .Y(_10460_));
 OAI21x1_ASAP7_75t_SL _18656_ (.A1(_10460_),
    .A2(_10448_),
    .B(_10260_),
    .Y(_10461_));
 NAND2x1_ASAP7_75t_SL _18657_ (.A(_10434_),
    .B(_10461_),
    .Y(_00027_));
 NOR2x1p5_ASAP7_75t_SL _18658_ (.A(_10288_),
    .B(_10154_),
    .Y(_10462_));
 NOR2x1_ASAP7_75t_SL _18659_ (.A(_10235_),
    .B(_10462_),
    .Y(_10463_));
 AO21x1_ASAP7_75t_R _18660_ (.A1(_10201_),
    .A2(_08968_),
    .B(_08975_),
    .Y(_10464_));
 OAI21x1_ASAP7_75t_R _18661_ (.A1(_10324_),
    .A2(_10464_),
    .B(_08982_),
    .Y(_10465_));
 OA21x2_ASAP7_75t_SL _18662_ (.A1(_10463_),
    .A2(_10465_),
    .B(_08988_),
    .Y(_10466_));
 INVx1_ASAP7_75t_SL _18663_ (.A(_10314_),
    .Y(_10467_));
 OR3x1_ASAP7_75t_L _18664_ (.A(_10103_),
    .B(_10104_),
    .C(_08968_),
    .Y(_10468_));
 NOR2x1_ASAP7_75t_R _18665_ (.A(_08975_),
    .B(_10274_),
    .Y(_10469_));
 NAND2x1_ASAP7_75t_R _18666_ (.A(_10468_),
    .B(_10469_),
    .Y(_10470_));
 AND2x2_ASAP7_75t_SL _18667_ (.A(_10206_),
    .B(_10456_),
    .Y(_10471_));
 AO21x1_ASAP7_75t_R _18668_ (.A1(_08958_),
    .A2(_08968_),
    .B(_08976_),
    .Y(_10472_));
 OA21x2_ASAP7_75t_SL _18669_ (.A1(_10471_),
    .A2(_10472_),
    .B(_10149_),
    .Y(_10473_));
 OAI21x1_ASAP7_75t_R _18670_ (.A1(_10467_),
    .A2(_10470_),
    .B(_10473_),
    .Y(_10474_));
 NAND2x1p5_ASAP7_75t_SL _18671_ (.A(_10474_),
    .B(_10466_),
    .Y(_10475_));
 NAND2x1_ASAP7_75t_R _18672_ (.A(_10176_),
    .B(_10116_),
    .Y(_10476_));
 OAI21x1_ASAP7_75t_R _18673_ (.A1(_10153_),
    .A2(_10116_),
    .B(_10476_),
    .Y(_10477_));
 AOI21x1_ASAP7_75t_SL _18674_ (.A1(_08975_),
    .A2(_10477_),
    .B(_10149_),
    .Y(_10478_));
 AND2x4_ASAP7_75t_L _18675_ (.A(_10120_),
    .B(_08968_),
    .Y(_10479_));
 NAND2x1_ASAP7_75t_SL _18676_ (.A(_10268_),
    .B(_10479_),
    .Y(_10480_));
 NOR2x1_ASAP7_75t_R _18677_ (.A(_08975_),
    .B(_10131_),
    .Y(_10481_));
 NAND2x1_ASAP7_75t_L _18678_ (.A(_10480_),
    .B(_10481_),
    .Y(_10482_));
 AOI21x1_ASAP7_75t_SL _18679_ (.A1(_10478_),
    .A2(_10482_),
    .B(_08988_),
    .Y(_10483_));
 NAND3x1_ASAP7_75t_R _18680_ (.A(_10419_),
    .B(_08968_),
    .C(_10139_),
    .Y(_10484_));
 AOI21x1_ASAP7_75t_SL _18681_ (.A1(_10197_),
    .A2(_10484_),
    .B(_08976_),
    .Y(_10485_));
 AO21x1_ASAP7_75t_R _18682_ (.A1(_10283_),
    .A2(_10268_),
    .B(_08968_),
    .Y(_10486_));
 AOI21x1_ASAP7_75t_R _18683_ (.A1(_10450_),
    .A2(_10486_),
    .B(_08975_),
    .Y(_10487_));
 OAI21x1_ASAP7_75t_R _18684_ (.A1(_10485_),
    .A2(_10487_),
    .B(_10149_),
    .Y(_10488_));
 AOI21x1_ASAP7_75t_R _18685_ (.A1(_10483_),
    .A2(_10488_),
    .B(_08992_),
    .Y(_10489_));
 NAND2x1_ASAP7_75t_SL _18686_ (.A(_10475_),
    .B(_10489_),
    .Y(_10490_));
 INVx2_ASAP7_75t_SL _18687_ (.A(_10395_),
    .Y(_10491_));
 NOR2x1_ASAP7_75t_R _18688_ (.A(_10170_),
    .B(_10175_),
    .Y(_10492_));
 AOI21x1_ASAP7_75t_SL _18689_ (.A1(_10491_),
    .A2(_10492_),
    .B(_10149_),
    .Y(_10493_));
 NOR2x1_ASAP7_75t_L _18690_ (.A(_08968_),
    .B(_10243_),
    .Y(_10494_));
 AO21x1_ASAP7_75t_L _18691_ (.A1(_10400_),
    .A2(_10494_),
    .B(_10126_),
    .Y(_10495_));
 NAND2x1_ASAP7_75t_L _18692_ (.A(_10493_),
    .B(_10495_),
    .Y(_10496_));
 NOR2x1_ASAP7_75t_R _18693_ (.A(_10104_),
    .B(_01046_),
    .Y(_10497_));
 OAI21x1_ASAP7_75t_R _18694_ (.A1(_10129_),
    .A2(_10497_),
    .B(_08968_),
    .Y(_10498_));
 AOI21x1_ASAP7_75t_R _18695_ (.A1(_10344_),
    .A2(_10498_),
    .B(_08975_),
    .Y(_10499_));
 OAI21x1_ASAP7_75t_R _18696_ (.A1(_10144_),
    .A2(_10497_),
    .B(_08968_),
    .Y(_10500_));
 AOI21x1_ASAP7_75t_R _18697_ (.A1(_10500_),
    .A2(_10301_),
    .B(_08976_),
    .Y(_10501_));
 OAI21x1_ASAP7_75t_R _18698_ (.A1(_10499_),
    .A2(_10501_),
    .B(_10149_),
    .Y(_10502_));
 AOI21x1_ASAP7_75t_SL _18699_ (.A1(_10496_),
    .A2(_10502_),
    .B(_08988_),
    .Y(_10503_));
 NAND2x1_ASAP7_75t_R _18700_ (.A(_10207_),
    .B(_10391_),
    .Y(_10504_));
 AOI21x1_ASAP7_75t_R _18701_ (.A1(_10315_),
    .A2(_10504_),
    .B(_08976_),
    .Y(_10505_));
 NOR2x1_ASAP7_75t_L _18702_ (.A(_08958_),
    .B(_01046_),
    .Y(_10506_));
 OAI21x1_ASAP7_75t_R _18703_ (.A1(_10196_),
    .A2(_10506_),
    .B(_08968_),
    .Y(_10507_));
 OAI21x1_ASAP7_75t_R _18704_ (.A1(_10209_),
    .A2(_10236_),
    .B(_10116_),
    .Y(_10508_));
 AOI21x1_ASAP7_75t_SL _18705_ (.A1(_10507_),
    .A2(_10508_),
    .B(_08975_),
    .Y(_10509_));
 OAI21x1_ASAP7_75t_R _18706_ (.A1(_10505_),
    .A2(_10509_),
    .B(_10149_),
    .Y(_10510_));
 OA21x2_ASAP7_75t_R _18707_ (.A1(_10479_),
    .A2(_10113_),
    .B(_08976_),
    .Y(_10511_));
 NAND2x1_ASAP7_75t_R _18708_ (.A(_10217_),
    .B(_10187_),
    .Y(_10512_));
 AOI21x1_ASAP7_75t_SL _18709_ (.A1(_10309_),
    .A2(_10512_),
    .B(_08976_),
    .Y(_10513_));
 OAI21x1_ASAP7_75t_R _18710_ (.A1(_10511_),
    .A2(_10513_),
    .B(_08982_),
    .Y(_10514_));
 AOI21x1_ASAP7_75t_R _18711_ (.A1(_10510_),
    .A2(_10514_),
    .B(_08987_),
    .Y(_10515_));
 OAI21x1_ASAP7_75t_SL _18712_ (.A1(_10503_),
    .A2(_10515_),
    .B(_08992_),
    .Y(_10516_));
 NAND2x1_ASAP7_75t_SL _18713_ (.A(_10516_),
    .B(_10490_),
    .Y(_00028_));
 NAND2x1_ASAP7_75t_R _18714_ (.A(_08968_),
    .B(_10103_),
    .Y(_10517_));
 AOI21x1_ASAP7_75t_R _18715_ (.A1(_10517_),
    .A2(_10508_),
    .B(_08976_),
    .Y(_10518_));
 AO21x1_ASAP7_75t_R _18716_ (.A1(_10267_),
    .A2(_10133_),
    .B(_10116_),
    .Y(_10519_));
 AO21x1_ASAP7_75t_R _18717_ (.A1(_10283_),
    .A2(_10255_),
    .B(_08968_),
    .Y(_10520_));
 AOI21x1_ASAP7_75t_R _18718_ (.A1(_10519_),
    .A2(_10520_),
    .B(_08975_),
    .Y(_10521_));
 OAI21x1_ASAP7_75t_R _18719_ (.A1(_10518_),
    .A2(_10521_),
    .B(_08982_),
    .Y(_10522_));
 INVx1_ASAP7_75t_R _18720_ (.A(_10506_),
    .Y(_10523_));
 AO21x1_ASAP7_75t_L _18721_ (.A1(_10523_),
    .A2(_10324_),
    .B(_10395_),
    .Y(_10524_));
 OA21x2_ASAP7_75t_R _18722_ (.A1(_10358_),
    .A2(_08968_),
    .B(_08975_),
    .Y(_10525_));
 AO21x1_ASAP7_75t_SL _18723_ (.A1(_10152_),
    .A2(_10104_),
    .B(_10223_),
    .Y(_10526_));
 AOI21x1_ASAP7_75t_R _18724_ (.A1(_10525_),
    .A2(_10526_),
    .B(_08982_),
    .Y(_10527_));
 AOI21x1_ASAP7_75t_SL _18725_ (.A1(_10524_),
    .A2(_10527_),
    .B(_08988_),
    .Y(_10528_));
 NAND2x1_ASAP7_75t_L _18726_ (.A(_10522_),
    .B(_10528_),
    .Y(_10529_));
 NAND3x1_ASAP7_75t_R _18727_ (.A(_10288_),
    .B(_08976_),
    .C(_10291_),
    .Y(_10530_));
 NOR2x1p5_ASAP7_75t_SL _18728_ (.A(_08976_),
    .B(_10202_),
    .Y(_10531_));
 AOI21x1_ASAP7_75t_SL _18729_ (.A1(_10455_),
    .A2(_10531_),
    .B(_08982_),
    .Y(_10532_));
 AOI21x1_ASAP7_75t_SL _18730_ (.A1(_10530_),
    .A2(_10532_),
    .B(_08987_),
    .Y(_10533_));
 AO21x1_ASAP7_75t_R _18731_ (.A1(_10193_),
    .A2(_10456_),
    .B(_08976_),
    .Y(_10534_));
 AO21x1_ASAP7_75t_SL _18732_ (.A1(_10284_),
    .A2(_10174_),
    .B(_10116_),
    .Y(_10535_));
 AOI21x1_ASAP7_75t_SL _18733_ (.A1(_10120_),
    .A2(_10140_),
    .B(_08975_),
    .Y(_10536_));
 AOI21x1_ASAP7_75t_R _18734_ (.A1(_10535_),
    .A2(_10536_),
    .B(_10149_),
    .Y(_10537_));
 OAI21x1_ASAP7_75t_R _18735_ (.A1(_10237_),
    .A2(_10534_),
    .B(_10537_),
    .Y(_10538_));
 AOI21x1_ASAP7_75t_SL _18736_ (.A1(_10538_),
    .A2(_10533_),
    .B(_10260_),
    .Y(_10539_));
 NAND2x1_ASAP7_75t_SL _18737_ (.A(_10539_),
    .B(_10529_),
    .Y(_10540_));
 NOR2x1p5_ASAP7_75t_SL _18738_ (.A(_10186_),
    .B(_10362_),
    .Y(_10541_));
 NAND2x1_ASAP7_75t_R _18739_ (.A(_10435_),
    .B(_10367_),
    .Y(_10542_));
 OAI22x1_ASAP7_75t_R _18740_ (.A1(_10476_),
    .A2(_08958_),
    .B1(_01047_),
    .B2(_10116_),
    .Y(_10543_));
 AOI21x1_ASAP7_75t_R _18741_ (.A1(_08975_),
    .A2(_10543_),
    .B(_08982_),
    .Y(_10544_));
 OAI21x1_ASAP7_75t_SL _18742_ (.A1(_10542_),
    .A2(_10541_),
    .B(_10544_),
    .Y(_10545_));
 OR3x1_ASAP7_75t_L _18743_ (.A(_10269_),
    .B(_08975_),
    .C(_10175_),
    .Y(_10546_));
 OA21x2_ASAP7_75t_R _18744_ (.A1(_10350_),
    .A2(_10116_),
    .B(_10291_),
    .Y(_10547_));
 AOI21x1_ASAP7_75t_R _18745_ (.A1(_10547_),
    .A2(_10328_),
    .B(_10149_),
    .Y(_10548_));
 AOI21x1_ASAP7_75t_R _18746_ (.A1(_10546_),
    .A2(_10548_),
    .B(_08988_),
    .Y(_10549_));
 AOI21x1_ASAP7_75t_SL _18747_ (.A1(_10549_),
    .A2(_10545_),
    .B(_08992_),
    .Y(_10550_));
 OR3x1_ASAP7_75t_L _18748_ (.A(_10239_),
    .B(_08968_),
    .C(_10121_),
    .Y(_10551_));
 OA21x2_ASAP7_75t_SL _18749_ (.A1(_10161_),
    .A2(_10253_),
    .B(_08976_),
    .Y(_10552_));
 AO21x1_ASAP7_75t_R _18750_ (.A1(_10110_),
    .A2(_08968_),
    .B(_08976_),
    .Y(_10553_));
 OAI21x1_ASAP7_75t_R _18751_ (.A1(_10553_),
    .A2(_10208_),
    .B(_08982_),
    .Y(_10554_));
 AO21x1_ASAP7_75t_SL _18752_ (.A1(_10551_),
    .A2(_10552_),
    .B(_10554_),
    .Y(_10555_));
 AOI22x1_ASAP7_75t_R _18753_ (.A1(_10116_),
    .A2(_10177_),
    .B1(_10232_),
    .B2(_01047_),
    .Y(_10556_));
 AOI21x1_ASAP7_75t_R _18754_ (.A1(_10367_),
    .A2(_10556_),
    .B(_08982_),
    .Y(_10557_));
 NAND2x1_ASAP7_75t_R _18755_ (.A(_10174_),
    .B(_10351_),
    .Y(_10558_));
 AO21x1_ASAP7_75t_SL _18756_ (.A1(_10116_),
    .A2(_10558_),
    .B(_10235_),
    .Y(_10559_));
 AOI21x1_ASAP7_75t_R _18757_ (.A1(_10557_),
    .A2(_10559_),
    .B(_08987_),
    .Y(_10560_));
 NAND2x1_ASAP7_75t_SL _18758_ (.A(_10555_),
    .B(_10560_),
    .Y(_10561_));
 NAND2x1_ASAP7_75t_SL _18759_ (.A(_10561_),
    .B(_10550_),
    .Y(_10562_));
 NAND2x1_ASAP7_75t_SL _18760_ (.A(_10562_),
    .B(_10540_),
    .Y(_00029_));
 OA21x2_ASAP7_75t_R _18761_ (.A1(_10103_),
    .A2(_08968_),
    .B(_08975_),
    .Y(_10563_));
 AO21x1_ASAP7_75t_SL _18762_ (.A1(_10283_),
    .A2(_10268_),
    .B(_10116_),
    .Y(_10564_));
 NAND2x1_ASAP7_75t_R _18763_ (.A(_10563_),
    .B(_10564_),
    .Y(_10565_));
 AO21x1_ASAP7_75t_SL _18764_ (.A1(_10349_),
    .A2(_10442_),
    .B(_10116_),
    .Y(_10566_));
 AOI21x1_ASAP7_75t_R _18765_ (.A1(_10469_),
    .A2(_10566_),
    .B(_08987_),
    .Y(_10567_));
 NAND2x1_ASAP7_75t_R _18766_ (.A(_10565_),
    .B(_10567_),
    .Y(_10568_));
 AOI21x1_ASAP7_75t_SL _18767_ (.A1(_10264_),
    .A2(_10324_),
    .B(_08976_),
    .Y(_10569_));
 OAI21x1_ASAP7_75t_R _18768_ (.A1(_10239_),
    .A2(_10253_),
    .B(_10569_),
    .Y(_10570_));
 OA21x2_ASAP7_75t_R _18769_ (.A1(_10383_),
    .A2(_10116_),
    .B(_08976_),
    .Y(_10571_));
 AO21x1_ASAP7_75t_SL _18770_ (.A1(_10291_),
    .A2(_10264_),
    .B(_08968_),
    .Y(_10572_));
 AOI21x1_ASAP7_75t_SL _18771_ (.A1(_10572_),
    .A2(_10571_),
    .B(_08988_),
    .Y(_10573_));
 AOI21x1_ASAP7_75t_SL _18772_ (.A1(_10573_),
    .A2(_10570_),
    .B(_10149_),
    .Y(_10574_));
 AOI21x1_ASAP7_75t_SL _18773_ (.A1(_10574_),
    .A2(_10568_),
    .B(_10260_),
    .Y(_10575_));
 AO21x1_ASAP7_75t_R _18774_ (.A1(_10113_),
    .A2(_08968_),
    .B(_08976_),
    .Y(_10576_));
 AOI221x1_ASAP7_75t_R _18775_ (.A1(_01040_),
    .A2(_10232_),
    .B1(_10120_),
    .B2(_10494_),
    .C(_10576_),
    .Y(_10577_));
 AND2x2_ASAP7_75t_SL _18776_ (.A(_10455_),
    .B(_08976_),
    .Y(_10578_));
 NAND2x1_ASAP7_75t_L _18777_ (.A(_10153_),
    .B(_10206_),
    .Y(_10579_));
 AO21x1_ASAP7_75t_SL _18778_ (.A1(_10579_),
    .A2(_10578_),
    .B(_08987_),
    .Y(_10580_));
 AOI21x1_ASAP7_75t_SL _18779_ (.A1(_10206_),
    .A2(_10153_),
    .B(_08976_),
    .Y(_10581_));
 OAI21x1_ASAP7_75t_SL _18780_ (.A1(_10145_),
    .A2(_10123_),
    .B(_10581_),
    .Y(_10582_));
 NOR2x1_ASAP7_75t_SL _18781_ (.A(_10123_),
    .B(_10497_),
    .Y(_10583_));
 OA21x2_ASAP7_75t_SL _18782_ (.A1(_10583_),
    .A2(_10134_),
    .B(_08987_),
    .Y(_10584_));
 AOI21x1_ASAP7_75t_SL _18783_ (.A1(_10584_),
    .A2(_10582_),
    .B(_08982_),
    .Y(_10585_));
 OAI21x1_ASAP7_75t_R _18784_ (.A1(_10577_),
    .A2(_10580_),
    .B(_10585_),
    .Y(_10586_));
 NAND2x1_ASAP7_75t_SL _18785_ (.A(_10575_),
    .B(_10586_),
    .Y(_10587_));
 OAI21x1_ASAP7_75t_R _18786_ (.A1(_10250_),
    .A2(_10240_),
    .B(_10297_),
    .Y(_10588_));
 OA21x2_ASAP7_75t_SL _18787_ (.A1(_08968_),
    .A2(_10264_),
    .B(_08975_),
    .Y(_10589_));
 AOI21x1_ASAP7_75t_SL _18788_ (.A1(_10455_),
    .A2(_10589_),
    .B(_08982_),
    .Y(_10590_));
 AOI21x1_ASAP7_75t_SL _18789_ (.A1(_10590_),
    .A2(_10588_),
    .B(_08987_),
    .Y(_10591_));
 AO21x1_ASAP7_75t_R _18790_ (.A1(_10207_),
    .A2(_10139_),
    .B(_10116_),
    .Y(_10592_));
 AO21x1_ASAP7_75t_R _18791_ (.A1(_10268_),
    .A2(_10291_),
    .B(_08968_),
    .Y(_10593_));
 AOI21x1_ASAP7_75t_R _18792_ (.A1(_10592_),
    .A2(_10593_),
    .B(_08976_),
    .Y(_10594_));
 INVx1_ASAP7_75t_R _18793_ (.A(_10494_),
    .Y(_10595_));
 AO21x1_ASAP7_75t_SL _18794_ (.A1(_10419_),
    .A2(_10351_),
    .B(_10116_),
    .Y(_10596_));
 INVx1_ASAP7_75t_R _18795_ (.A(_10273_),
    .Y(_10597_));
 AOI21x1_ASAP7_75t_SL _18796_ (.A1(_10595_),
    .A2(_10596_),
    .B(_10597_),
    .Y(_10598_));
 OAI21x1_ASAP7_75t_R _18797_ (.A1(_10594_),
    .A2(_10598_),
    .B(_08982_),
    .Y(_10599_));
 NAND2x1_ASAP7_75t_SL _18798_ (.A(_10599_),
    .B(_10591_),
    .Y(_10600_));
 AO21x1_ASAP7_75t_R _18799_ (.A1(_01046_),
    .A2(_10104_),
    .B(_08968_),
    .Y(_10601_));
 OA21x2_ASAP7_75t_R _18800_ (.A1(_01053_),
    .A2(_10116_),
    .B(_08975_),
    .Y(_10602_));
 OAI21x1_ASAP7_75t_R _18801_ (.A1(_10121_),
    .A2(_10601_),
    .B(_10602_),
    .Y(_10603_));
 NAND2x1p5_ASAP7_75t_L _18802_ (.A(_10264_),
    .B(_10269_),
    .Y(_10604_));
 AOI21x1_ASAP7_75t_R _18803_ (.A1(_10273_),
    .A2(_10604_),
    .B(_10149_),
    .Y(_10605_));
 AOI21x1_ASAP7_75t_R _18804_ (.A1(_10603_),
    .A2(_10605_),
    .B(_08988_),
    .Y(_10606_));
 AO21x1_ASAP7_75t_R _18805_ (.A1(_08958_),
    .A2(_10185_),
    .B(_08968_),
    .Y(_10607_));
 AOI21x1_ASAP7_75t_SL _18806_ (.A1(_10480_),
    .A2(_10607_),
    .B(_08975_),
    .Y(_10608_));
 OAI21x1_ASAP7_75t_R _18807_ (.A1(_10340_),
    .A2(_10608_),
    .B(_10149_),
    .Y(_10609_));
 AOI21x1_ASAP7_75t_SL _18808_ (.A1(_10609_),
    .A2(_10606_),
    .B(_08992_),
    .Y(_10610_));
 NAND2x1_ASAP7_75t_SL _18809_ (.A(_10600_),
    .B(_10610_),
    .Y(_10611_));
 NAND2x1_ASAP7_75t_SL _18810_ (.A(_10587_),
    .B(_10611_),
    .Y(_00030_));
 AOI221x1_ASAP7_75t_R _18811_ (.A1(_10120_),
    .A2(_10494_),
    .B1(_10313_),
    .B2(_10187_),
    .C(_08982_),
    .Y(_10612_));
 NOR2x1_ASAP7_75t_L _18812_ (.A(_10149_),
    .B(_10494_),
    .Y(_10613_));
 AO21x1_ASAP7_75t_R _18813_ (.A1(_10480_),
    .A2(_10613_),
    .B(_08976_),
    .Y(_10614_));
 OAI21x1_ASAP7_75t_R _18814_ (.A1(_10129_),
    .A2(_10145_),
    .B(_10116_),
    .Y(_10615_));
 NAND2x1_ASAP7_75t_R _18815_ (.A(_10143_),
    .B(_10104_),
    .Y(_10616_));
 AOI21x1_ASAP7_75t_SL _18816_ (.A1(_10616_),
    .A2(_10263_),
    .B(_10149_),
    .Y(_10617_));
 AOI21x1_ASAP7_75t_R _18817_ (.A1(_10615_),
    .A2(_10617_),
    .B(_08975_),
    .Y(_10618_));
 OAI21x1_ASAP7_75t_SL _18818_ (.A1(_10216_),
    .A2(_10243_),
    .B(_10445_),
    .Y(_10619_));
 AOI21x1_ASAP7_75t_SL _18819_ (.A1(_10619_),
    .A2(_10618_),
    .B(_08987_),
    .Y(_10620_));
 OAI21x1_ASAP7_75t_SL _18820_ (.A1(_10612_),
    .A2(_10614_),
    .B(_10620_),
    .Y(_10621_));
 NAND2x1_ASAP7_75t_R _18821_ (.A(_10435_),
    .B(_10234_),
    .Y(_10622_));
 AND2x2_ASAP7_75t_L _18822_ (.A(_10123_),
    .B(_08976_),
    .Y(_10623_));
 NAND2x1_ASAP7_75t_R _18823_ (.A(_10201_),
    .B(_10218_),
    .Y(_10624_));
 AOI21x1_ASAP7_75t_SL _18824_ (.A1(_10623_),
    .A2(_10624_),
    .B(_08982_),
    .Y(_10625_));
 AOI21x1_ASAP7_75t_R _18825_ (.A1(_10622_),
    .A2(_10625_),
    .B(_08988_),
    .Y(_10626_));
 INVx1_ASAP7_75t_R _18826_ (.A(_10201_),
    .Y(_10627_));
 OAI21x1_ASAP7_75t_R _18827_ (.A1(_10627_),
    .A2(_10601_),
    .B(_10392_),
    .Y(_10628_));
 NAND2x1_ASAP7_75t_R _18828_ (.A(_01043_),
    .B(_10116_),
    .Y(_10629_));
 OAI21x1_ASAP7_75t_R _18829_ (.A1(_10497_),
    .A2(_10188_),
    .B(_10629_),
    .Y(_10630_));
 AOI21x1_ASAP7_75t_R _18830_ (.A1(_08976_),
    .A2(_10630_),
    .B(_10149_),
    .Y(_10631_));
 NAND2x1_ASAP7_75t_SL _18831_ (.A(_10628_),
    .B(_10631_),
    .Y(_10632_));
 AOI21x1_ASAP7_75t_SL _18832_ (.A1(_10626_),
    .A2(_10632_),
    .B(_08992_),
    .Y(_10633_));
 NAND2x1_ASAP7_75t_SL _18833_ (.A(_10633_),
    .B(_10621_),
    .Y(_10634_));
 AND3x1_ASAP7_75t_R _18834_ (.A(_01046_),
    .B(_08958_),
    .C(_08968_),
    .Y(_10635_));
 NOR2x1_ASAP7_75t_R _18835_ (.A(_08968_),
    .B(_10349_),
    .Y(_10636_));
 OR3x1_ASAP7_75t_R _18836_ (.A(_10636_),
    .B(_08982_),
    .C(_10144_),
    .Y(_10637_));
 AO21x1_ASAP7_75t_SL _18837_ (.A1(_10275_),
    .A2(_10133_),
    .B(_10116_),
    .Y(_10638_));
 AND2x2_ASAP7_75t_R _18838_ (.A(_10201_),
    .B(_10116_),
    .Y(_10639_));
 AOI21x1_ASAP7_75t_SL _18839_ (.A1(_10616_),
    .A2(_10639_),
    .B(_10149_),
    .Y(_10640_));
 AOI21x1_ASAP7_75t_R _18840_ (.A1(_10638_),
    .A2(_10640_),
    .B(_08976_),
    .Y(_10641_));
 OAI21x1_ASAP7_75t_SL _18841_ (.A1(_10635_),
    .A2(_10637_),
    .B(_10641_),
    .Y(_10642_));
 OA21x2_ASAP7_75t_R _18842_ (.A1(_01045_),
    .A2(_08968_),
    .B(_10149_),
    .Y(_10643_));
 NAND2x1_ASAP7_75t_R _18843_ (.A(_10643_),
    .B(_10564_),
    .Y(_10644_));
 NAND2x1_ASAP7_75t_R _18844_ (.A(_10201_),
    .B(_10182_),
    .Y(_10645_));
 AOI21x1_ASAP7_75t_R _18845_ (.A1(_10351_),
    .A2(_10479_),
    .B(_10149_),
    .Y(_10646_));
 AOI21x1_ASAP7_75t_R _18846_ (.A1(_10645_),
    .A2(_10646_),
    .B(_08975_),
    .Y(_10647_));
 AOI21x1_ASAP7_75t_R _18847_ (.A1(_10644_),
    .A2(_10647_),
    .B(_08987_),
    .Y(_10648_));
 NAND2x1_ASAP7_75t_L _18848_ (.A(_10642_),
    .B(_10648_),
    .Y(_10649_));
 NAND2x1_ASAP7_75t_R _18849_ (.A(_10468_),
    .B(_10481_),
    .Y(_10650_));
 AO21x1_ASAP7_75t_R _18850_ (.A1(_01040_),
    .A2(_08968_),
    .B(_08976_),
    .Y(_10651_));
 OA21x2_ASAP7_75t_R _18851_ (.A1(_10651_),
    .A2(_10636_),
    .B(_08982_),
    .Y(_10652_));
 OAI21x1_ASAP7_75t_R _18852_ (.A1(_10467_),
    .A2(_10650_),
    .B(_10652_),
    .Y(_10653_));
 OA21x2_ASAP7_75t_R _18853_ (.A1(_01059_),
    .A2(_10116_),
    .B(_08975_),
    .Y(_10654_));
 AO21x1_ASAP7_75t_R _18854_ (.A1(_10442_),
    .A2(_10400_),
    .B(_08968_),
    .Y(_10655_));
 AOI21x1_ASAP7_75t_R _18855_ (.A1(_10654_),
    .A2(_10655_),
    .B(_08982_),
    .Y(_10656_));
 NAND2x1_ASAP7_75t_SL _18856_ (.A(_10264_),
    .B(_10215_),
    .Y(_10657_));
 NAND3x1_ASAP7_75t_SL _18857_ (.A(_10273_),
    .B(_10657_),
    .C(_10403_),
    .Y(_10658_));
 AOI21x1_ASAP7_75t_R _18858_ (.A1(_10656_),
    .A2(_10658_),
    .B(_08988_),
    .Y(_10659_));
 AOI21x1_ASAP7_75t_R _18859_ (.A1(_10653_),
    .A2(_10659_),
    .B(_10260_),
    .Y(_10660_));
 NAND2x1_ASAP7_75t_SL _18860_ (.A(_10649_),
    .B(_10660_),
    .Y(_10661_));
 NAND2x1_ASAP7_75t_SL _18861_ (.A(_10661_),
    .B(_10634_),
    .Y(_00031_));
 NOR2x1_ASAP7_75t_R _18865_ (.A(_00444_),
    .B(_00574_),
    .Y(_10665_));
 XNOR2x2_ASAP7_75t_SL _18866_ (.A(_00575_),
    .B(_00582_),
    .Y(_10666_));
 XOR2x2_ASAP7_75t_SL _18867_ (.A(_00640_),
    .B(_00608_),
    .Y(_10667_));
 XOR2x2_ASAP7_75t_SL _18868_ (.A(_10667_),
    .B(_10666_),
    .Y(_10668_));
 XOR2x2_ASAP7_75t_SL _18869_ (.A(_00614_),
    .B(_00607_),
    .Y(_10669_));
 XOR2x2_ASAP7_75t_SL _18870_ (.A(_00672_),
    .B(_10669_),
    .Y(_10670_));
 INVx1_ASAP7_75t_R _18871_ (.A(_10670_),
    .Y(_10671_));
 NAND2x1_ASAP7_75t_L _18872_ (.A(_10668_),
    .B(_10671_),
    .Y(_10672_));
 INVx2_ASAP7_75t_SL _18873_ (.A(_10668_),
    .Y(_10673_));
 NAND2x1p5_ASAP7_75t_L _18874_ (.A(_10670_),
    .B(_10673_),
    .Y(_10674_));
 INVx3_ASAP7_75t_SL _18875_ (.A(_00574_),
    .Y(_10675_));
 AOI21x1_ASAP7_75t_SL _18878_ (.A1(_10674_),
    .A2(_10672_),
    .B(_10675_),
    .Y(_10678_));
 OAI21x1_ASAP7_75t_SL _18879_ (.A1(_10678_),
    .A2(_10665_),
    .B(_00855_),
    .Y(_10679_));
 AND2x2_ASAP7_75t_R _18881_ (.A(_10675_),
    .B(_00444_),
    .Y(_10681_));
 XOR2x1_ASAP7_75t_SL _18883_ (.A(_10670_),
    .Y(_10683_),
    .B(_10668_));
 NOR2x1_ASAP7_75t_SL _18884_ (.A(_10675_),
    .B(_10683_),
    .Y(_10684_));
 INVx1_ASAP7_75t_R _18885_ (.A(_00855_),
    .Y(_10685_));
 OAI21x1_ASAP7_75t_SL _18886_ (.A1(_10684_),
    .A2(_10681_),
    .B(_10685_),
    .Y(_10686_));
 NAND2x2_ASAP7_75t_SL _18887_ (.A(_10686_),
    .B(_10679_),
    .Y(_10687_));
 INVx1_ASAP7_75t_R _18892_ (.A(_00671_),
    .Y(_10691_));
 XOR2x2_ASAP7_75t_L _18893_ (.A(_00582_),
    .B(_00614_),
    .Y(_10692_));
 NAND2x1_ASAP7_75t_SL _18894_ (.A(_10691_),
    .B(_10692_),
    .Y(_10693_));
 XNOR2x2_ASAP7_75t_SL _18895_ (.A(_00582_),
    .B(_00614_),
    .Y(_10694_));
 NAND2x1_ASAP7_75t_SL _18896_ (.A(_00671_),
    .B(_10694_),
    .Y(_10695_));
 XOR2x2_ASAP7_75t_SL _18897_ (.A(_00607_),
    .B(_00639_),
    .Y(_10696_));
 INVx1_ASAP7_75t_SL _18898_ (.A(_10696_),
    .Y(_10697_));
 AOI21x1_ASAP7_75t_SL _18899_ (.A1(_10695_),
    .A2(_10693_),
    .B(_10697_),
    .Y(_10698_));
 NAND2x1_ASAP7_75t_SL _18900_ (.A(_00671_),
    .B(_10692_),
    .Y(_10699_));
 NAND2x1_ASAP7_75t_SL _18901_ (.A(_10691_),
    .B(_10694_),
    .Y(_10700_));
 AOI21x1_ASAP7_75t_SL _18902_ (.A1(_10700_),
    .A2(_10699_),
    .B(_10696_),
    .Y(_10701_));
 NOR2x1_ASAP7_75t_SL _18903_ (.A(_10698_),
    .B(_10701_),
    .Y(_10702_));
 AND2x2_ASAP7_75t_SL _18904_ (.A(_10675_),
    .B(_00445_),
    .Y(_10703_));
 AOI21x1_ASAP7_75t_SL _18905_ (.A1(_00574_),
    .A2(_10702_),
    .B(_10703_),
    .Y(_10704_));
 XNOR2x2_ASAP7_75t_SL _18906_ (.A(_00854_),
    .B(_10704_),
    .Y(_01067_));
 INVx1_ASAP7_75t_R _18907_ (.A(_00609_),
    .Y(_10705_));
 XOR2x2_ASAP7_75t_SL _18908_ (.A(_00576_),
    .B(_00608_),
    .Y(_10706_));
 NAND2x1_ASAP7_75t_L _18909_ (.A(_10705_),
    .B(_10706_),
    .Y(_10707_));
 XNOR2x2_ASAP7_75t_SL _18910_ (.A(_00576_),
    .B(_00608_),
    .Y(_10708_));
 NAND2x1_ASAP7_75t_R _18911_ (.A(_00609_),
    .B(_10708_),
    .Y(_10709_));
 XNOR2x2_ASAP7_75t_SL _18912_ (.A(_00641_),
    .B(_00673_),
    .Y(_10710_));
 AOI21x1_ASAP7_75t_SL _18913_ (.A1(_10707_),
    .A2(_10709_),
    .B(_10710_),
    .Y(_10711_));
 NAND2x1_ASAP7_75t_L _18914_ (.A(_00609_),
    .B(_10706_),
    .Y(_10712_));
 NAND2x1_ASAP7_75t_SL _18915_ (.A(_10705_),
    .B(_10708_),
    .Y(_10713_));
 XOR2x1_ASAP7_75t_SL _18916_ (.A(_00641_),
    .Y(_10714_),
    .B(_00673_));
 AOI21x1_ASAP7_75t_SL _18917_ (.A1(_10712_),
    .A2(_10713_),
    .B(_10714_),
    .Y(_10715_));
 OAI21x1_ASAP7_75t_SL _18918_ (.A1(_10711_),
    .A2(_10715_),
    .B(_00574_),
    .Y(_10716_));
 OR2x2_ASAP7_75t_SL _18919_ (.A(_00574_),
    .B(_00446_),
    .Y(_10717_));
 NAND3x1_ASAP7_75t_SL _18920_ (.A(_10716_),
    .B(_00856_),
    .C(_10717_),
    .Y(_10718_));
 AOI21x1_ASAP7_75t_SL _18921_ (.A1(_10717_),
    .A2(_10716_),
    .B(_00856_),
    .Y(_10719_));
 INVx2_ASAP7_75t_SL _18922_ (.A(_10719_),
    .Y(_10720_));
 NAND2x2_ASAP7_75t_SL _18923_ (.A(_10718_),
    .B(_10720_),
    .Y(_10721_));
 XOR2x2_ASAP7_75t_SL _18926_ (.A(_00854_),
    .B(_10704_),
    .Y(_10723_));
 INVx1_ASAP7_75t_R _18928_ (.A(_00856_),
    .Y(_10724_));
 NAND3x1_ASAP7_75t_SL _18929_ (.A(_10716_),
    .B(_10724_),
    .C(_10717_),
    .Y(_10725_));
 AOI21x1_ASAP7_75t_SL _18930_ (.A1(_10717_),
    .A2(_10716_),
    .B(_10724_),
    .Y(_10726_));
 INVx2_ASAP7_75t_SL _18931_ (.A(_10726_),
    .Y(_10727_));
 NAND2x2_ASAP7_75t_SL _18932_ (.A(_10725_),
    .B(_10727_),
    .Y(_10728_));
 XOR2x2_ASAP7_75t_SL _18935_ (.A(_00613_),
    .B(_00645_),
    .Y(_10730_));
 XOR2x2_ASAP7_75t_R _18936_ (.A(_10730_),
    .B(_00677_),
    .Y(_10731_));
 XOR2x2_ASAP7_75t_R _18937_ (.A(_00580_),
    .B(_00612_),
    .Y(_10732_));
 INVx1_ASAP7_75t_SL _18938_ (.A(_10732_),
    .Y(_10733_));
 XOR2x2_ASAP7_75t_SL _18939_ (.A(_10731_),
    .B(_10733_),
    .Y(_10734_));
 NOR2x1_ASAP7_75t_SL _18945_ (.A(_00574_),
    .B(_00550_),
    .Y(_10740_));
 AO21x1_ASAP7_75t_SL _18946_ (.A1(_10734_),
    .A2(_00574_),
    .B(_10740_),
    .Y(_10741_));
 XOR2x2_ASAP7_75t_SL _18947_ (.A(_10741_),
    .B(_00861_),
    .Y(_10742_));
 XNOR2x2_ASAP7_75t_SL _18950_ (.A(_00643_),
    .B(_00675_),
    .Y(_10745_));
 XOR2x2_ASAP7_75t_SL _18951_ (.A(_00610_),
    .B(_00614_),
    .Y(_10746_));
 XOR2x2_ASAP7_75t_R _18952_ (.A(_10745_),
    .B(_10746_),
    .Y(_10747_));
 XOR2x2_ASAP7_75t_L _18953_ (.A(_00578_),
    .B(_00582_),
    .Y(_10748_));
 XOR2x2_ASAP7_75t_R _18954_ (.A(_10748_),
    .B(_00611_),
    .Y(_10749_));
 XOR2x2_ASAP7_75t_SL _18955_ (.A(_10747_),
    .B(_10749_),
    .Y(_10750_));
 NOR2x1_ASAP7_75t_R _18958_ (.A(_00574_),
    .B(_00552_),
    .Y(_10753_));
 AOI21x1_ASAP7_75t_SL _18959_ (.A1(_00574_),
    .A2(_10750_),
    .B(_10753_),
    .Y(_10754_));
 XNOR2x2_ASAP7_75t_SL _18960_ (.A(_00858_),
    .B(_10754_),
    .Y(_10755_));
 AO21x1_ASAP7_75t_R _18963_ (.A1(_10720_),
    .A2(_10718_),
    .B(_01063_),
    .Y(_10758_));
 XOR2x2_ASAP7_75t_SL _18966_ (.A(_00577_),
    .B(_00582_),
    .Y(_10761_));
 XNOR2x2_ASAP7_75t_L _18967_ (.A(_00610_),
    .B(_10761_),
    .Y(_10762_));
 XNOR2x2_ASAP7_75t_R _18968_ (.A(_00642_),
    .B(_00674_),
    .Y(_10763_));
 XOR2x2_ASAP7_75t_SL _18969_ (.A(_00609_),
    .B(_00614_),
    .Y(_10764_));
 XOR2x2_ASAP7_75t_SL _18970_ (.A(_10763_),
    .B(_10764_),
    .Y(_10765_));
 XNOR2x2_ASAP7_75t_SL _18971_ (.A(_10762_),
    .B(_10765_),
    .Y(_10766_));
 NOR2x1_ASAP7_75t_R _18973_ (.A(_00574_),
    .B(_00553_),
    .Y(_10768_));
 AOI21x1_ASAP7_75t_SL _18974_ (.A1(_00574_),
    .A2(_10766_),
    .B(_10768_),
    .Y(_10769_));
 XOR2x2_ASAP7_75t_SL _18975_ (.A(_10769_),
    .B(_00857_),
    .Y(_10770_));
 AOI21x1_ASAP7_75t_SL _18977_ (.A1(_10728_),
    .A2(_10687_),
    .B(_10770_),
    .Y(_10772_));
 NAND2x1_ASAP7_75t_SL _18978_ (.A(_10758_),
    .B(_10772_),
    .Y(_10773_));
 NOR2x2_ASAP7_75t_SL _18979_ (.A(_10721_),
    .B(_10723_),
    .Y(_10774_));
 INVx1_ASAP7_75t_SL _18980_ (.A(_10774_),
    .Y(_10775_));
 INVx1_ASAP7_75t_SL _18981_ (.A(_01068_),
    .Y(_10776_));
 AO21x1_ASAP7_75t_SL _18982_ (.A1(_10720_),
    .A2(_10718_),
    .B(_10776_),
    .Y(_10777_));
 XNOR2x2_ASAP7_75t_SL _18983_ (.A(_00857_),
    .B(_10769_),
    .Y(_10778_));
 AO21x1_ASAP7_75t_SL _18986_ (.A1(_10775_),
    .A2(_10777_),
    .B(_10778_),
    .Y(_10781_));
 NAND2x1_ASAP7_75t_SL _18987_ (.A(_10773_),
    .B(_10781_),
    .Y(_10782_));
 INVx2_ASAP7_75t_SL _18988_ (.A(_01066_),
    .Y(_10783_));
 NOR2x1_ASAP7_75t_SL _18989_ (.A(_10783_),
    .B(_10721_),
    .Y(_10784_));
 NOR2x1_ASAP7_75t_SL _18990_ (.A(_10778_),
    .B(_10784_),
    .Y(_10785_));
 INVx1_ASAP7_75t_L _18991_ (.A(_10785_),
    .Y(_10786_));
 NAND2x1_ASAP7_75t_R _18994_ (.A(_00446_),
    .B(_10675_),
    .Y(_10789_));
 NOR2x1_ASAP7_75t_R _18995_ (.A(_10711_),
    .B(_10715_),
    .Y(_10790_));
 NAND2x1_ASAP7_75t_L _18996_ (.A(_00574_),
    .B(_10790_),
    .Y(_10791_));
 AOI21x1_ASAP7_75t_R _18997_ (.A1(_10789_),
    .A2(_10791_),
    .B(_00856_),
    .Y(_10792_));
 INVx2_ASAP7_75t_SL _18998_ (.A(_01064_),
    .Y(_10793_));
 OAI21x1_ASAP7_75t_SL _18999_ (.A1(_10726_),
    .A2(_10792_),
    .B(_10793_),
    .Y(_10794_));
 AOI21x1_ASAP7_75t_R _19000_ (.A1(_10789_),
    .A2(_10791_),
    .B(_10724_),
    .Y(_10795_));
 OAI21x1_ASAP7_75t_SL _19001_ (.A1(_10719_),
    .A2(_10795_),
    .B(_01062_),
    .Y(_10796_));
 AO21x1_ASAP7_75t_SL _19003_ (.A1(_10794_),
    .A2(_10796_),
    .B(_10770_),
    .Y(_10798_));
 AOI21x1_ASAP7_75t_R _19005_ (.A1(_10786_),
    .A2(_10798_),
    .B(_10755_),
    .Y(_10800_));
 AOI21x1_ASAP7_75t_R _19006_ (.A1(_10755_),
    .A2(_10782_),
    .B(_10800_),
    .Y(_10801_));
 NOR2x1_ASAP7_75t_R _19007_ (.A(_10742_),
    .B(_10801_),
    .Y(_10802_));
 NAND2x1_ASAP7_75t_SL _19008_ (.A(_10723_),
    .B(_10687_),
    .Y(_10803_));
 INVx1_ASAP7_75t_R _19009_ (.A(_10803_),
    .Y(_10804_));
 NAND2x1_ASAP7_75t_SL _19010_ (.A(_10728_),
    .B(_10804_),
    .Y(_10805_));
 AOI21x1_ASAP7_75t_SL _19011_ (.A1(_10718_),
    .A2(_10720_),
    .B(_01068_),
    .Y(_10806_));
 NOR2x1_ASAP7_75t_SL _19012_ (.A(_10806_),
    .B(_10770_),
    .Y(_10807_));
 INVx2_ASAP7_75t_SL _19015_ (.A(_10755_),
    .Y(_10810_));
 OAI21x1_ASAP7_75t_R _19017_ (.A1(_10778_),
    .A2(_10794_),
    .B(_10810_),
    .Y(_10812_));
 AO21x1_ASAP7_75t_R _19018_ (.A1(_10805_),
    .A2(_10807_),
    .B(_10812_),
    .Y(_10813_));
 OAI21x1_ASAP7_75t_SL _19020_ (.A1(_10770_),
    .A2(_10794_),
    .B(_10755_),
    .Y(_10815_));
 INVx1_ASAP7_75t_R _19021_ (.A(_10815_),
    .Y(_10816_));
 INVx1_ASAP7_75t_SL _19022_ (.A(_01069_),
    .Y(_10817_));
 AOI21x1_ASAP7_75t_SL _19023_ (.A1(_10718_),
    .A2(_10720_),
    .B(_10817_),
    .Y(_10818_));
 NOR2x1_ASAP7_75t_R _19024_ (.A(_10818_),
    .B(_10778_),
    .Y(_10819_));
 OAI21x1_ASAP7_75t_SL _19025_ (.A1(_10721_),
    .A2(_10803_),
    .B(_10819_),
    .Y(_10820_));
 INVx1_ASAP7_75t_SL _19026_ (.A(_10742_),
    .Y(_10821_));
 AOI21x1_ASAP7_75t_R _19027_ (.A1(_10816_),
    .A2(_10820_),
    .B(_10821_),
    .Y(_10822_));
 NOR2x1_ASAP7_75t_R _19028_ (.A(_00574_),
    .B(_00551_),
    .Y(_10823_));
 INVx1_ASAP7_75t_R _19029_ (.A(_10823_),
    .Y(_10824_));
 XOR2x2_ASAP7_75t_SL _19031_ (.A(_00612_),
    .B(_00644_),
    .Y(_10826_));
 XOR2x2_ASAP7_75t_L _19032_ (.A(_10826_),
    .B(_00676_),
    .Y(_10827_));
 XNOR2x2_ASAP7_75t_R _19033_ (.A(_00579_),
    .B(_00611_),
    .Y(_10828_));
 XOR2x2_ASAP7_75t_R _19034_ (.A(_10827_),
    .B(_10828_),
    .Y(_10829_));
 NAND2x1_ASAP7_75t_R _19035_ (.A(_00574_),
    .B(_10829_),
    .Y(_10830_));
 INVx1_ASAP7_75t_R _19036_ (.A(_00859_),
    .Y(_10831_));
 AOI21x1_ASAP7_75t_R _19037_ (.A1(_10824_),
    .A2(_10830_),
    .B(_10831_),
    .Y(_10832_));
 AO21x1_ASAP7_75t_R _19038_ (.A1(_10829_),
    .A2(_00574_),
    .B(_10823_),
    .Y(_10833_));
 NOR2x1_ASAP7_75t_SL _19039_ (.A(_00859_),
    .B(_10833_),
    .Y(_10834_));
 NOR2x1_ASAP7_75t_SL _19040_ (.A(_10832_),
    .B(_10834_),
    .Y(_10835_));
 AO21x1_ASAP7_75t_R _19042_ (.A1(_10813_),
    .A2(_10822_),
    .B(_10835_),
    .Y(_10837_));
 OAI21x1_ASAP7_75t_SL _19043_ (.A1(_10719_),
    .A2(_10795_),
    .B(_10783_),
    .Y(_10838_));
 OAI21x1_ASAP7_75t_R _19044_ (.A1(_10770_),
    .A2(_10838_),
    .B(_10755_),
    .Y(_10839_));
 INVx1_ASAP7_75t_SL _19045_ (.A(_10839_),
    .Y(_10840_));
 NAND2x2_ASAP7_75t_SL _19046_ (.A(_10721_),
    .B(_01067_),
    .Y(_10841_));
 INVx1_ASAP7_75t_SL _19047_ (.A(_10841_),
    .Y(_10842_));
 AOI21x1_ASAP7_75t_SL _19048_ (.A1(_01067_),
    .A2(_10687_),
    .B(_10721_),
    .Y(_10843_));
 OAI21x1_ASAP7_75t_SL _19050_ (.A1(_10842_),
    .A2(_10843_),
    .B(_10770_),
    .Y(_10845_));
 NAND2x1_ASAP7_75t_R _19051_ (.A(_10840_),
    .B(_10845_),
    .Y(_10846_));
 OA21x2_ASAP7_75t_SL _19053_ (.A1(_10770_),
    .A2(_10838_),
    .B(_10810_),
    .Y(_10848_));
 INVx1_ASAP7_75t_SL _19054_ (.A(_01063_),
    .Y(_10849_));
 AOI21x1_ASAP7_75t_SL _19055_ (.A1(_10725_),
    .A2(_10727_),
    .B(_10849_),
    .Y(_10850_));
 NOR2x2_ASAP7_75t_SL _19056_ (.A(_10778_),
    .B(_10850_),
    .Y(_10851_));
 AO21x1_ASAP7_75t_R _19057_ (.A1(_10727_),
    .A2(_10725_),
    .B(_01069_),
    .Y(_10852_));
 NOR2x1_ASAP7_75t_SL _19059_ (.A(_10770_),
    .B(_10852_),
    .Y(_10854_));
 NOR2x1p5_ASAP7_75t_SL _19060_ (.A(_10854_),
    .B(_10851_),
    .Y(_10855_));
 AOI21x1_ASAP7_75t_SL _19061_ (.A1(_10855_),
    .A2(_10848_),
    .B(_10742_),
    .Y(_10856_));
 NAND2x1_ASAP7_75t_SL _19062_ (.A(_10846_),
    .B(_10856_),
    .Y(_10857_));
 OR2x2_ASAP7_75t_R _19064_ (.A(_10778_),
    .B(_01076_),
    .Y(_10859_));
 NOR2x1_ASAP7_75t_SL _19065_ (.A(_01063_),
    .B(_10728_),
    .Y(_10860_));
 AOI21x1_ASAP7_75t_SL _19066_ (.A1(_10778_),
    .A2(_10860_),
    .B(_10755_),
    .Y(_10861_));
 AOI21x1_ASAP7_75t_R _19067_ (.A1(_10859_),
    .A2(_10861_),
    .B(_10821_),
    .Y(_10862_));
 INVx2_ASAP7_75t_R _19068_ (.A(_10838_),
    .Y(_10863_));
 AOI21x1_ASAP7_75t_SL _19069_ (.A1(_10723_),
    .A2(_10687_),
    .B(_10721_),
    .Y(_10864_));
 OAI21x1_ASAP7_75t_SL _19071_ (.A1(_10863_),
    .A2(_10864_),
    .B(_10778_),
    .Y(_10866_));
 INVx1_ASAP7_75t_R _19073_ (.A(_01062_),
    .Y(_10868_));
 AO21x1_ASAP7_75t_L _19074_ (.A1(_10727_),
    .A2(_10725_),
    .B(_10868_),
    .Y(_10869_));
 NAND2x1_ASAP7_75t_SL _19075_ (.A(_10869_),
    .B(_10841_),
    .Y(_10870_));
 OAI21x1_ASAP7_75t_SL _19076_ (.A1(_10719_),
    .A2(_10795_),
    .B(_10793_),
    .Y(_10871_));
 OAI21x1_ASAP7_75t_SL _19077_ (.A1(_10770_),
    .A2(_10871_),
    .B(_10755_),
    .Y(_10872_));
 AOI21x1_ASAP7_75t_R _19078_ (.A1(_10770_),
    .A2(_10870_),
    .B(_10872_),
    .Y(_10873_));
 NAND2x1_ASAP7_75t_SL _19079_ (.A(_10866_),
    .B(_10873_),
    .Y(_10874_));
 INVx2_ASAP7_75t_SL _19080_ (.A(_10835_),
    .Y(_10875_));
 AOI21x1_ASAP7_75t_L _19082_ (.A1(_10862_),
    .A2(_10874_),
    .B(_10875_),
    .Y(_10877_));
 XNOR2x2_ASAP7_75t_R _19083_ (.A(_00581_),
    .B(_00613_),
    .Y(_10878_));
 INVx2_ASAP7_75t_R _19084_ (.A(_00678_),
    .Y(_10879_));
 XOR2x2_ASAP7_75t_R _19085_ (.A(_10878_),
    .B(_10879_),
    .Y(_10880_));
 XNOR2x2_ASAP7_75t_R _19086_ (.A(_00614_),
    .B(_00646_),
    .Y(_10881_));
 XOR2x2_ASAP7_75t_SL _19087_ (.A(_10880_),
    .B(_10881_),
    .Y(_10882_));
 NOR2x1_ASAP7_75t_SL _19090_ (.A(_00574_),
    .B(_00549_),
    .Y(_10885_));
 AO21x1_ASAP7_75t_SL _19091_ (.A1(_10882_),
    .A2(_00574_),
    .B(_10885_),
    .Y(_10886_));
 XOR2x2_ASAP7_75t_SL _19092_ (.A(_10886_),
    .B(_00862_),
    .Y(_10887_));
 AOI21x1_ASAP7_75t_SL _19093_ (.A1(_10857_),
    .A2(_10877_),
    .B(_10887_),
    .Y(_10888_));
 OAI21x1_ASAP7_75t_SL _19094_ (.A1(_10802_),
    .A2(_10837_),
    .B(_10888_),
    .Y(_10889_));
 OAI21x1_ASAP7_75t_R _19095_ (.A1(_10728_),
    .A2(_10687_),
    .B(_10723_),
    .Y(_10890_));
 NAND2x1_ASAP7_75t_SL _19096_ (.A(_10778_),
    .B(_10890_),
    .Y(_10891_));
 INVx1_ASAP7_75t_SL _19097_ (.A(_01071_),
    .Y(_10892_));
 AO21x1_ASAP7_75t_R _19098_ (.A1(_10720_),
    .A2(_10718_),
    .B(_10892_),
    .Y(_10893_));
 AOI21x1_ASAP7_75t_SL _19100_ (.A1(_10851_),
    .A2(_10893_),
    .B(_10755_),
    .Y(_10895_));
 AOI21x1_ASAP7_75t_SL _19103_ (.A1(_10895_),
    .A2(_10891_),
    .B(_10835_),
    .Y(_10898_));
 NAND3x1_ASAP7_75t_SL _19104_ (.A(_10687_),
    .B(_10723_),
    .C(_10721_),
    .Y(_10899_));
 INVx1_ASAP7_75t_SL _19105_ (.A(_10899_),
    .Y(_10900_));
 NOR2x1_ASAP7_75t_SL _19107_ (.A(_10728_),
    .B(_01067_),
    .Y(_10902_));
 NOR2x1_ASAP7_75t_SL _19108_ (.A(_10770_),
    .B(_10902_),
    .Y(_10903_));
 NOR2x1_ASAP7_75t_R _19109_ (.A(_10810_),
    .B(_10903_),
    .Y(_10904_));
 OAI21x1_ASAP7_75t_R _19110_ (.A1(_10900_),
    .A2(_10786_),
    .B(_10904_),
    .Y(_10905_));
 AOI21x1_ASAP7_75t_SL _19111_ (.A1(_10905_),
    .A2(_10898_),
    .B(_10742_),
    .Y(_10906_));
 NOR2x1_ASAP7_75t_SL _19112_ (.A(_10892_),
    .B(_10721_),
    .Y(_10907_));
 INVx1_ASAP7_75t_R _19113_ (.A(_10907_),
    .Y(_10908_));
 NAND2x1_ASAP7_75t_SL _19114_ (.A(_10721_),
    .B(_10723_),
    .Y(_10909_));
 AND3x1_ASAP7_75t_R _19116_ (.A(_10908_),
    .B(_10909_),
    .C(_10770_),
    .Y(_10911_));
 OA21x2_ASAP7_75t_SL _19117_ (.A1(_10687_),
    .A2(_10721_),
    .B(_10778_),
    .Y(_10912_));
 AO21x1_ASAP7_75t_R _19118_ (.A1(_10912_),
    .A2(_10899_),
    .B(_10755_),
    .Y(_10913_));
 NOR2x2_ASAP7_75t_L _19120_ (.A(_10728_),
    .B(_10687_),
    .Y(_10915_));
 AOI21x1_ASAP7_75t_SL _19121_ (.A1(_10778_),
    .A2(_10915_),
    .B(_10815_),
    .Y(_10916_));
 AOI21x1_ASAP7_75t_SL _19123_ (.A1(_10845_),
    .A2(_10916_),
    .B(_10875_),
    .Y(_10918_));
 OAI21x1_ASAP7_75t_R _19124_ (.A1(_10911_),
    .A2(_10913_),
    .B(_10918_),
    .Y(_10919_));
 INVx2_ASAP7_75t_SL _19125_ (.A(_10887_),
    .Y(_10920_));
 AOI21x1_ASAP7_75t_SL _19126_ (.A1(_10919_),
    .A2(_10906_),
    .B(_10920_),
    .Y(_10921_));
 OAI21x1_ASAP7_75t_SL _19127_ (.A1(_10726_),
    .A2(_10792_),
    .B(_10849_),
    .Y(_10922_));
 AO21x1_ASAP7_75t_R _19128_ (.A1(_10922_),
    .A2(_10796_),
    .B(_10778_),
    .Y(_10923_));
 AO21x1_ASAP7_75t_R _19129_ (.A1(_10869_),
    .A2(_10777_),
    .B(_10770_),
    .Y(_10924_));
 AOI21x1_ASAP7_75t_R _19132_ (.A1(_10923_),
    .A2(_10924_),
    .B(_10810_),
    .Y(_10927_));
 NOR2x1p5_ASAP7_75t_SL _19133_ (.A(_10849_),
    .B(_10728_),
    .Y(_10928_));
 NOR2x1_ASAP7_75t_SL _19134_ (.A(_10778_),
    .B(_10928_),
    .Y(_10929_));
 NOR2x1_ASAP7_75t_SL _19135_ (.A(_10755_),
    .B(_10929_),
    .Y(_10930_));
 INVx1_ASAP7_75t_SL _19136_ (.A(_10930_),
    .Y(_10931_));
 OA21x2_ASAP7_75t_R _19137_ (.A1(_10850_),
    .A2(_10915_),
    .B(_10778_),
    .Y(_10932_));
 NOR2x1_ASAP7_75t_R _19138_ (.A(_10931_),
    .B(_10932_),
    .Y(_10933_));
 OAI21x1_ASAP7_75t_R _19139_ (.A1(_10927_),
    .A2(_10933_),
    .B(_10835_),
    .Y(_10934_));
 INVx4_ASAP7_75t_SL _19140_ (.A(_10687_),
    .Y(_01061_));
 NAND2x1_ASAP7_75t_R _19141_ (.A(_10723_),
    .B(_01061_),
    .Y(_10935_));
 NOR2x1_ASAP7_75t_SL _19142_ (.A(_10770_),
    .B(_10774_),
    .Y(_10936_));
 NAND2x1_ASAP7_75t_SL _19143_ (.A(_10935_),
    .B(_10936_),
    .Y(_10937_));
 AOI21x1_ASAP7_75t_SL _19144_ (.A1(_10723_),
    .A2(_10687_),
    .B(_10778_),
    .Y(_10938_));
 AOI21x1_ASAP7_75t_R _19146_ (.A1(_10841_),
    .A2(_10938_),
    .B(_10755_),
    .Y(_10940_));
 NAND2x1_ASAP7_75t_SL _19147_ (.A(_10937_),
    .B(_10940_),
    .Y(_10941_));
 NAND2x1_ASAP7_75t_L _19148_ (.A(_01067_),
    .B(_10687_),
    .Y(_10942_));
 NOR2x1_ASAP7_75t_L _19149_ (.A(_10850_),
    .B(_10770_),
    .Y(_10943_));
 OAI21x1_ASAP7_75t_R _19150_ (.A1(_10728_),
    .A2(_10942_),
    .B(_10943_),
    .Y(_10944_));
 OAI21x1_ASAP7_75t_SL _19151_ (.A1(_10776_),
    .A2(_10721_),
    .B(_10796_),
    .Y(_10945_));
 AOI21x1_ASAP7_75t_R _19152_ (.A1(_10770_),
    .A2(_10945_),
    .B(_10810_),
    .Y(_10946_));
 AOI21x1_ASAP7_75t_R _19153_ (.A1(_10944_),
    .A2(_10946_),
    .B(_10835_),
    .Y(_10947_));
 NAND2x1_ASAP7_75t_SL _19154_ (.A(_10941_),
    .B(_10947_),
    .Y(_10948_));
 NAND3x1_ASAP7_75t_SL _19155_ (.A(_10934_),
    .B(_10948_),
    .C(_10742_),
    .Y(_10949_));
 NAND2x1_ASAP7_75t_SL _19156_ (.A(_10949_),
    .B(_10921_),
    .Y(_10950_));
 NAND2x1_ASAP7_75t_SL _19157_ (.A(_10889_),
    .B(_10950_),
    .Y(_00032_));
 NOR2x1_ASAP7_75t_SL _19158_ (.A(_10728_),
    .B(_10778_),
    .Y(_10951_));
 NAND2x1_ASAP7_75t_SL _19159_ (.A(_10803_),
    .B(_10951_),
    .Y(_10952_));
 NAND2x1_ASAP7_75t_SL _19160_ (.A(_10935_),
    .B(_10772_),
    .Y(_10953_));
 AOI21x1_ASAP7_75t_SL _19161_ (.A1(_10952_),
    .A2(_10953_),
    .B(_10810_),
    .Y(_10954_));
 NAND2x1_ASAP7_75t_SL _19162_ (.A(_10909_),
    .B(_10851_),
    .Y(_10955_));
 OAI21x1_ASAP7_75t_R _19163_ (.A1(_10726_),
    .A2(_10792_),
    .B(_10783_),
    .Y(_10956_));
 AO21x1_ASAP7_75t_SL _19164_ (.A1(_10909_),
    .A2(_10956_),
    .B(_10770_),
    .Y(_10957_));
 AOI21x1_ASAP7_75t_SL _19165_ (.A1(_10955_),
    .A2(_10957_),
    .B(_10755_),
    .Y(_10958_));
 OAI21x1_ASAP7_75t_SL _19166_ (.A1(_10954_),
    .A2(_10958_),
    .B(_10875_),
    .Y(_10959_));
 AOI21x1_ASAP7_75t_SL _19167_ (.A1(_10908_),
    .A2(_10929_),
    .B(_10810_),
    .Y(_10960_));
 NAND2x1_ASAP7_75t_SL _19168_ (.A(_10866_),
    .B(_10960_),
    .Y(_10961_));
 NOR2x1_ASAP7_75t_SL _19169_ (.A(_10721_),
    .B(_10687_),
    .Y(_10962_));
 AOI21x1_ASAP7_75t_SL _19170_ (.A1(_10721_),
    .A2(_10687_),
    .B(_10778_),
    .Y(_10963_));
 NOR2x1_ASAP7_75t_SL _19171_ (.A(_10962_),
    .B(_10963_),
    .Y(_10964_));
 AOI21x1_ASAP7_75t_SL _19173_ (.A1(_10848_),
    .A2(_10964_),
    .B(_10875_),
    .Y(_10966_));
 AOI21x1_ASAP7_75t_SL _19175_ (.A1(_10961_),
    .A2(_10966_),
    .B(_10821_),
    .Y(_10968_));
 AOI21x1_ASAP7_75t_SL _19176_ (.A1(_10959_),
    .A2(_10968_),
    .B(_10887_),
    .Y(_10969_));
 AND2x2_ASAP7_75t_SL _19177_ (.A(_10843_),
    .B(_10778_),
    .Y(_10970_));
 INVx2_ASAP7_75t_SL _19178_ (.A(_10962_),
    .Y(_10971_));
 AOI21x1_ASAP7_75t_SL _19179_ (.A1(_01071_),
    .A2(_10721_),
    .B(_10778_),
    .Y(_10972_));
 AOI21x1_ASAP7_75t_SL _19180_ (.A1(_10971_),
    .A2(_10972_),
    .B(_10755_),
    .Y(_10973_));
 INVx1_ASAP7_75t_SL _19181_ (.A(_10973_),
    .Y(_10974_));
 OA21x2_ASAP7_75t_SL _19182_ (.A1(_10956_),
    .A2(_10770_),
    .B(_10755_),
    .Y(_10975_));
 AOI21x1_ASAP7_75t_SL _19183_ (.A1(_01067_),
    .A2(_10687_),
    .B(_10728_),
    .Y(_10976_));
 OAI21x1_ASAP7_75t_SL _19184_ (.A1(_10850_),
    .A2(_10976_),
    .B(_10770_),
    .Y(_10977_));
 AOI21x1_ASAP7_75t_SL _19185_ (.A1(_10975_),
    .A2(_10977_),
    .B(_10835_),
    .Y(_10978_));
 OAI21x1_ASAP7_75t_SL _19186_ (.A1(_10970_),
    .A2(_10974_),
    .B(_10978_),
    .Y(_10979_));
 AND2x2_ASAP7_75t_SL _19187_ (.A(_10838_),
    .B(_10851_),
    .Y(_10980_));
 NOR2x1_ASAP7_75t_SL _19188_ (.A(_10770_),
    .B(_10870_),
    .Y(_10981_));
 OAI21x1_ASAP7_75t_SL _19190_ (.A1(_10980_),
    .A2(_10981_),
    .B(_10810_),
    .Y(_10983_));
 NAND2x1_ASAP7_75t_SL _19191_ (.A(_10728_),
    .B(_10723_),
    .Y(_10984_));
 AO21x1_ASAP7_75t_SL _19192_ (.A1(_10942_),
    .A2(_10984_),
    .B(_10778_),
    .Y(_10985_));
 NAND2x1_ASAP7_75t_SL _19193_ (.A(_10778_),
    .B(_10758_),
    .Y(_10986_));
 INVx1_ASAP7_75t_L _19194_ (.A(_10986_),
    .Y(_10987_));
 AOI21x1_ASAP7_75t_SL _19195_ (.A1(_10984_),
    .A2(_10987_),
    .B(_10810_),
    .Y(_10988_));
 AOI21x1_ASAP7_75t_SL _19196_ (.A1(_10985_),
    .A2(_10988_),
    .B(_10875_),
    .Y(_10989_));
 AOI21x1_ASAP7_75t_SL _19197_ (.A1(_10989_),
    .A2(_10983_),
    .B(_10742_),
    .Y(_10990_));
 NAND2x1_ASAP7_75t_SL _19198_ (.A(_10990_),
    .B(_10979_),
    .Y(_10991_));
 NAND2x1_ASAP7_75t_SL _19199_ (.A(_10969_),
    .B(_10991_),
    .Y(_10992_));
 AO21x1_ASAP7_75t_SL _19200_ (.A1(_10869_),
    .A2(_10758_),
    .B(_10778_),
    .Y(_10993_));
 AO21x1_ASAP7_75t_SL _19201_ (.A1(_10841_),
    .A2(_10794_),
    .B(_10770_),
    .Y(_10994_));
 AOI21x1_ASAP7_75t_SL _19202_ (.A1(_10993_),
    .A2(_10994_),
    .B(_10755_),
    .Y(_10995_));
 INVx1_ASAP7_75t_SL _19203_ (.A(_10915_),
    .Y(_10996_));
 NAND2x1_ASAP7_75t_SL _19204_ (.A(_10996_),
    .B(_10785_),
    .Y(_10997_));
 AO21x1_ASAP7_75t_SL _19205_ (.A1(_10984_),
    .A2(_10796_),
    .B(_10770_),
    .Y(_10998_));
 AOI21x1_ASAP7_75t_SL _19206_ (.A1(_10997_),
    .A2(_10998_),
    .B(_10810_),
    .Y(_10999_));
 OAI21x1_ASAP7_75t_SL _19207_ (.A1(_10995_),
    .A2(_10999_),
    .B(_10875_),
    .Y(_11000_));
 AO21x1_ASAP7_75t_SL _19208_ (.A1(_10727_),
    .A2(_10725_),
    .B(_01071_),
    .Y(_11001_));
 NAND2x1_ASAP7_75t_SL _19209_ (.A(_10871_),
    .B(_11001_),
    .Y(_11002_));
 AOI21x1_ASAP7_75t_SL _19210_ (.A1(_10778_),
    .A2(_11002_),
    .B(_10755_),
    .Y(_11003_));
 NAND2x1_ASAP7_75t_SL _19211_ (.A(_11003_),
    .B(_10977_),
    .Y(_11004_));
 NOR2x1_ASAP7_75t_SL _19212_ (.A(_10810_),
    .B(_10851_),
    .Y(_11005_));
 NAND3x1_ASAP7_75t_SL _19213_ (.A(_10687_),
    .B(_01067_),
    .C(_10728_),
    .Y(_11006_));
 NAND2x1_ASAP7_75t_SL _19214_ (.A(_10903_),
    .B(_11006_),
    .Y(_11007_));
 AOI21x1_ASAP7_75t_SL _19215_ (.A1(_11005_),
    .A2(_11007_),
    .B(_10875_),
    .Y(_11008_));
 AOI21x1_ASAP7_75t_SL _19216_ (.A1(_11004_),
    .A2(_11008_),
    .B(_10742_),
    .Y(_11009_));
 AOI21x1_ASAP7_75t_SL _19217_ (.A1(_11000_),
    .A2(_11009_),
    .B(_10920_),
    .Y(_11010_));
 NAND2x1_ASAP7_75t_SL _19218_ (.A(_01078_),
    .B(_10835_),
    .Y(_11011_));
 AOI21x1_ASAP7_75t_SL _19219_ (.A1(_10807_),
    .A2(_11006_),
    .B(_10810_),
    .Y(_11012_));
 OA21x2_ASAP7_75t_SL _19220_ (.A1(_10778_),
    .A2(_11011_),
    .B(_11012_),
    .Y(_11013_));
 NAND2x1_ASAP7_75t_SL _19221_ (.A(_10721_),
    .B(_10687_),
    .Y(_11014_));
 AOI21x1_ASAP7_75t_SL _19222_ (.A1(_11014_),
    .A2(_10936_),
    .B(_10875_),
    .Y(_11015_));
 NAND2x1_ASAP7_75t_SL _19223_ (.A(_10997_),
    .B(_11015_),
    .Y(_11016_));
 NAND2x1_ASAP7_75t_SL _19224_ (.A(_10770_),
    .B(_11006_),
    .Y(_11017_));
 AOI21x1_ASAP7_75t_SL _19225_ (.A1(_10868_),
    .A2(_10721_),
    .B(_10770_),
    .Y(_11018_));
 AOI21x1_ASAP7_75t_SL _19226_ (.A1(_10984_),
    .A2(_11018_),
    .B(_10835_),
    .Y(_11019_));
 OAI21x1_ASAP7_75t_SL _19227_ (.A1(_10900_),
    .A2(_11017_),
    .B(_11019_),
    .Y(_11020_));
 AOI21x1_ASAP7_75t_SL _19228_ (.A1(_11016_),
    .A2(_11020_),
    .B(_10755_),
    .Y(_11021_));
 OAI21x1_ASAP7_75t_SL _19229_ (.A1(_11013_),
    .A2(_11021_),
    .B(_10742_),
    .Y(_11022_));
 NAND2x1_ASAP7_75t_SL _19230_ (.A(_11010_),
    .B(_11022_),
    .Y(_11023_));
 NAND2x1_ASAP7_75t_SL _19231_ (.A(_10992_),
    .B(_11023_),
    .Y(_00033_));
 NOR2x1_ASAP7_75t_SL _19232_ (.A(_10854_),
    .B(_10839_),
    .Y(_11024_));
 NAND2x1_ASAP7_75t_SL _19233_ (.A(_10728_),
    .B(_10687_),
    .Y(_11025_));
 AO21x1_ASAP7_75t_SL _19234_ (.A1(_11025_),
    .A2(_10838_),
    .B(_10778_),
    .Y(_11026_));
 NAND2x1_ASAP7_75t_SL _19235_ (.A(_11024_),
    .B(_11026_),
    .Y(_11027_));
 NAND2x1_ASAP7_75t_L _19236_ (.A(_10770_),
    .B(_10838_),
    .Y(_11028_));
 OAI21x1_ASAP7_75t_R _19237_ (.A1(_10719_),
    .A2(_10795_),
    .B(_10892_),
    .Y(_11029_));
 NAND2x1p5_ASAP7_75t_L _19238_ (.A(_10778_),
    .B(_11029_),
    .Y(_11030_));
 OAI21x1_ASAP7_75t_SL _19239_ (.A1(_10774_),
    .A2(_11028_),
    .B(_11030_),
    .Y(_11031_));
 NOR2x1_ASAP7_75t_SL _19240_ (.A(_10755_),
    .B(_10854_),
    .Y(_11032_));
 AOI21x1_ASAP7_75t_SL _19241_ (.A1(_11031_),
    .A2(_11032_),
    .B(_10875_),
    .Y(_11033_));
 NAND2x1_ASAP7_75t_SL _19242_ (.A(_11027_),
    .B(_11033_),
    .Y(_11034_));
 NAND2x1_ASAP7_75t_R _19243_ (.A(_10770_),
    .B(_10852_),
    .Y(_11035_));
 NOR2x1_ASAP7_75t_SL _19244_ (.A(_10915_),
    .B(_11035_),
    .Y(_11036_));
 OAI21x1_ASAP7_75t_SL _19245_ (.A1(_10774_),
    .A2(_11030_),
    .B(_10810_),
    .Y(_11037_));
 NOR2x1_ASAP7_75t_SL _19246_ (.A(_11036_),
    .B(_11037_),
    .Y(_11038_));
 NOR2x1_ASAP7_75t_R _19247_ (.A(_10818_),
    .B(_10770_),
    .Y(_11039_));
 NAND2x1_ASAP7_75t_SL _19248_ (.A(_10984_),
    .B(_11039_),
    .Y(_11040_));
 NAND2x1_ASAP7_75t_SL _19249_ (.A(_10758_),
    .B(_10851_),
    .Y(_11041_));
 AOI21x1_ASAP7_75t_SL _19250_ (.A1(_11040_),
    .A2(_11041_),
    .B(_10810_),
    .Y(_11042_));
 OAI21x1_ASAP7_75t_SL _19251_ (.A1(_11038_),
    .A2(_11042_),
    .B(_10875_),
    .Y(_11043_));
 AOI21x1_ASAP7_75t_SL _19252_ (.A1(_11034_),
    .A2(_11043_),
    .B(_10742_),
    .Y(_11044_));
 OAI21x1_ASAP7_75t_SL _19253_ (.A1(_10863_),
    .A2(_10864_),
    .B(_10770_),
    .Y(_11045_));
 AO21x1_ASAP7_75t_SL _19254_ (.A1(_11025_),
    .A2(_10758_),
    .B(_10770_),
    .Y(_11046_));
 AOI21x1_ASAP7_75t_SL _19255_ (.A1(_11045_),
    .A2(_11046_),
    .B(_10810_),
    .Y(_11047_));
 OAI21x1_ASAP7_75t_SL _19256_ (.A1(_10723_),
    .A2(_10728_),
    .B(_10687_),
    .Y(_11048_));
 AOI21x1_ASAP7_75t_R _19257_ (.A1(_11029_),
    .A2(_10956_),
    .B(_10770_),
    .Y(_11049_));
 AOI21x1_ASAP7_75t_SL _19258_ (.A1(_10770_),
    .A2(_11048_),
    .B(_11049_),
    .Y(_11050_));
 OAI21x1_ASAP7_75t_SL _19259_ (.A1(_10755_),
    .A2(_11050_),
    .B(_10835_),
    .Y(_11051_));
 NOR2x1_ASAP7_75t_SL _19260_ (.A(_11047_),
    .B(_11051_),
    .Y(_11052_));
 INVx1_ASAP7_75t_R _19261_ (.A(_10871_),
    .Y(_11053_));
 NOR3x1_ASAP7_75t_SL _19262_ (.A(_10774_),
    .B(_11053_),
    .C(_10778_),
    .Y(_11054_));
 NAND2x1_ASAP7_75t_SL _19263_ (.A(_10778_),
    .B(_10922_),
    .Y(_11055_));
 OAI21x1_ASAP7_75t_SL _19264_ (.A1(_10915_),
    .A2(_11055_),
    .B(_10810_),
    .Y(_11056_));
 OAI21x1_ASAP7_75t_SL _19265_ (.A1(_11054_),
    .A2(_11056_),
    .B(_10875_),
    .Y(_11057_));
 AOI21x1_ASAP7_75t_SL _19266_ (.A1(_10687_),
    .A2(_10902_),
    .B(_10770_),
    .Y(_11058_));
 INVx1_ASAP7_75t_SL _19267_ (.A(_11058_),
    .Y(_11059_));
 INVx1_ASAP7_75t_R _19268_ (.A(_11001_),
    .Y(_11060_));
 OAI21x1_ASAP7_75t_SL _19269_ (.A1(_11060_),
    .A2(_10976_),
    .B(_10770_),
    .Y(_11061_));
 AOI21x1_ASAP7_75t_SL _19270_ (.A1(_11059_),
    .A2(_11061_),
    .B(_10810_),
    .Y(_11062_));
 OAI21x1_ASAP7_75t_SL _19271_ (.A1(_11057_),
    .A2(_11062_),
    .B(_10742_),
    .Y(_11063_));
 NOR2x1_ASAP7_75t_SL _19272_ (.A(_11052_),
    .B(_11063_),
    .Y(_11064_));
 OAI21x1_ASAP7_75t_SL _19273_ (.A1(_11044_),
    .A2(_11064_),
    .B(_10887_),
    .Y(_11065_));
 NOR2x1_ASAP7_75t_SL _19274_ (.A(_10770_),
    .B(_11011_),
    .Y(_11066_));
 AOI21x1_ASAP7_75t_R _19275_ (.A1(_10723_),
    .A2(_01061_),
    .B(_10778_),
    .Y(_11067_));
 AOI21x1_ASAP7_75t_SL _19276_ (.A1(_11025_),
    .A2(_11067_),
    .B(_10810_),
    .Y(_11068_));
 NOR2x1_ASAP7_75t_SL _19277_ (.A(_10875_),
    .B(_11068_),
    .Y(_11069_));
 NOR2x1_ASAP7_75t_SL _19278_ (.A(_10776_),
    .B(_10721_),
    .Y(_11070_));
 NOR3x1_ASAP7_75t_SL _19279_ (.A(_11070_),
    .B(_10860_),
    .C(_10778_),
    .Y(_11071_));
 AND2x2_ASAP7_75t_SL _19280_ (.A(_10772_),
    .B(_10796_),
    .Y(_11072_));
 OAI21x1_ASAP7_75t_SL _19281_ (.A1(_11071_),
    .A2(_11072_),
    .B(_10810_),
    .Y(_11073_));
 OAI21x1_ASAP7_75t_SL _19282_ (.A1(_11066_),
    .A2(_11069_),
    .B(_11073_),
    .Y(_11074_));
 OAI21x1_ASAP7_75t_SL _19283_ (.A1(_10728_),
    .A2(_10687_),
    .B(_10770_),
    .Y(_11075_));
 INVx1_ASAP7_75t_SL _19284_ (.A(_11075_),
    .Y(_11076_));
 NAND2x1_ASAP7_75t_SL _19285_ (.A(_10984_),
    .B(_11076_),
    .Y(_11077_));
 NAND3x1_ASAP7_75t_SL _19286_ (.A(_11077_),
    .B(_10810_),
    .C(_10773_),
    .Y(_11078_));
 OA21x2_ASAP7_75t_SL _19287_ (.A1(_10770_),
    .A2(_01076_),
    .B(_10755_),
    .Y(_11079_));
 NAND2x1_ASAP7_75t_SL _19288_ (.A(_10929_),
    .B(_10805_),
    .Y(_11080_));
 AOI21x1_ASAP7_75t_SL _19289_ (.A1(_11079_),
    .A2(_11080_),
    .B(_10835_),
    .Y(_11081_));
 AOI21x1_ASAP7_75t_SL _19290_ (.A1(_11078_),
    .A2(_11081_),
    .B(_10742_),
    .Y(_11082_));
 NAND2x1_ASAP7_75t_SL _19291_ (.A(_11074_),
    .B(_11082_),
    .Y(_11083_));
 AO21x1_ASAP7_75t_SL _19292_ (.A1(_10922_),
    .A2(_10838_),
    .B(_10778_),
    .Y(_11084_));
 NOR2x1_ASAP7_75t_R _19293_ (.A(_10770_),
    .B(_10869_),
    .Y(_11085_));
 NOR2x1_ASAP7_75t_SL _19294_ (.A(_10835_),
    .B(_11085_),
    .Y(_11086_));
 AOI21x1_ASAP7_75t_SL _19295_ (.A1(_11084_),
    .A2(_11086_),
    .B(_10810_),
    .Y(_11087_));
 AND2x2_ASAP7_75t_SL _19296_ (.A(_10770_),
    .B(_01075_),
    .Y(_11088_));
 NOR2x1_ASAP7_75t_SL _19297_ (.A(_11088_),
    .B(_11058_),
    .Y(_11089_));
 NAND2x1_ASAP7_75t_SL _19298_ (.A(_10835_),
    .B(_11089_),
    .Y(_11090_));
 NAND2x1_ASAP7_75t_SL _19299_ (.A(_11087_),
    .B(_11090_),
    .Y(_11091_));
 NAND2x1_ASAP7_75t_SL _19300_ (.A(_10770_),
    .B(_11048_),
    .Y(_11092_));
 OA21x2_ASAP7_75t_SL _19301_ (.A1(_01080_),
    .A2(_10770_),
    .B(_10835_),
    .Y(_11093_));
 AOI21x1_ASAP7_75t_SL _19302_ (.A1(_11092_),
    .A2(_11093_),
    .B(_10755_),
    .Y(_11094_));
 NOR2x1_ASAP7_75t_SL _19303_ (.A(_10778_),
    .B(_10794_),
    .Y(_11095_));
 AOI21x1_ASAP7_75t_SL _19304_ (.A1(_10942_),
    .A2(_10951_),
    .B(_11095_),
    .Y(_11096_));
 NOR2x1_ASAP7_75t_SL _19305_ (.A(_10721_),
    .B(_10778_),
    .Y(_11097_));
 AOI21x1_ASAP7_75t_SL _19306_ (.A1(_10783_),
    .A2(_11097_),
    .B(_10835_),
    .Y(_11098_));
 OAI21x1_ASAP7_75t_SL _19307_ (.A1(_10721_),
    .A2(_10942_),
    .B(_10807_),
    .Y(_11099_));
 NAND3x1_ASAP7_75t_SL _19308_ (.A(_11096_),
    .B(_11098_),
    .C(_11099_),
    .Y(_11100_));
 AOI21x1_ASAP7_75t_SL _19309_ (.A1(_11094_),
    .A2(_11100_),
    .B(_10821_),
    .Y(_11101_));
 AOI21x1_ASAP7_75t_SL _19310_ (.A1(_11091_),
    .A2(_11101_),
    .B(_10887_),
    .Y(_11102_));
 NAND2x1_ASAP7_75t_SL _19311_ (.A(_11083_),
    .B(_11102_),
    .Y(_11103_));
 NAND2x1_ASAP7_75t_SL _19312_ (.A(_11065_),
    .B(_11103_),
    .Y(_00034_));
 NAND2x1_ASAP7_75t_SL _19313_ (.A(_10893_),
    .B(_10943_),
    .Y(_11104_));
 AO21x1_ASAP7_75t_SL _19314_ (.A1(_10909_),
    .A2(_10852_),
    .B(_10778_),
    .Y(_11105_));
 AOI21x1_ASAP7_75t_SL _19315_ (.A1(_11104_),
    .A2(_11105_),
    .B(_10755_),
    .Y(_11106_));
 AO21x1_ASAP7_75t_SL _19316_ (.A1(_10841_),
    .A2(_10869_),
    .B(_10778_),
    .Y(_11107_));
 AOI21x1_ASAP7_75t_SL _19317_ (.A1(_10953_),
    .A2(_11107_),
    .B(_10810_),
    .Y(_11108_));
 OAI21x1_ASAP7_75t_SL _19318_ (.A1(_11106_),
    .A2(_11108_),
    .B(_10875_),
    .Y(_11109_));
 NOR2x1_ASAP7_75t_SL _19319_ (.A(_10774_),
    .B(_11030_),
    .Y(_11110_));
 AOI21x1_ASAP7_75t_SL _19320_ (.A1(_10810_),
    .A2(_11110_),
    .B(_10875_),
    .Y(_11111_));
 NAND2x1_ASAP7_75t_SL _19321_ (.A(_01064_),
    .B(_10784_),
    .Y(_11112_));
 NAND2x1_ASAP7_75t_SL _19322_ (.A(_10819_),
    .B(_11112_),
    .Y(_11113_));
 NAND2x1_ASAP7_75t_SL _19323_ (.A(_11113_),
    .B(_11012_),
    .Y(_11114_));
 AOI21x1_ASAP7_75t_SL _19324_ (.A1(_11111_),
    .A2(_11114_),
    .B(_10742_),
    .Y(_11115_));
 AOI21x1_ASAP7_75t_SL _19325_ (.A1(_11109_),
    .A2(_11115_),
    .B(_10920_),
    .Y(_11116_));
 OA21x2_ASAP7_75t_SL _19326_ (.A1(_10778_),
    .A2(_10852_),
    .B(_10875_),
    .Y(_11117_));
 AOI21x1_ASAP7_75t_SL _19327_ (.A1(_11040_),
    .A2(_11117_),
    .B(_10810_),
    .Y(_11118_));
 OAI21x1_ASAP7_75t_R _19328_ (.A1(_10793_),
    .A2(_10783_),
    .B(_10728_),
    .Y(_11119_));
 AO21x1_ASAP7_75t_SL _19329_ (.A1(_11119_),
    .A2(_11029_),
    .B(_10778_),
    .Y(_11120_));
 AO21x1_ASAP7_75t_SL _19330_ (.A1(_10841_),
    .A2(_10922_),
    .B(_10770_),
    .Y(_11121_));
 NAND3x1_ASAP7_75t_SL _19331_ (.A(_11120_),
    .B(_11121_),
    .C(_10835_),
    .Y(_11122_));
 AOI21x1_ASAP7_75t_SL _19332_ (.A1(_11118_),
    .A2(_11122_),
    .B(_10821_),
    .Y(_11123_));
 NAND2x1_ASAP7_75t_SL _19333_ (.A(_11025_),
    .B(_10807_),
    .Y(_11124_));
 NAND2x1_ASAP7_75t_SL _19334_ (.A(_10770_),
    .B(_10928_),
    .Y(_11125_));
 AO21x1_ASAP7_75t_SL _19335_ (.A1(_11124_),
    .A2(_11125_),
    .B(_10875_),
    .Y(_11126_));
 NAND2x1p5_ASAP7_75t_SL _19336_ (.A(_10850_),
    .B(_10778_),
    .Y(_11127_));
 OA22x2_ASAP7_75t_SL _19337_ (.A1(_10778_),
    .A2(_10794_),
    .B1(_11127_),
    .B2(_10835_),
    .Y(_11128_));
 AO21x1_ASAP7_75t_SL _19338_ (.A1(_11126_),
    .A2(_11128_),
    .B(_10755_),
    .Y(_11129_));
 NAND2x1_ASAP7_75t_SL _19339_ (.A(_11123_),
    .B(_11129_),
    .Y(_11130_));
 NAND2x1_ASAP7_75t_SL _19340_ (.A(_11116_),
    .B(_11130_),
    .Y(_11131_));
 AO21x1_ASAP7_75t_SL _19341_ (.A1(_01069_),
    .A2(_10721_),
    .B(_11055_),
    .Y(_11132_));
 NAND2x1_ASAP7_75t_SL _19342_ (.A(_11132_),
    .B(_10973_),
    .Y(_11133_));
 INVx1_ASAP7_75t_SL _19343_ (.A(_11097_),
    .Y(_11134_));
 AOI211x1_ASAP7_75t_SL _19344_ (.A1(_01061_),
    .A2(_10723_),
    .B(_10842_),
    .C(_10810_),
    .Y(_11135_));
 NAND2x1_ASAP7_75t_SL _19345_ (.A(_11134_),
    .B(_11135_),
    .Y(_11136_));
 AOI21x1_ASAP7_75t_SL _19346_ (.A1(_11133_),
    .A2(_11136_),
    .B(_10875_),
    .Y(_11137_));
 OAI21x1_ASAP7_75t_SL _19347_ (.A1(_10986_),
    .A2(_10843_),
    .B(_10755_),
    .Y(_11138_));
 OAI21x1_ASAP7_75t_SL _19348_ (.A1(_10776_),
    .A2(_10721_),
    .B(_10841_),
    .Y(_11139_));
 NOR2x1_ASAP7_75t_SL _19349_ (.A(_11075_),
    .B(_11139_),
    .Y(_11140_));
 NOR2x1_ASAP7_75t_SL _19350_ (.A(_11138_),
    .B(_11140_),
    .Y(_11141_));
 INVx1_ASAP7_75t_SL _19351_ (.A(_10777_),
    .Y(_11142_));
 INVx2_ASAP7_75t_SL _19352_ (.A(_10850_),
    .Y(_11143_));
 NAND2x1_ASAP7_75t_SL _19353_ (.A(_10778_),
    .B(_11143_),
    .Y(_11144_));
 OAI21x1_ASAP7_75t_SL _19354_ (.A1(_11142_),
    .A2(_11144_),
    .B(_10810_),
    .Y(_11145_));
 AOI21x1_ASAP7_75t_SL _19355_ (.A1(_10775_),
    .A2(_10935_),
    .B(_10778_),
    .Y(_11146_));
 OAI21x1_ASAP7_75t_SL _19356_ (.A1(_11145_),
    .A2(_11146_),
    .B(_10875_),
    .Y(_11147_));
 OAI21x1_ASAP7_75t_SL _19357_ (.A1(_11141_),
    .A2(_11147_),
    .B(_10821_),
    .Y(_11148_));
 NOR2x1_ASAP7_75t_SL _19358_ (.A(_11137_),
    .B(_11148_),
    .Y(_11149_));
 AO21x1_ASAP7_75t_SL _19359_ (.A1(_10775_),
    .A2(_11014_),
    .B(_10770_),
    .Y(_11150_));
 NAND2x1_ASAP7_75t_SL _19360_ (.A(_10930_),
    .B(_11150_),
    .Y(_11151_));
 NAND2x1_ASAP7_75t_SL _19361_ (.A(_10803_),
    .B(_10936_),
    .Y(_11152_));
 AOI21x1_ASAP7_75t_SL _19362_ (.A1(_10851_),
    .A2(_10996_),
    .B(_10810_),
    .Y(_11153_));
 AOI21x1_ASAP7_75t_SL _19363_ (.A1(_11152_),
    .A2(_11153_),
    .B(_10875_),
    .Y(_11154_));
 NAND2x1_ASAP7_75t_SL _19364_ (.A(_11151_),
    .B(_11154_),
    .Y(_11155_));
 INVx1_ASAP7_75t_SL _19365_ (.A(_10869_),
    .Y(_11156_));
 OAI21x1_ASAP7_75t_SL _19366_ (.A1(_10928_),
    .A2(_11156_),
    .B(_10770_),
    .Y(_11157_));
 OAI21x1_ASAP7_75t_SL _19367_ (.A1(_11070_),
    .A2(_10842_),
    .B(_10778_),
    .Y(_11158_));
 AOI21x1_ASAP7_75t_SL _19368_ (.A1(_11157_),
    .A2(_11158_),
    .B(_10755_),
    .Y(_11159_));
 AO21x1_ASAP7_75t_SL _19369_ (.A1(_11001_),
    .A2(_10838_),
    .B(_10778_),
    .Y(_11160_));
 INVx1_ASAP7_75t_SL _19370_ (.A(_11055_),
    .Y(_11161_));
 NAND2x1_ASAP7_75t_SL _19371_ (.A(_10996_),
    .B(_11161_),
    .Y(_11162_));
 AOI21x1_ASAP7_75t_SL _19372_ (.A1(_11160_),
    .A2(_11162_),
    .B(_10810_),
    .Y(_11163_));
 OAI21x1_ASAP7_75t_SL _19373_ (.A1(_11159_),
    .A2(_11163_),
    .B(_10875_),
    .Y(_11164_));
 AOI21x1_ASAP7_75t_SL _19374_ (.A1(_11155_),
    .A2(_11164_),
    .B(_10821_),
    .Y(_11165_));
 OAI21x1_ASAP7_75t_SL _19375_ (.A1(_11149_),
    .A2(_11165_),
    .B(_10920_),
    .Y(_11166_));
 NAND2x1_ASAP7_75t_SL _19376_ (.A(_11131_),
    .B(_11166_),
    .Y(_00035_));
 AO21x1_ASAP7_75t_SL _19377_ (.A1(_01066_),
    .A2(_10728_),
    .B(_10770_),
    .Y(_11167_));
 NOR2x1_ASAP7_75t_SL _19378_ (.A(_10860_),
    .B(_11167_),
    .Y(_11168_));
 NAND2x1_ASAP7_75t_SL _19379_ (.A(_10755_),
    .B(_10845_),
    .Y(_11169_));
 OAI21x1_ASAP7_75t_SL _19380_ (.A1(_10728_),
    .A2(_10942_),
    .B(_10770_),
    .Y(_11170_));
 NOR2x1_ASAP7_75t_SL _19381_ (.A(_10793_),
    .B(_10728_),
    .Y(_11171_));
 OA21x2_ASAP7_75t_SL _19382_ (.A1(_11171_),
    .A2(_10770_),
    .B(_10810_),
    .Y(_11172_));
 AOI21x1_ASAP7_75t_SL _19383_ (.A1(_11170_),
    .A2(_11172_),
    .B(_10835_),
    .Y(_11173_));
 OAI21x1_ASAP7_75t_SL _19384_ (.A1(_11168_),
    .A2(_11169_),
    .B(_11173_),
    .Y(_11174_));
 NOR2x1_ASAP7_75t_SL _19385_ (.A(_10810_),
    .B(_10951_),
    .Y(_11175_));
 AO21x1_ASAP7_75t_SL _19386_ (.A1(_10984_),
    .A2(_11029_),
    .B(_10770_),
    .Y(_11176_));
 AOI21x1_ASAP7_75t_SL _19387_ (.A1(_11175_),
    .A2(_11176_),
    .B(_10875_),
    .Y(_11177_));
 AOI21x1_ASAP7_75t_SL _19388_ (.A1(_10778_),
    .A2(_10915_),
    .B(_10755_),
    .Y(_11178_));
 AOI21x1_ASAP7_75t_SL _19389_ (.A1(_10996_),
    .A2(_10785_),
    .B(_11085_),
    .Y(_11179_));
 NAND2x1_ASAP7_75t_SL _19390_ (.A(_11178_),
    .B(_11179_),
    .Y(_11180_));
 AOI21x1_ASAP7_75t_SL _19391_ (.A1(_11177_),
    .A2(_11180_),
    .B(_10742_),
    .Y(_11181_));
 AOI21x1_ASAP7_75t_SL _19392_ (.A1(_11174_),
    .A2(_11181_),
    .B(_10920_),
    .Y(_11182_));
 OAI21x1_ASAP7_75t_SL _19393_ (.A1(_10818_),
    .A2(_10774_),
    .B(_10770_),
    .Y(_11183_));
 NAND2x1_ASAP7_75t_SL _19394_ (.A(_10942_),
    .B(_10912_),
    .Y(_11184_));
 AOI21x1_ASAP7_75t_SL _19395_ (.A1(_11183_),
    .A2(_11184_),
    .B(_10755_),
    .Y(_11185_));
 AOI21x1_ASAP7_75t_SL _19396_ (.A1(_10841_),
    .A2(_10938_),
    .B(_10810_),
    .Y(_11186_));
 AO21x1_ASAP7_75t_SL _19397_ (.A1(_11186_),
    .A2(_10798_),
    .B(_10875_),
    .Y(_11187_));
 NAND2x1_ASAP7_75t_SL _19398_ (.A(_10778_),
    .B(_10864_),
    .Y(_11188_));
 AOI21x1_ASAP7_75t_SL _19399_ (.A1(_10819_),
    .A2(_10971_),
    .B(_10755_),
    .Y(_11189_));
 NAND2x1_ASAP7_75t_SL _19400_ (.A(_11188_),
    .B(_11189_),
    .Y(_11190_));
 AO21x1_ASAP7_75t_SL _19401_ (.A1(_10778_),
    .A2(_01070_),
    .B(_10810_),
    .Y(_11191_));
 NOR2x1_ASAP7_75t_SL _19402_ (.A(_10778_),
    .B(_10860_),
    .Y(_11192_));
 OA21x2_ASAP7_75t_SL _19403_ (.A1(_11191_),
    .A2(_11192_),
    .B(_10875_),
    .Y(_11193_));
 AOI21x1_ASAP7_75t_SL _19404_ (.A1(_11190_),
    .A2(_11193_),
    .B(_10821_),
    .Y(_11194_));
 OAI21x1_ASAP7_75t_SL _19405_ (.A1(_11185_),
    .A2(_11187_),
    .B(_11194_),
    .Y(_11195_));
 NAND2x1_ASAP7_75t_SL _19406_ (.A(_11182_),
    .B(_11195_),
    .Y(_11196_));
 OA21x2_ASAP7_75t_SL _19407_ (.A1(_10758_),
    .A2(_10778_),
    .B(_10852_),
    .Y(_11197_));
 AOI21x1_ASAP7_75t_SL _19408_ (.A1(_10848_),
    .A2(_11197_),
    .B(_10835_),
    .Y(_11198_));
 INVx1_ASAP7_75t_SL _19409_ (.A(_10928_),
    .Y(_11199_));
 NOR2x1_ASAP7_75t_SL _19410_ (.A(_10770_),
    .B(_10907_),
    .Y(_11200_));
 AOI21x1_ASAP7_75t_SL _19411_ (.A1(_11199_),
    .A2(_11200_),
    .B(_10810_),
    .Y(_11201_));
 NAND2x1_ASAP7_75t_SL _19412_ (.A(_10820_),
    .B(_11201_),
    .Y(_11202_));
 AOI21x1_ASAP7_75t_SL _19413_ (.A1(_11198_),
    .A2(_11202_),
    .B(_10821_),
    .Y(_11203_));
 AO21x1_ASAP7_75t_SL _19414_ (.A1(_11156_),
    .A2(_10770_),
    .B(_10810_),
    .Y(_11204_));
 NAND2x1_ASAP7_75t_SL _19415_ (.A(_10770_),
    .B(_10687_),
    .Y(_11205_));
 OAI21x1_ASAP7_75t_SL _19416_ (.A1(_10728_),
    .A2(_11205_),
    .B(_10866_),
    .Y(_11206_));
 NOR2x1_ASAP7_75t_SL _19417_ (.A(_10755_),
    .B(_11049_),
    .Y(_11207_));
 INVx1_ASAP7_75t_SL _19418_ (.A(_11014_),
    .Y(_11208_));
 OAI21x1_ASAP7_75t_SL _19419_ (.A1(_11208_),
    .A2(_10864_),
    .B(_10770_),
    .Y(_11209_));
 AOI21x1_ASAP7_75t_SL _19420_ (.A1(_11207_),
    .A2(_11209_),
    .B(_10875_),
    .Y(_11210_));
 OAI21x1_ASAP7_75t_SL _19421_ (.A1(_11204_),
    .A2(_11206_),
    .B(_11210_),
    .Y(_11211_));
 AOI21x1_ASAP7_75t_SL _19422_ (.A1(_11203_),
    .A2(_11211_),
    .B(_10887_),
    .Y(_11212_));
 AOI21x1_ASAP7_75t_SL _19423_ (.A1(_10984_),
    .A2(_10963_),
    .B(_10810_),
    .Y(_11213_));
 NOR2x1_ASAP7_75t_SL _19424_ (.A(_10755_),
    .B(_10835_),
    .Y(_11214_));
 INVx1_ASAP7_75t_SL _19425_ (.A(_10819_),
    .Y(_11215_));
 AND3x1_ASAP7_75t_SL _19426_ (.A(_11214_),
    .B(_10794_),
    .C(_11215_),
    .Y(_11216_));
 AO21x1_ASAP7_75t_SL _19427_ (.A1(_11019_),
    .A2(_11213_),
    .B(_11216_),
    .Y(_11217_));
 NAND2x1_ASAP7_75t_SL _19428_ (.A(_11014_),
    .B(_10936_),
    .Y(_11218_));
 NAND2x1_ASAP7_75t_SL _19429_ (.A(_11218_),
    .B(_11068_),
    .Y(_11219_));
 AO21x1_ASAP7_75t_SL _19430_ (.A1(_11025_),
    .A2(_10796_),
    .B(_10778_),
    .Y(_11220_));
 AOI21x1_ASAP7_75t_SL _19431_ (.A1(_10942_),
    .A2(_10912_),
    .B(_10755_),
    .Y(_11221_));
 NAND2x1_ASAP7_75t_SL _19432_ (.A(_11220_),
    .B(_11221_),
    .Y(_11222_));
 AOI21x1_ASAP7_75t_SL _19433_ (.A1(_11219_),
    .A2(_11222_),
    .B(_10875_),
    .Y(_11223_));
 OAI21x1_ASAP7_75t_SL _19434_ (.A1(_11217_),
    .A2(_11223_),
    .B(_10821_),
    .Y(_11224_));
 NAND2x1_ASAP7_75t_SL _19435_ (.A(_11212_),
    .B(_11224_),
    .Y(_11225_));
 NAND2x1_ASAP7_75t_SL _19436_ (.A(_11196_),
    .B(_11225_),
    .Y(_00036_));
 OAI21x1_ASAP7_75t_SL _19437_ (.A1(_11053_),
    .A2(_10962_),
    .B(_10778_),
    .Y(_11226_));
 OA21x2_ASAP7_75t_SL _19438_ (.A1(_10758_),
    .A2(_10778_),
    .B(_10810_),
    .Y(_11227_));
 AOI21x1_ASAP7_75t_SL _19439_ (.A1(_11226_),
    .A2(_11227_),
    .B(_10875_),
    .Y(_11228_));
 NAND2x1p5_ASAP7_75t_SL _19440_ (.A(_10851_),
    .B(_10796_),
    .Y(_11229_));
 AO21x1_ASAP7_75t_SL _19441_ (.A1(_11030_),
    .A2(_11229_),
    .B(_10810_),
    .Y(_11230_));
 AOI21x1_ASAP7_75t_SL _19442_ (.A1(_11228_),
    .A2(_11230_),
    .B(_10821_),
    .Y(_11231_));
 OAI21x1_ASAP7_75t_SL _19443_ (.A1(_11142_),
    .A2(_10843_),
    .B(_10770_),
    .Y(_11232_));
 AO21x1_ASAP7_75t_SL _19444_ (.A1(_10942_),
    .A2(_10909_),
    .B(_10770_),
    .Y(_11233_));
 AOI21x1_ASAP7_75t_SL _19445_ (.A1(_11232_),
    .A2(_11233_),
    .B(_10755_),
    .Y(_11234_));
 AOI21x1_ASAP7_75t_SL _19446_ (.A1(_11205_),
    .A2(_11184_),
    .B(_10810_),
    .Y(_11235_));
 OAI21x1_ASAP7_75t_SL _19447_ (.A1(_11234_),
    .A2(_11235_),
    .B(_10875_),
    .Y(_11236_));
 NAND2x1_ASAP7_75t_SL _19448_ (.A(_11236_),
    .B(_11231_),
    .Y(_11237_));
 NAND3x1_ASAP7_75t_SL _19449_ (.A(_10952_),
    .B(_11167_),
    .C(_10810_),
    .Y(_11238_));
 NAND2x1_ASAP7_75t_SL _19450_ (.A(_11127_),
    .B(_11035_),
    .Y(_11239_));
 AOI21x1_ASAP7_75t_SL _19451_ (.A1(_10723_),
    .A2(_10951_),
    .B(_10810_),
    .Y(_11240_));
 AOI21x1_ASAP7_75t_SL _19452_ (.A1(_11239_),
    .A2(_11240_),
    .B(_10875_),
    .Y(_11241_));
 AOI21x1_ASAP7_75t_SL _19453_ (.A1(_11238_),
    .A2(_11241_),
    .B(_10742_),
    .Y(_11242_));
 INVx1_ASAP7_75t_SL _19454_ (.A(_10972_),
    .Y(_11243_));
 OAI21x1_ASAP7_75t_SL _19455_ (.A1(_11243_),
    .A2(_10784_),
    .B(_10916_),
    .Y(_11244_));
 OAI21x1_ASAP7_75t_SL _19456_ (.A1(_10721_),
    .A2(_10803_),
    .B(_11039_),
    .Y(_11245_));
 AOI211x1_ASAP7_75t_SL _19457_ (.A1(_10783_),
    .A2(_10770_),
    .B(_11095_),
    .C(_10755_),
    .Y(_11246_));
 AOI21x1_ASAP7_75t_SL _19458_ (.A1(_11245_),
    .A2(_11246_),
    .B(_10835_),
    .Y(_11247_));
 NAND2x1_ASAP7_75t_SL _19459_ (.A(_11244_),
    .B(_11247_),
    .Y(_11248_));
 AOI21x1_ASAP7_75t_SL _19460_ (.A1(_11242_),
    .A2(_11248_),
    .B(_10887_),
    .Y(_11249_));
 NAND2x1_ASAP7_75t_SL _19461_ (.A(_11237_),
    .B(_11249_),
    .Y(_11250_));
 NAND2x1_ASAP7_75t_SL _19462_ (.A(_10778_),
    .B(_10774_),
    .Y(_11251_));
 AND3x1_ASAP7_75t_SL _19463_ (.A(_10845_),
    .B(_10840_),
    .C(_11251_),
    .Y(_11252_));
 AO21x1_ASAP7_75t_SL _19464_ (.A1(_11142_),
    .A2(_10770_),
    .B(_10755_),
    .Y(_11253_));
 AND3x1_ASAP7_75t_SL _19465_ (.A(_11006_),
    .B(_10778_),
    .C(_10893_),
    .Y(_11254_));
 OAI21x1_ASAP7_75t_SL _19466_ (.A1(_11253_),
    .A2(_11254_),
    .B(_10835_),
    .Y(_11255_));
 NOR2x1_ASAP7_75t_SL _19467_ (.A(_11252_),
    .B(_11255_),
    .Y(_11256_));
 OA21x2_ASAP7_75t_SL _19468_ (.A1(_10778_),
    .A2(_10723_),
    .B(_10755_),
    .Y(_11257_));
 AO21x1_ASAP7_75t_SL _19469_ (.A1(_10937_),
    .A2(_11257_),
    .B(_10835_),
    .Y(_11258_));
 INVx2_ASAP7_75t_SL _19470_ (.A(_10851_),
    .Y(_11259_));
 AOI21x1_ASAP7_75t_SL _19471_ (.A1(_11039_),
    .A2(_10971_),
    .B(_10755_),
    .Y(_11260_));
 OA21x2_ASAP7_75t_SL _19472_ (.A1(_10900_),
    .A2(_11259_),
    .B(_11260_),
    .Y(_11261_));
 OAI21x1_ASAP7_75t_SL _19473_ (.A1(_11258_),
    .A2(_11261_),
    .B(_10821_),
    .Y(_11262_));
 NOR2x1_ASAP7_75t_SL _19474_ (.A(_10806_),
    .B(_11259_),
    .Y(_11263_));
 AO21x1_ASAP7_75t_SL _19475_ (.A1(_11161_),
    .A2(_10893_),
    .B(_10755_),
    .Y(_11264_));
 OA21x2_ASAP7_75t_SL _19476_ (.A1(_10778_),
    .A2(_10776_),
    .B(_10755_),
    .Y(_11265_));
 NOR2x1_ASAP7_75t_SL _19477_ (.A(_01067_),
    .B(_10770_),
    .Y(_11266_));
 NOR2x1_ASAP7_75t_SL _19478_ (.A(_11266_),
    .B(_10772_),
    .Y(_11267_));
 AOI21x1_ASAP7_75t_SL _19479_ (.A1(_11265_),
    .A2(_11267_),
    .B(_10875_),
    .Y(_11268_));
 OAI21x1_ASAP7_75t_SL _19480_ (.A1(_11263_),
    .A2(_11264_),
    .B(_11268_),
    .Y(_11269_));
 AOI21x1_ASAP7_75t_SL _19481_ (.A1(_11243_),
    .A2(_10848_),
    .B(_10835_),
    .Y(_11270_));
 AOI21x1_ASAP7_75t_SL _19482_ (.A1(_10770_),
    .A2(_11112_),
    .B(_10810_),
    .Y(_11271_));
 NAND2x1_ASAP7_75t_SL _19483_ (.A(_11006_),
    .B(_11058_),
    .Y(_11272_));
 NAND2x1_ASAP7_75t_SL _19484_ (.A(_11271_),
    .B(_11272_),
    .Y(_11273_));
 AOI21x1_ASAP7_75t_SL _19485_ (.A1(_11270_),
    .A2(_11273_),
    .B(_10821_),
    .Y(_11274_));
 AOI21x1_ASAP7_75t_SL _19486_ (.A1(_11269_),
    .A2(_11274_),
    .B(_10920_),
    .Y(_11275_));
 OAI21x1_ASAP7_75t_SL _19487_ (.A1(_11256_),
    .A2(_11262_),
    .B(_11275_),
    .Y(_11276_));
 NAND2x1_ASAP7_75t_SL _19488_ (.A(_11250_),
    .B(_11276_),
    .Y(_00037_));
 INVx1_ASAP7_75t_SL _19489_ (.A(_10807_),
    .Y(_11277_));
 AOI21x1_ASAP7_75t_SL _19490_ (.A1(_11277_),
    .A2(_11189_),
    .B(_10875_),
    .Y(_11278_));
 OR4x1_ASAP7_75t_SL _19491_ (.A(_11028_),
    .B(_10962_),
    .C(_10810_),
    .D(_10774_),
    .Y(_11279_));
 NAND2x1_ASAP7_75t_SL _19492_ (.A(_11278_),
    .B(_11279_),
    .Y(_11280_));
 AO21x1_ASAP7_75t_SL _19493_ (.A1(_11143_),
    .A2(_11029_),
    .B(_10778_),
    .Y(_11281_));
 OA21x2_ASAP7_75t_SL _19494_ (.A1(_10841_),
    .A2(_10770_),
    .B(_10810_),
    .Y(_11282_));
 AOI21x1_ASAP7_75t_SL _19495_ (.A1(_11281_),
    .A2(_11282_),
    .B(_10835_),
    .Y(_11283_));
 AO21x1_ASAP7_75t_SL _19496_ (.A1(_10770_),
    .A2(_01074_),
    .B(_10810_),
    .Y(_11284_));
 AO21x1_ASAP7_75t_SL _19497_ (.A1(_10971_),
    .A2(_11039_),
    .B(_11284_),
    .Y(_11285_));
 AOI21x1_ASAP7_75t_SL _19498_ (.A1(_11283_),
    .A2(_11285_),
    .B(_10821_),
    .Y(_11286_));
 NAND2x1_ASAP7_75t_SL _19499_ (.A(_11280_),
    .B(_11286_),
    .Y(_11287_));
 OA21x2_ASAP7_75t_SL _19500_ (.A1(_11067_),
    .A2(_11200_),
    .B(_10841_),
    .Y(_11288_));
 NOR2x1_ASAP7_75t_SL _19501_ (.A(_10755_),
    .B(_11288_),
    .Y(_11289_));
 NAND2x1_ASAP7_75t_SL _19502_ (.A(_10778_),
    .B(_01061_),
    .Y(_11290_));
 AO21x1_ASAP7_75t_SL _19503_ (.A1(_11135_),
    .A2(_11290_),
    .B(_10835_),
    .Y(_11291_));
 NOR2x1_ASAP7_75t_SL _19504_ (.A(_10755_),
    .B(_10963_),
    .Y(_11292_));
 NAND2x1_ASAP7_75t_SL _19505_ (.A(_10891_),
    .B(_11292_),
    .Y(_11293_));
 NAND2x1_ASAP7_75t_SL _19506_ (.A(_11055_),
    .B(_11035_),
    .Y(_11294_));
 AOI21x1_ASAP7_75t_SL _19507_ (.A1(_11294_),
    .A2(_11240_),
    .B(_10875_),
    .Y(_11295_));
 AOI21x1_ASAP7_75t_SL _19508_ (.A1(_11293_),
    .A2(_11295_),
    .B(_10742_),
    .Y(_11296_));
 OAI21x1_ASAP7_75t_SL _19509_ (.A1(_11289_),
    .A2(_11291_),
    .B(_11296_),
    .Y(_11297_));
 AOI21x1_ASAP7_75t_SL _19510_ (.A1(_11287_),
    .A2(_11297_),
    .B(_10920_),
    .Y(_11298_));
 NAND2x1_ASAP7_75t_SL _19511_ (.A(_10908_),
    .B(_11039_),
    .Y(_11299_));
 AOI21x1_ASAP7_75t_SL _19512_ (.A1(_11299_),
    .A2(_11096_),
    .B(_10810_),
    .Y(_11300_));
 NAND2x1_ASAP7_75t_R _19513_ (.A(_10871_),
    .B(_10852_),
    .Y(_11301_));
 NOR2x1_ASAP7_75t_SL _19514_ (.A(_11028_),
    .B(_11301_),
    .Y(_11302_));
 NAND2x1_ASAP7_75t_SL _19515_ (.A(_11251_),
    .B(_10861_),
    .Y(_11303_));
 OAI21x1_ASAP7_75t_SL _19516_ (.A1(_11302_),
    .A2(_11303_),
    .B(_10835_),
    .Y(_11304_));
 NOR2x1_ASAP7_75t_SL _19517_ (.A(_11300_),
    .B(_11304_),
    .Y(_11305_));
 OAI21x1_ASAP7_75t_SL _19518_ (.A1(_10770_),
    .A2(_10869_),
    .B(_10810_),
    .Y(_11306_));
 AOI21x1_ASAP7_75t_SL _19519_ (.A1(_10871_),
    .A2(_10852_),
    .B(_10778_),
    .Y(_11307_));
 NOR2x1_ASAP7_75t_SL _19520_ (.A(_11306_),
    .B(_11307_),
    .Y(_11308_));
 AND2x2_ASAP7_75t_R _19521_ (.A(_01079_),
    .B(_01073_),
    .Y(_11309_));
 OAI21x1_ASAP7_75t_SL _19522_ (.A1(_11309_),
    .A2(_10770_),
    .B(_10755_),
    .Y(_11310_));
 AOI21x1_ASAP7_75t_SL _19523_ (.A1(_10803_),
    .A2(_11076_),
    .B(_11310_),
    .Y(_11311_));
 OAI21x1_ASAP7_75t_SL _19524_ (.A1(_11308_),
    .A2(_11311_),
    .B(_10875_),
    .Y(_11312_));
 NAND2x1_ASAP7_75t_SL _19525_ (.A(_10821_),
    .B(_11312_),
    .Y(_11313_));
 OAI21x1_ASAP7_75t_SL _19526_ (.A1(_11305_),
    .A2(_11313_),
    .B(_10920_),
    .Y(_11314_));
 AO21x1_ASAP7_75t_SL _19527_ (.A1(_11143_),
    .A2(_10871_),
    .B(_10770_),
    .Y(_11315_));
 NOR2x1_ASAP7_75t_SL _19528_ (.A(_10778_),
    .B(_10962_),
    .Y(_11316_));
 NAND2x1_ASAP7_75t_SL _19529_ (.A(_10899_),
    .B(_11316_),
    .Y(_11317_));
 AOI21x1_ASAP7_75t_SL _19530_ (.A1(_11315_),
    .A2(_11317_),
    .B(_10810_),
    .Y(_11318_));
 AO21x1_ASAP7_75t_SL _19531_ (.A1(_10778_),
    .A2(_10850_),
    .B(_10755_),
    .Y(_11319_));
 OAI21x1_ASAP7_75t_SL _19532_ (.A1(_11319_),
    .A2(_11089_),
    .B(_10875_),
    .Y(_11320_));
 OAI21x1_ASAP7_75t_SL _19533_ (.A1(_11318_),
    .A2(_11320_),
    .B(_10742_),
    .Y(_11321_));
 AO21x1_ASAP7_75t_SL _19534_ (.A1(_11142_),
    .A2(_10778_),
    .B(_10755_),
    .Y(_11322_));
 AO21x1_ASAP7_75t_SL _19535_ (.A1(_10803_),
    .A2(_10963_),
    .B(_11322_),
    .Y(_11323_));
 AND3x1_ASAP7_75t_SL _19536_ (.A(_10770_),
    .B(_10723_),
    .C(_10721_),
    .Y(_11324_));
 AOI21x1_ASAP7_75t_SL _19537_ (.A1(_10987_),
    .A2(_11112_),
    .B(_11324_),
    .Y(_11325_));
 NAND2x1_ASAP7_75t_SL _19538_ (.A(_11186_),
    .B(_11325_),
    .Y(_11326_));
 AOI21x1_ASAP7_75t_SL _19539_ (.A1(_11323_),
    .A2(_11326_),
    .B(_10875_),
    .Y(_11327_));
 NOR2x1_ASAP7_75t_SL _19540_ (.A(_11321_),
    .B(_11327_),
    .Y(_11328_));
 NOR2x1_ASAP7_75t_SL _19541_ (.A(_11314_),
    .B(_11328_),
    .Y(_11329_));
 NOR2x1_ASAP7_75t_SL _19542_ (.A(_11298_),
    .B(_11329_),
    .Y(_00038_));
 OAI21x1_ASAP7_75t_SL _19543_ (.A1(_10770_),
    .A2(_10687_),
    .B(_10810_),
    .Y(_11330_));
 AOI21x1_ASAP7_75t_SL _19544_ (.A1(_10721_),
    .A2(_11266_),
    .B(_11330_),
    .Y(_11331_));
 AO21x1_ASAP7_75t_SL _19545_ (.A1(_11331_),
    .A2(_11113_),
    .B(_10835_),
    .Y(_11332_));
 NOR2x1_ASAP7_75t_SL _19546_ (.A(_11156_),
    .B(_10976_),
    .Y(_11333_));
 AOI22x1_ASAP7_75t_SL _19547_ (.A1(_10851_),
    .A2(_10777_),
    .B1(_11333_),
    .B2(_10778_),
    .Y(_11334_));
 NOR2x1_ASAP7_75t_SL _19548_ (.A(_10810_),
    .B(_11334_),
    .Y(_11335_));
 NOR2x1_ASAP7_75t_SL _19549_ (.A(_11332_),
    .B(_11335_),
    .Y(_11336_));
 INVx1_ASAP7_75t_SL _19550_ (.A(_10872_),
    .Y(_11337_));
 AOI21x1_ASAP7_75t_SL _19551_ (.A1(_10770_),
    .A2(_10915_),
    .B(_11156_),
    .Y(_11338_));
 AOI21x1_ASAP7_75t_SL _19552_ (.A1(_11337_),
    .A2(_11338_),
    .B(_10875_),
    .Y(_11339_));
 AO21x1_ASAP7_75t_SL _19553_ (.A1(_10778_),
    .A2(_10783_),
    .B(_10755_),
    .Y(_11340_));
 AO21x1_ASAP7_75t_SL _19554_ (.A1(_11076_),
    .A2(_10803_),
    .B(_11340_),
    .Y(_11341_));
 AO21x1_ASAP7_75t_SL _19555_ (.A1(_11339_),
    .A2(_11341_),
    .B(_10742_),
    .Y(_11342_));
 INVx1_ASAP7_75t_SL _19556_ (.A(_10997_),
    .Y(_11343_));
 AO21x1_ASAP7_75t_SL _19557_ (.A1(_10778_),
    .A2(_10774_),
    .B(_11330_),
    .Y(_11344_));
 AND2x2_ASAP7_75t_SL _19558_ (.A(_10770_),
    .B(_01070_),
    .Y(_11345_));
 OA21x2_ASAP7_75t_SL _19559_ (.A1(_10872_),
    .A2(_11345_),
    .B(_10875_),
    .Y(_11346_));
 OAI21x1_ASAP7_75t_SL _19560_ (.A1(_11343_),
    .A2(_11344_),
    .B(_11346_),
    .Y(_11347_));
 NAND2x1_ASAP7_75t_SL _19561_ (.A(_10778_),
    .B(_10928_),
    .Y(_11348_));
 OAI21x1_ASAP7_75t_SL _19562_ (.A1(_01079_),
    .A2(_10778_),
    .B(_10755_),
    .Y(_11349_));
 NOR2x1_ASAP7_75t_SL _19563_ (.A(_11349_),
    .B(_10854_),
    .Y(_11350_));
 AOI21x1_ASAP7_75t_SL _19564_ (.A1(_11348_),
    .A2(_11350_),
    .B(_10875_),
    .Y(_11351_));
 NAND2x1_ASAP7_75t_SL _19565_ (.A(_10971_),
    .B(_10903_),
    .Y(_11352_));
 AOI21x1_ASAP7_75t_SL _19566_ (.A1(_10922_),
    .A2(_10929_),
    .B(_10755_),
    .Y(_11353_));
 NAND2x1_ASAP7_75t_SL _19567_ (.A(_11352_),
    .B(_11353_),
    .Y(_11354_));
 AOI21x1_ASAP7_75t_SL _19568_ (.A1(_11351_),
    .A2(_11354_),
    .B(_10821_),
    .Y(_11355_));
 AOI21x1_ASAP7_75t_SL _19569_ (.A1(_11347_),
    .A2(_11355_),
    .B(_10887_),
    .Y(_11356_));
 OAI21x1_ASAP7_75t_SL _19570_ (.A1(_11336_),
    .A2(_11342_),
    .B(_11356_),
    .Y(_11357_));
 NAND2x1_ASAP7_75t_SL _19571_ (.A(_10819_),
    .B(_10971_),
    .Y(_11358_));
 NOR2x1_ASAP7_75t_SL _19572_ (.A(_10810_),
    .B(_11200_),
    .Y(_11359_));
 AOI21x1_ASAP7_75t_SL _19573_ (.A1(_11358_),
    .A2(_11359_),
    .B(_10835_),
    .Y(_11360_));
 OAI21x1_ASAP7_75t_SL _19574_ (.A1(_10721_),
    .A2(_10687_),
    .B(_10723_),
    .Y(_11361_));
 AOI21x1_ASAP7_75t_SL _19575_ (.A1(_10778_),
    .A2(_11361_),
    .B(_10755_),
    .Y(_11362_));
 OAI21x1_ASAP7_75t_SL _19576_ (.A1(_10778_),
    .A2(_11333_),
    .B(_11362_),
    .Y(_11363_));
 AOI21x1_ASAP7_75t_SL _19577_ (.A1(_11360_),
    .A2(_11363_),
    .B(_10742_),
    .Y(_11364_));
 AO21x1_ASAP7_75t_SL _19578_ (.A1(_11001_),
    .A2(_10758_),
    .B(_10778_),
    .Y(_11365_));
 AOI21x1_ASAP7_75t_SL _19579_ (.A1(_11365_),
    .A2(_11121_),
    .B(_10755_),
    .Y(_11366_));
 AOI21x1_ASAP7_75t_SL _19580_ (.A1(_11299_),
    .A2(_11077_),
    .B(_10810_),
    .Y(_11367_));
 OAI21x1_ASAP7_75t_SL _19581_ (.A1(_11366_),
    .A2(_11367_),
    .B(_10835_),
    .Y(_11368_));
 AOI21x1_ASAP7_75t_SL _19582_ (.A1(_11364_),
    .A2(_11368_),
    .B(_10920_),
    .Y(_11369_));
 OAI21x1_ASAP7_75t_SL _19583_ (.A1(_10728_),
    .A2(_10942_),
    .B(_10912_),
    .Y(_11370_));
 NAND2x1_ASAP7_75t_SL _19584_ (.A(_11068_),
    .B(_11370_),
    .Y(_11371_));
 AO21x1_ASAP7_75t_SL _19585_ (.A1(_10963_),
    .A2(_10984_),
    .B(_11266_),
    .Y(_11372_));
 AOI21x1_ASAP7_75t_SL _19586_ (.A1(_10810_),
    .A2(_11372_),
    .B(_10835_),
    .Y(_11373_));
 NAND2x1_ASAP7_75t_SL _19587_ (.A(_11371_),
    .B(_11373_),
    .Y(_11374_));
 AND2x2_ASAP7_75t_SL _19588_ (.A(_11097_),
    .B(_10942_),
    .Y(_11375_));
 NAND2x1_ASAP7_75t_SL _19589_ (.A(_10755_),
    .B(_11127_),
    .Y(_11376_));
 OA21x2_ASAP7_75t_SL _19590_ (.A1(_11375_),
    .A2(_11376_),
    .B(_10835_),
    .Y(_11377_));
 AO21x1_ASAP7_75t_SL _19591_ (.A1(_11208_),
    .A2(_01067_),
    .B(_11055_),
    .Y(_11378_));
 AOI21x1_ASAP7_75t_SL _19592_ (.A1(_10770_),
    .A2(_10805_),
    .B(_10755_),
    .Y(_11379_));
 NAND2x1_ASAP7_75t_SL _19593_ (.A(_11378_),
    .B(_11379_),
    .Y(_11380_));
 AOI21x1_ASAP7_75t_SL _19594_ (.A1(_11377_),
    .A2(_11380_),
    .B(_10821_),
    .Y(_11381_));
 NAND2x1_ASAP7_75t_SL _19595_ (.A(_11374_),
    .B(_11381_),
    .Y(_11382_));
 NAND2x1_ASAP7_75t_SL _19596_ (.A(_11369_),
    .B(_11382_),
    .Y(_11383_));
 NAND2x1_ASAP7_75t_SL _19597_ (.A(_11357_),
    .B(_11383_),
    .Y(_00039_));
 NOR2x1_ASAP7_75t_R _19599_ (.A(_00574_),
    .B(_00447_),
    .Y(_11385_));
 XOR2x2_ASAP7_75t_SL _19600_ (.A(_00622_),
    .B(_00615_),
    .Y(_11386_));
 XOR2x2_ASAP7_75t_SL _19601_ (.A(_00680_),
    .B(_11386_),
    .Y(_11387_));
 XOR2x2_ASAP7_75t_SL _19602_ (.A(_00590_),
    .B(_00583_),
    .Y(_11388_));
 XOR2x2_ASAP7_75t_SL _19603_ (.A(_00648_),
    .B(_00616_),
    .Y(_11389_));
 XOR2x2_ASAP7_75t_SL _19604_ (.A(_11389_),
    .B(_11388_),
    .Y(_11390_));
 NAND2x1p5_ASAP7_75t_SL _19605_ (.A(_11387_),
    .B(_11390_),
    .Y(_11391_));
 INVx1_ASAP7_75t_R _19606_ (.A(_00680_),
    .Y(_11392_));
 XOR2x2_ASAP7_75t_SL _19607_ (.A(_11392_),
    .B(_11386_),
    .Y(_11393_));
 XNOR2x2_ASAP7_75t_SL _19608_ (.A(_00590_),
    .B(_00583_),
    .Y(_11394_));
 XOR2x2_ASAP7_75t_SL _19609_ (.A(_11389_),
    .B(_11394_),
    .Y(_11395_));
 NAND2x1p5_ASAP7_75t_SL _19610_ (.A(_11393_),
    .B(_11395_),
    .Y(_11396_));
 AOI21x1_ASAP7_75t_SL _19613_ (.A1(_11396_),
    .A2(_11391_),
    .B(_10675_),
    .Y(_11399_));
 OAI21x1_ASAP7_75t_SL _19614_ (.A1(_11399_),
    .A2(_11385_),
    .B(_00887_),
    .Y(_11400_));
 AND2x2_ASAP7_75t_R _19615_ (.A(_10675_),
    .B(_00447_),
    .Y(_11401_));
 NAND2x1p5_ASAP7_75t_SL _19616_ (.A(_11393_),
    .B(_11390_),
    .Y(_11402_));
 NAND2x1p5_ASAP7_75t_SL _19617_ (.A(_11387_),
    .B(_11395_),
    .Y(_11403_));
 AOI21x1_ASAP7_75t_SL _19619_ (.A1(_11403_),
    .A2(_11402_),
    .B(_10675_),
    .Y(_11405_));
 OAI21x1_ASAP7_75t_SL _19620_ (.A1(_11405_),
    .A2(_11401_),
    .B(_08768_),
    .Y(_11406_));
 NAND2x2_ASAP7_75t_SL _19621_ (.A(_11406_),
    .B(_11400_),
    .Y(_11407_));
 INVx1_ASAP7_75t_R _19623_ (.A(_00679_),
    .Y(_11408_));
 XOR2x2_ASAP7_75t_SL _19624_ (.A(_00622_),
    .B(_00590_),
    .Y(_11409_));
 NAND2x1_ASAP7_75t_R _19625_ (.A(_11408_),
    .B(_11409_),
    .Y(_11410_));
 XNOR2x2_ASAP7_75t_L _19626_ (.A(_00590_),
    .B(_00622_),
    .Y(_11411_));
 NAND2x1_ASAP7_75t_L _19627_ (.A(_00679_),
    .B(_11411_),
    .Y(_11412_));
 XNOR2x2_ASAP7_75t_L _19628_ (.A(_00647_),
    .B(_00615_),
    .Y(_11413_));
 AOI21x1_ASAP7_75t_R _19629_ (.A1(_11410_),
    .A2(_11412_),
    .B(_11413_),
    .Y(_11414_));
 NAND2x1_ASAP7_75t_R _19630_ (.A(_00679_),
    .B(_11409_),
    .Y(_11415_));
 NAND2x1_ASAP7_75t_L _19631_ (.A(_11408_),
    .B(_11411_),
    .Y(_11416_));
 XOR2x2_ASAP7_75t_SL _19632_ (.A(_00647_),
    .B(_00615_),
    .Y(_11417_));
 AOI21x1_ASAP7_75t_R _19633_ (.A1(_11415_),
    .A2(_11416_),
    .B(_11417_),
    .Y(_11418_));
 OAI21x1_ASAP7_75t_SL _19634_ (.A1(_11418_),
    .A2(_11414_),
    .B(_00574_),
    .Y(_11419_));
 NOR2x1_ASAP7_75t_L _19635_ (.A(_00574_),
    .B(_00448_),
    .Y(_11420_));
 INVx1_ASAP7_75t_R _19636_ (.A(_11420_),
    .Y(_11421_));
 NAND3x1_ASAP7_75t_R _19637_ (.A(_11419_),
    .B(_10106_),
    .C(_11421_),
    .Y(_11422_));
 INVx2_ASAP7_75t_SL _19638_ (.A(_11419_),
    .Y(_11423_));
 OAI21x1_ASAP7_75t_R _19639_ (.A1(_11420_),
    .A2(_11423_),
    .B(_00886_),
    .Y(_11424_));
 NAND2x2_ASAP7_75t_SL _19640_ (.A(_11424_),
    .B(_11422_),
    .Y(_01088_));
 NOR2x1_ASAP7_75t_SL _19641_ (.A(_00574_),
    .B(_00449_),
    .Y(_11425_));
 XOR2x2_ASAP7_75t_SL _19642_ (.A(_00616_),
    .B(_00584_),
    .Y(_11426_));
 NOR2x1_ASAP7_75t_R _19643_ (.A(_00617_),
    .B(_11426_),
    .Y(_11427_));
 NAND2x1_ASAP7_75t_SL _19644_ (.A(_00617_),
    .B(_11426_),
    .Y(_11428_));
 INVx1_ASAP7_75t_R _19645_ (.A(_11428_),
    .Y(_11429_));
 XNOR2x1_ASAP7_75t_SL _19646_ (.B(_00681_),
    .Y(_11430_),
    .A(_00649_));
 OAI21x1_ASAP7_75t_SL _19647_ (.A1(_11427_),
    .A2(_11429_),
    .B(_11430_),
    .Y(_11431_));
 INVx1_ASAP7_75t_R _19648_ (.A(_00617_),
    .Y(_11432_));
 NAND2x1_ASAP7_75t_SL _19649_ (.A(_11432_),
    .B(_11426_),
    .Y(_11433_));
 XNOR2x2_ASAP7_75t_SL _19650_ (.A(_00616_),
    .B(_00584_),
    .Y(_11434_));
 NAND2x1_ASAP7_75t_R _19651_ (.A(_00617_),
    .B(_11434_),
    .Y(_11435_));
 AOI21x1_ASAP7_75t_SL _19652_ (.A1(_11433_),
    .A2(_11435_),
    .B(_11430_),
    .Y(_11436_));
 INVx1_ASAP7_75t_SL _19653_ (.A(_11436_),
    .Y(_11437_));
 AOI21x1_ASAP7_75t_SL _19654_ (.A1(_11431_),
    .A2(_11437_),
    .B(_10675_),
    .Y(_11438_));
 OAI21x1_ASAP7_75t_R _19655_ (.A1(_11425_),
    .A2(_11438_),
    .B(_08953_),
    .Y(_11439_));
 NAND2x1_ASAP7_75t_R _19656_ (.A(_11432_),
    .B(_11434_),
    .Y(_11440_));
 XOR2x1_ASAP7_75t_SL _19657_ (.A(_00649_),
    .Y(_11441_),
    .B(_00681_));
 AOI21x1_ASAP7_75t_R _19658_ (.A1(_11428_),
    .A2(_11440_),
    .B(_11441_),
    .Y(_11442_));
 OAI21x1_ASAP7_75t_SL _19659_ (.A1(_11436_),
    .A2(_11442_),
    .B(_00574_),
    .Y(_11443_));
 INVx1_ASAP7_75t_SL _19660_ (.A(_11425_),
    .Y(_11444_));
 NAND3x1_ASAP7_75t_SL _19661_ (.A(_11443_),
    .B(_00888_),
    .C(_11444_),
    .Y(_11445_));
 NAND2x2_ASAP7_75t_SL _19662_ (.A(_11439_),
    .B(_11445_),
    .Y(_11446_));
 NAND3x1_ASAP7_75t_L _19664_ (.A(_11419_),
    .B(_00886_),
    .C(_11421_),
    .Y(_11447_));
 OAI21x1_ASAP7_75t_SL _19665_ (.A1(_11423_),
    .A2(_11420_),
    .B(_10106_),
    .Y(_11448_));
 NAND2x2_ASAP7_75t_SL _19666_ (.A(_11448_),
    .B(_11447_),
    .Y(_11449_));
 OAI21x1_ASAP7_75t_SL _19668_ (.A1(_11425_),
    .A2(_11438_),
    .B(_00888_),
    .Y(_11450_));
 NAND3x1_ASAP7_75t_SL _19669_ (.A(_11443_),
    .B(_08953_),
    .C(_11444_),
    .Y(_11451_));
 NAND2x2_ASAP7_75t_SL _19670_ (.A(_11450_),
    .B(_11451_),
    .Y(_11452_));
 XOR2x2_ASAP7_75t_L _19673_ (.A(_00617_),
    .B(_00622_),
    .Y(_11454_));
 XOR2x2_ASAP7_75t_R _19674_ (.A(_00650_),
    .B(_00682_),
    .Y(_11455_));
 XOR2x2_ASAP7_75t_L _19675_ (.A(_11454_),
    .B(_11455_),
    .Y(_11456_));
 XOR2x2_ASAP7_75t_SL _19676_ (.A(_00585_),
    .B(_00590_),
    .Y(_11457_));
 XOR2x2_ASAP7_75t_R _19677_ (.A(_11457_),
    .B(_00618_),
    .Y(_11458_));
 AND2x2_ASAP7_75t_SL _19678_ (.A(_11456_),
    .B(_11458_),
    .Y(_11459_));
 OAI21x1_ASAP7_75t_R _19679_ (.A1(_11458_),
    .A2(_11456_),
    .B(_00574_),
    .Y(_11460_));
 NAND2x1_ASAP7_75t_R _19680_ (.A(_00494_),
    .B(_10675_),
    .Y(_11461_));
 OAI21x1_ASAP7_75t_SL _19681_ (.A1(_11459_),
    .A2(_11460_),
    .B(_11461_),
    .Y(_11462_));
 XOR2x2_ASAP7_75t_SL _19682_ (.A(_11462_),
    .B(_08963_),
    .Y(_11463_));
 INVx4_ASAP7_75t_SL _19684_ (.A(_11407_),
    .Y(_01082_));
 NAND2x1_ASAP7_75t_R _19685_ (.A(_11463_),
    .B(_01082_),
    .Y(_11465_));
 OAI21x1_ASAP7_75t_SL _19686_ (.A1(_11452_),
    .A2(_01088_),
    .B(_11463_),
    .Y(_11466_));
 NAND2x1_ASAP7_75t_SL _19687_ (.A(_11452_),
    .B(_11449_),
    .Y(_11467_));
 INVx1_ASAP7_75t_R _19688_ (.A(_11467_),
    .Y(_11468_));
 AO21x1_ASAP7_75t_SL _19689_ (.A1(_11465_),
    .A2(_11466_),
    .B(_11468_),
    .Y(_11469_));
 XOR2x2_ASAP7_75t_SL _19690_ (.A(_11462_),
    .B(_00889_),
    .Y(_11470_));
 INVx1_ASAP7_75t_SL _19695_ (.A(_01092_),
    .Y(_11475_));
 AO21x1_ASAP7_75t_SL _19696_ (.A1(_11445_),
    .A2(_11439_),
    .B(_11475_),
    .Y(_11476_));
 NAND2x1_ASAP7_75t_SL _19697_ (.A(_11470_),
    .B(_11476_),
    .Y(_11477_));
 INVx1_ASAP7_75t_SL _19698_ (.A(_01084_),
    .Y(_11478_));
 AOI21x1_ASAP7_75t_SL _19699_ (.A1(_11450_),
    .A2(_11451_),
    .B(_11478_),
    .Y(_11479_));
 XOR2x2_ASAP7_75t_R _19701_ (.A(_00618_),
    .B(_00622_),
    .Y(_11481_));
 XOR2x2_ASAP7_75t_R _19702_ (.A(_00651_),
    .B(_00683_),
    .Y(_11482_));
 XOR2x2_ASAP7_75t_SL _19703_ (.A(_11481_),
    .B(_11482_),
    .Y(_11483_));
 XOR2x2_ASAP7_75t_SL _19704_ (.A(_00586_),
    .B(_00590_),
    .Y(_11484_));
 XNOR2x2_ASAP7_75t_R _19705_ (.A(_00619_),
    .B(_11484_),
    .Y(_11485_));
 XOR2x2_ASAP7_75t_SL _19706_ (.A(_11483_),
    .B(_11485_),
    .Y(_11486_));
 NOR2x1_ASAP7_75t_R _19707_ (.A(_00574_),
    .B(_00493_),
    .Y(_11487_));
 AOI21x1_ASAP7_75t_SL _19708_ (.A1(_00574_),
    .A2(_11486_),
    .B(_11487_),
    .Y(_11488_));
 XOR2x2_ASAP7_75t_SL _19709_ (.A(_11488_),
    .B(_00890_),
    .Y(_11489_));
 OA21x2_ASAP7_75t_R _19712_ (.A1(_11477_),
    .A2(_11479_),
    .B(_11489_),
    .Y(_11492_));
 XOR2x2_ASAP7_75t_SL _19713_ (.A(_11488_),
    .B(_08775_),
    .Y(_11493_));
 NAND2x1_ASAP7_75t_R _19715_ (.A(_11493_),
    .B(_11466_),
    .Y(_11495_));
 AOI21x1_ASAP7_75t_SL _19717_ (.A1(_01087_),
    .A2(_11452_),
    .B(_11463_),
    .Y(_11497_));
 INVx1_ASAP7_75t_L _19718_ (.A(_11497_),
    .Y(_11498_));
 NAND2x1_ASAP7_75t_SL _19719_ (.A(_11449_),
    .B(_11407_),
    .Y(_11499_));
 NOR2x1_ASAP7_75t_SL _19721_ (.A(_11452_),
    .B(_11499_),
    .Y(_11501_));
 NOR2x1_ASAP7_75t_SL _19722_ (.A(_11498_),
    .B(_11501_),
    .Y(_11502_));
 XOR2x2_ASAP7_75t_SL _19723_ (.A(_00588_),
    .B(_00620_),
    .Y(_11503_));
 XOR2x2_ASAP7_75t_R _19724_ (.A(_00621_),
    .B(_00653_),
    .Y(_11504_));
 XOR2x2_ASAP7_75t_R _19725_ (.A(_11504_),
    .B(_00685_),
    .Y(_11505_));
 XNOR2x2_ASAP7_75t_R _19726_ (.A(_11503_),
    .B(_11505_),
    .Y(_11506_));
 NOR2x1_ASAP7_75t_R _19730_ (.A(_00574_),
    .B(_00491_),
    .Y(_11510_));
 AO21x1_ASAP7_75t_SL _19731_ (.A1(_11506_),
    .A2(_00574_),
    .B(_11510_),
    .Y(_11511_));
 XOR2x2_ASAP7_75t_SL _19732_ (.A(_11511_),
    .B(_00893_),
    .Y(_11512_));
 INVx2_ASAP7_75t_SL _19733_ (.A(_11512_),
    .Y(_11513_));
 OAI21x1_ASAP7_75t_R _19735_ (.A1(_11495_),
    .A2(_11502_),
    .B(_11513_),
    .Y(_11515_));
 AOI21x1_ASAP7_75t_R _19736_ (.A1(_11469_),
    .A2(_11492_),
    .B(_11515_),
    .Y(_11516_));
 AOI21x1_ASAP7_75t_SL _19737_ (.A1(_01088_),
    .A2(_11407_),
    .B(_11452_),
    .Y(_11517_));
 INVx1_ASAP7_75t_SL _19738_ (.A(_11517_),
    .Y(_11518_));
 AO21x2_ASAP7_75t_SL _19739_ (.A1(_11451_),
    .A2(_11450_),
    .B(_01084_),
    .Y(_11519_));
 AO21x1_ASAP7_75t_R _19741_ (.A1(_11518_),
    .A2(_11519_),
    .B(_11470_),
    .Y(_11521_));
 INVx1_ASAP7_75t_R _19742_ (.A(_01083_),
    .Y(_11522_));
 AO21x1_ASAP7_75t_R _19743_ (.A1(_11445_),
    .A2(_11439_),
    .B(_11522_),
    .Y(_11523_));
 INVx1_ASAP7_75t_SL _19745_ (.A(_01089_),
    .Y(_11525_));
 AO21x1_ASAP7_75t_SL _19746_ (.A1(_11451_),
    .A2(_11450_),
    .B(_11525_),
    .Y(_11526_));
 AOI21x1_ASAP7_75t_R _19748_ (.A1(_11523_),
    .A2(_11526_),
    .B(_11463_),
    .Y(_11528_));
 NOR2x1_ASAP7_75t_R _19749_ (.A(_11489_),
    .B(_11528_),
    .Y(_11529_));
 NAND2x1_ASAP7_75t_SL _19750_ (.A(_11449_),
    .B(_01082_),
    .Y(_11530_));
 NOR2x1_ASAP7_75t_SL _19751_ (.A(_11446_),
    .B(_11449_),
    .Y(_11531_));
 NOR2x1_ASAP7_75t_SL _19752_ (.A(_11470_),
    .B(_11531_),
    .Y(_11532_));
 NAND2x1_ASAP7_75t_SL _19753_ (.A(_11530_),
    .B(_11532_),
    .Y(_11533_));
 INVx1_ASAP7_75t_SL _19754_ (.A(_11533_),
    .Y(_11534_));
 NAND2x2_ASAP7_75t_SL _19757_ (.A(_11446_),
    .B(_01088_),
    .Y(_11537_));
 NAND2x1_ASAP7_75t_SL _19758_ (.A(_11537_),
    .B(_11499_),
    .Y(_11538_));
 OAI21x1_ASAP7_75t_SL _19759_ (.A1(_11463_),
    .A2(_11538_),
    .B(_11489_),
    .Y(_11539_));
 OAI21x1_ASAP7_75t_R _19761_ (.A1(_11534_),
    .A2(_11539_),
    .B(_11512_),
    .Y(_11541_));
 AOI21x1_ASAP7_75t_R _19762_ (.A1(_11521_),
    .A2(_11529_),
    .B(_11541_),
    .Y(_11542_));
 XOR2x2_ASAP7_75t_SL _19763_ (.A(_00620_),
    .B(_00652_),
    .Y(_11543_));
 XOR2x2_ASAP7_75t_R _19764_ (.A(_11543_),
    .B(_00684_),
    .Y(_11544_));
 XNOR2x2_ASAP7_75t_R _19765_ (.A(_00587_),
    .B(_00619_),
    .Y(_11545_));
 XOR2x2_ASAP7_75t_L _19766_ (.A(_11544_),
    .B(_11545_),
    .Y(_11546_));
 NAND2x1_ASAP7_75t_R _19767_ (.A(_00574_),
    .B(_11546_),
    .Y(_11547_));
 OA21x2_ASAP7_75t_SL _19768_ (.A1(_00574_),
    .A2(_00492_),
    .B(_11547_),
    .Y(_11548_));
 XOR2x2_ASAP7_75t_SL _19769_ (.A(_11548_),
    .B(_00891_),
    .Y(_11549_));
 OAI21x1_ASAP7_75t_R _19771_ (.A1(_11516_),
    .A2(_11542_),
    .B(_11549_),
    .Y(_11551_));
 NAND2x2_ASAP7_75t_SL _19772_ (.A(_11446_),
    .B(_11407_),
    .Y(_11552_));
 OA21x2_ASAP7_75t_SL _19773_ (.A1(_11446_),
    .A2(_01084_),
    .B(_11463_),
    .Y(_11553_));
 NAND2x1_ASAP7_75t_R _19774_ (.A(_11552_),
    .B(_11553_),
    .Y(_11554_));
 OA21x2_ASAP7_75t_SL _19777_ (.A1(_11452_),
    .A2(_11478_),
    .B(_11470_),
    .Y(_11557_));
 NOR2x1_ASAP7_75t_SL _19778_ (.A(_11493_),
    .B(_11557_),
    .Y(_11558_));
 AOI21x1_ASAP7_75t_R _19779_ (.A1(_11554_),
    .A2(_11558_),
    .B(_11513_),
    .Y(_11559_));
 AO21x1_ASAP7_75t_R _19781_ (.A1(_11519_),
    .A2(_11523_),
    .B(_11463_),
    .Y(_11561_));
 AO21x1_ASAP7_75t_SL _19782_ (.A1(_11445_),
    .A2(_11439_),
    .B(_11525_),
    .Y(_11562_));
 AO21x1_ASAP7_75t_R _19783_ (.A1(_11451_),
    .A2(_11450_),
    .B(_11522_),
    .Y(_11563_));
 AO21x1_ASAP7_75t_R _19785_ (.A1(_11562_),
    .A2(_11563_),
    .B(_11470_),
    .Y(_11565_));
 AO21x1_ASAP7_75t_R _19786_ (.A1(_11561_),
    .A2(_11565_),
    .B(_11489_),
    .Y(_11566_));
 AOI21x1_ASAP7_75t_R _19787_ (.A1(_11559_),
    .A2(_11566_),
    .B(_11549_),
    .Y(_11567_));
 AO21x1_ASAP7_75t_R _19788_ (.A1(_11451_),
    .A2(_11450_),
    .B(_01085_),
    .Y(_11568_));
 INVx1_ASAP7_75t_SL _19789_ (.A(_11568_),
    .Y(_11569_));
 NOR2x2_ASAP7_75t_SL _19790_ (.A(_11452_),
    .B(_11407_),
    .Y(_11570_));
 OA21x2_ASAP7_75t_R _19791_ (.A1(_11569_),
    .A2(_11570_),
    .B(_11463_),
    .Y(_11571_));
 NAND2x1_ASAP7_75t_SL _19792_ (.A(_11446_),
    .B(_11449_),
    .Y(_11572_));
 INVx1_ASAP7_75t_SL _19793_ (.A(_11572_),
    .Y(_11573_));
 NAND2x2_ASAP7_75t_SL _19794_ (.A(_01088_),
    .B(_11407_),
    .Y(_11574_));
 OAI21x1_ASAP7_75t_SL _19796_ (.A1(_11446_),
    .A2(_11574_),
    .B(_11470_),
    .Y(_11576_));
 NOR2x1_ASAP7_75t_SL _19797_ (.A(_11573_),
    .B(_11576_),
    .Y(_11577_));
 OAI21x1_ASAP7_75t_R _19800_ (.A1(_11571_),
    .A2(_11577_),
    .B(_11493_),
    .Y(_11580_));
 AO21x1_ASAP7_75t_SL _19801_ (.A1(_11451_),
    .A2(_11450_),
    .B(_11475_),
    .Y(_11581_));
 AND3x1_ASAP7_75t_R _19802_ (.A(_11572_),
    .B(_11470_),
    .C(_11581_),
    .Y(_11582_));
 NAND2x2_ASAP7_75t_SL _19803_ (.A(_11452_),
    .B(_11407_),
    .Y(_11583_));
 AO21x1_ASAP7_75t_SL _19804_ (.A1(_11407_),
    .A2(_11449_),
    .B(_11452_),
    .Y(_11584_));
 AOI21x1_ASAP7_75t_R _19805_ (.A1(_11583_),
    .A2(_11584_),
    .B(_11470_),
    .Y(_11585_));
 OAI21x1_ASAP7_75t_SL _19806_ (.A1(_11582_),
    .A2(_11585_),
    .B(_11489_),
    .Y(_11586_));
 NAND3x1_ASAP7_75t_SL _19807_ (.A(_11580_),
    .B(_11586_),
    .C(_11513_),
    .Y(_11587_));
 XNOR2x2_ASAP7_75t_R _19808_ (.A(_00589_),
    .B(_00621_),
    .Y(_11588_));
 INVx2_ASAP7_75t_R _19809_ (.A(_00686_),
    .Y(_11589_));
 XOR2x2_ASAP7_75t_SL _19810_ (.A(_11588_),
    .B(_11589_),
    .Y(_11590_));
 XNOR2x2_ASAP7_75t_SL _19811_ (.A(_00622_),
    .B(_00654_),
    .Y(_11591_));
 XOR2x2_ASAP7_75t_SL _19812_ (.A(_11590_),
    .B(_11591_),
    .Y(_11592_));
 NOR2x1_ASAP7_75t_SL _19813_ (.A(_00574_),
    .B(_00490_),
    .Y(_11593_));
 AO21x1_ASAP7_75t_SL _19814_ (.A1(_11592_),
    .A2(_00574_),
    .B(_11593_),
    .Y(_11594_));
 XOR2x2_ASAP7_75t_SL _19815_ (.A(_11594_),
    .B(_00894_),
    .Y(_11595_));
 INVx1_ASAP7_75t_SL _19816_ (.A(_11595_),
    .Y(_11596_));
 AOI21x1_ASAP7_75t_R _19817_ (.A1(_11567_),
    .A2(_11587_),
    .B(_11596_),
    .Y(_11597_));
 AO21x1_ASAP7_75t_SL _19819_ (.A1(_11537_),
    .A2(_11563_),
    .B(_11463_),
    .Y(_11599_));
 AND2x2_ASAP7_75t_SL _19820_ (.A(_01087_),
    .B(_01085_),
    .Y(_11600_));
 NOR2x1_ASAP7_75t_SL _19821_ (.A(_11600_),
    .B(_11452_),
    .Y(_11601_));
 AOI21x1_ASAP7_75t_SL _19822_ (.A1(_11449_),
    .A2(_11407_),
    .B(_11446_),
    .Y(_11602_));
 OAI21x1_ASAP7_75t_R _19823_ (.A1(_11601_),
    .A2(_11602_),
    .B(_11463_),
    .Y(_11603_));
 NAND2x1_ASAP7_75t_R _19824_ (.A(_11599_),
    .B(_11603_),
    .Y(_11604_));
 OR2x2_ASAP7_75t_R _19825_ (.A(_11463_),
    .B(_01097_),
    .Y(_11605_));
 AOI21x1_ASAP7_75t_SL _19826_ (.A1(_11439_),
    .A2(_11445_),
    .B(_01084_),
    .Y(_11606_));
 AOI21x1_ASAP7_75t_SL _19827_ (.A1(_11606_),
    .A2(_11463_),
    .B(_11493_),
    .Y(_11607_));
 AOI21x1_ASAP7_75t_R _19828_ (.A1(_11605_),
    .A2(_11607_),
    .B(_11513_),
    .Y(_11608_));
 OAI21x1_ASAP7_75t_R _19829_ (.A1(_11489_),
    .A2(_11604_),
    .B(_11608_),
    .Y(_11609_));
 AO21x1_ASAP7_75t_R _19831_ (.A1(_11445_),
    .A2(_11439_),
    .B(_01087_),
    .Y(_11611_));
 OAI21x1_ASAP7_75t_SL _19832_ (.A1(_11470_),
    .A2(_11611_),
    .B(_11493_),
    .Y(_11612_));
 INVx1_ASAP7_75t_SL _19833_ (.A(_11612_),
    .Y(_11613_));
 OAI21x1_ASAP7_75t_SL _19834_ (.A1(_11573_),
    .A2(_11576_),
    .B(_11613_),
    .Y(_11614_));
 NOR2x1_ASAP7_75t_SL _19836_ (.A(_01087_),
    .B(_11452_),
    .Y(_11616_));
 AOI21x1_ASAP7_75t_SL _19837_ (.A1(_11463_),
    .A2(_11616_),
    .B(_11493_),
    .Y(_11617_));
 NOR2x2_ASAP7_75t_SL _19838_ (.A(_11463_),
    .B(_11479_),
    .Y(_11618_));
 INVx1_ASAP7_75t_R _19839_ (.A(_01090_),
    .Y(_11619_));
 NAND3x1_ASAP7_75t_SL _19840_ (.A(_11445_),
    .B(_11619_),
    .C(_11439_),
    .Y(_11620_));
 NOR2x1_ASAP7_75t_L _19841_ (.A(_11470_),
    .B(_11620_),
    .Y(_11621_));
 NOR2x1p5_ASAP7_75t_SL _19842_ (.A(_11621_),
    .B(_11618_),
    .Y(_11622_));
 AOI21x1_ASAP7_75t_SL _19843_ (.A1(_11617_),
    .A2(_11622_),
    .B(_11512_),
    .Y(_11623_));
 AOI21x1_ASAP7_75t_SL _19844_ (.A1(_11623_),
    .A2(_11614_),
    .B(_11549_),
    .Y(_11624_));
 NAND2x1_ASAP7_75t_SL _19845_ (.A(_11624_),
    .B(_11609_),
    .Y(_11625_));
 INVx2_ASAP7_75t_SL _19846_ (.A(_11606_),
    .Y(_11626_));
 AOI21x1_ASAP7_75t_SL _19847_ (.A1(_11452_),
    .A2(_11407_),
    .B(_11470_),
    .Y(_11627_));
 NAND2x1p5_ASAP7_75t_SL _19848_ (.A(_11627_),
    .B(_11626_),
    .Y(_11628_));
 INVx1_ASAP7_75t_SL _19849_ (.A(_11562_),
    .Y(_11629_));
 OAI21x1_ASAP7_75t_R _19850_ (.A1(_11531_),
    .A2(_11629_),
    .B(_11470_),
    .Y(_11630_));
 AOI21x1_ASAP7_75t_SL _19852_ (.A1(_11628_),
    .A2(_11630_),
    .B(_11489_),
    .Y(_11632_));
 INVx1_ASAP7_75t_R _19853_ (.A(_11523_),
    .Y(_11633_));
 OAI21x1_ASAP7_75t_R _19854_ (.A1(_11633_),
    .A2(_11569_),
    .B(_11463_),
    .Y(_11634_));
 AOI21x1_ASAP7_75t_R _19855_ (.A1(_11498_),
    .A2(_11634_),
    .B(_11493_),
    .Y(_11635_));
 OAI21x1_ASAP7_75t_R _19856_ (.A1(_11632_),
    .A2(_11635_),
    .B(_11513_),
    .Y(_11636_));
 OA21x2_ASAP7_75t_R _19858_ (.A1(_11568_),
    .A2(_11470_),
    .B(_11493_),
    .Y(_11638_));
 NAND3x2_ASAP7_75t_SL _19859_ (.B(_11449_),
    .C(_11452_),
    .Y(_11639_),
    .A(_11407_));
 OA21x2_ASAP7_75t_SL _19860_ (.A1(_11452_),
    .A2(_11619_),
    .B(_11470_),
    .Y(_11640_));
 NAND2x1_ASAP7_75t_SL _19862_ (.A(_11639_),
    .B(_11640_),
    .Y(_11642_));
 NAND2x1_ASAP7_75t_L _19863_ (.A(_11638_),
    .B(_11642_),
    .Y(_11643_));
 AOI21x1_ASAP7_75t_SL _19864_ (.A1(_11470_),
    .A2(_11569_),
    .B(_11493_),
    .Y(_11644_));
 AOI21x1_ASAP7_75t_SL _19865_ (.A1(_11525_),
    .A2(_11446_),
    .B(_11470_),
    .Y(_11645_));
 NAND2x1_ASAP7_75t_R _19866_ (.A(_11645_),
    .B(_11639_),
    .Y(_11646_));
 AOI21x1_ASAP7_75t_R _19867_ (.A1(_11644_),
    .A2(_11646_),
    .B(_11513_),
    .Y(_11647_));
 XOR2x2_ASAP7_75t_SL _19868_ (.A(_11548_),
    .B(_08778_),
    .Y(_11648_));
 AOI21x1_ASAP7_75t_R _19870_ (.A1(_11643_),
    .A2(_11647_),
    .B(_11648_),
    .Y(_11650_));
 NAND2x1_ASAP7_75t_SL _19871_ (.A(_11636_),
    .B(_11650_),
    .Y(_11651_));
 AOI21x1_ASAP7_75t_SL _19872_ (.A1(_11651_),
    .A2(_11625_),
    .B(_11595_),
    .Y(_11652_));
 AOI21x1_ASAP7_75t_SL _19873_ (.A1(_11551_),
    .A2(_11597_),
    .B(_11652_),
    .Y(_00040_));
 AO21x1_ASAP7_75t_SL _19874_ (.A1(_11451_),
    .A2(_11450_),
    .B(_01087_),
    .Y(_11653_));
 OA21x2_ASAP7_75t_SL _19875_ (.A1(_11653_),
    .A2(_11470_),
    .B(_11493_),
    .Y(_11654_));
 OAI21x1_ASAP7_75t_SL _19876_ (.A1(_11479_),
    .A2(_11517_),
    .B(_11470_),
    .Y(_11655_));
 AOI21x1_ASAP7_75t_SL _19877_ (.A1(_11654_),
    .A2(_11655_),
    .B(_11648_),
    .Y(_11656_));
 AOI21x1_ASAP7_75t_SL _19878_ (.A1(_01088_),
    .A2(_11407_),
    .B(_11446_),
    .Y(_11657_));
 NAND2x1_ASAP7_75t_SL _19879_ (.A(_11463_),
    .B(_11657_),
    .Y(_11658_));
 AO21x1_ASAP7_75t_SL _19880_ (.A1(_11445_),
    .A2(_11439_),
    .B(_01092_),
    .Y(_11659_));
 NAND2x1_ASAP7_75t_SL _19882_ (.A(_11659_),
    .B(_11583_),
    .Y(_11661_));
 AOI21x1_ASAP7_75t_SL _19883_ (.A1(_11470_),
    .A2(_11661_),
    .B(_11493_),
    .Y(_11662_));
 NAND2x1_ASAP7_75t_SL _19884_ (.A(_11658_),
    .B(_11662_),
    .Y(_11663_));
 NAND2x1_ASAP7_75t_SL _19885_ (.A(_11656_),
    .B(_11663_),
    .Y(_11664_));
 NOR2x1p5_ASAP7_75t_SL _19887_ (.A(_11606_),
    .B(_11470_),
    .Y(_11666_));
 AOI21x1_ASAP7_75t_SL _19889_ (.A1(_11666_),
    .A2(_11467_),
    .B(_11489_),
    .Y(_11668_));
 AO21x1_ASAP7_75t_SL _19890_ (.A1(_11574_),
    .A2(_11467_),
    .B(_11463_),
    .Y(_11669_));
 AOI21x1_ASAP7_75t_SL _19892_ (.A1(_11668_),
    .A2(_11669_),
    .B(_11549_),
    .Y(_11671_));
 AND2x2_ASAP7_75t_SL _19893_ (.A(_11611_),
    .B(_11618_),
    .Y(_11672_));
 AND3x1_ASAP7_75t_SL _19894_ (.A(_11537_),
    .B(_11463_),
    .C(_11563_),
    .Y(_11673_));
 OAI21x1_ASAP7_75t_SL _19895_ (.A1(_11673_),
    .A2(_11672_),
    .B(_11489_),
    .Y(_11674_));
 NAND2x1_ASAP7_75t_SL _19896_ (.A(_11674_),
    .B(_11671_),
    .Y(_11675_));
 AOI21x1_ASAP7_75t_SL _19898_ (.A1(_11675_),
    .A2(_11664_),
    .B(_11512_),
    .Y(_11677_));
 INVx1_ASAP7_75t_SL _19899_ (.A(_11537_),
    .Y(_11678_));
 AO21x1_ASAP7_75t_SL _19900_ (.A1(_11452_),
    .A2(_01087_),
    .B(_11470_),
    .Y(_11679_));
 NOR2x1_ASAP7_75t_SL _19901_ (.A(_11678_),
    .B(_11679_),
    .Y(_11680_));
 AO21x1_ASAP7_75t_SL _19903_ (.A1(_11572_),
    .A2(_11618_),
    .B(_11493_),
    .Y(_11682_));
 NOR2x2_ASAP7_75t_SL _19904_ (.A(_11452_),
    .B(_11463_),
    .Y(_11683_));
 AOI21x1_ASAP7_75t_SL _19905_ (.A1(_11683_),
    .A2(_11499_),
    .B(_11489_),
    .Y(_11684_));
 NAND2x1_ASAP7_75t_SL _19906_ (.A(_11530_),
    .B(_11627_),
    .Y(_11685_));
 AOI21x1_ASAP7_75t_SL _19908_ (.A1(_11684_),
    .A2(_11685_),
    .B(_11648_),
    .Y(_11687_));
 OAI21x1_ASAP7_75t_SL _19909_ (.A1(_11680_),
    .A2(_11682_),
    .B(_11687_),
    .Y(_11688_));
 AOI21x1_ASAP7_75t_SL _19910_ (.A1(_11446_),
    .A2(_11407_),
    .B(_11463_),
    .Y(_11689_));
 NOR2x1_ASAP7_75t_SL _19911_ (.A(_11446_),
    .B(_11407_),
    .Y(_11690_));
 AOI211x1_ASAP7_75t_SL _19912_ (.A1(_11463_),
    .A2(_11616_),
    .B(_11689_),
    .C(_11690_),
    .Y(_11691_));
 NAND2x1_ASAP7_75t_SL _19913_ (.A(_11489_),
    .B(_11691_),
    .Y(_11692_));
 OAI21x1_ASAP7_75t_SL _19914_ (.A1(_11616_),
    .A2(_11602_),
    .B(_11463_),
    .Y(_11693_));
 AOI21x1_ASAP7_75t_SL _19915_ (.A1(_11581_),
    .A2(_11557_),
    .B(_11489_),
    .Y(_11694_));
 AOI21x1_ASAP7_75t_SL _19916_ (.A1(_11693_),
    .A2(_11694_),
    .B(_11549_),
    .Y(_11695_));
 NAND2x1_ASAP7_75t_SL _19917_ (.A(_11692_),
    .B(_11695_),
    .Y(_11696_));
 AOI21x1_ASAP7_75t_SL _19918_ (.A1(_11688_),
    .A2(_11696_),
    .B(_11513_),
    .Y(_11697_));
 OAI21x1_ASAP7_75t_SL _19919_ (.A1(_11697_),
    .A2(_11677_),
    .B(_11596_),
    .Y(_11698_));
 NOR2x1_ASAP7_75t_SL _19920_ (.A(_11501_),
    .B(_11576_),
    .Y(_11699_));
 OA21x2_ASAP7_75t_SL _19921_ (.A1(_11452_),
    .A2(_01083_),
    .B(_11463_),
    .Y(_11700_));
 AO21x1_ASAP7_75t_SL _19922_ (.A1(_11700_),
    .A2(_11467_),
    .B(_11648_),
    .Y(_11701_));
 INVx2_ASAP7_75t_SL _19923_ (.A(_11570_),
    .Y(_11702_));
 NAND2x1_ASAP7_75t_SL _19924_ (.A(_11497_),
    .B(_11702_),
    .Y(_11703_));
 AOI21x1_ASAP7_75t_SL _19925_ (.A1(_11552_),
    .A2(_11532_),
    .B(_11549_),
    .Y(_11704_));
 NAND2x1_ASAP7_75t_SL _19926_ (.A(_11703_),
    .B(_11704_),
    .Y(_11705_));
 OAI21x1_ASAP7_75t_SL _19927_ (.A1(_11699_),
    .A2(_11701_),
    .B(_11705_),
    .Y(_11706_));
 INVx1_ASAP7_75t_SL _19928_ (.A(_11645_),
    .Y(_11707_));
 NOR2x1_ASAP7_75t_SL _19929_ (.A(_11446_),
    .B(_11574_),
    .Y(_11708_));
 OAI21x1_ASAP7_75t_SL _19930_ (.A1(_11707_),
    .A2(_11708_),
    .B(_11493_),
    .Y(_11709_));
 AND3x1_ASAP7_75t_SL _19931_ (.A(_11648_),
    .B(_01099_),
    .C(_11470_),
    .Y(_11710_));
 OAI21x1_ASAP7_75t_SL _19932_ (.A1(_11709_),
    .A2(_11710_),
    .B(_11512_),
    .Y(_11711_));
 AOI21x1_ASAP7_75t_SL _19933_ (.A1(_11489_),
    .A2(_11706_),
    .B(_11711_),
    .Y(_11712_));
 AO21x1_ASAP7_75t_SL _19934_ (.A1(_11451_),
    .A2(_11450_),
    .B(_01092_),
    .Y(_11713_));
 AO21x1_ASAP7_75t_SL _19935_ (.A1(_11445_),
    .A2(_11439_),
    .B(_01085_),
    .Y(_11714_));
 AO21x1_ASAP7_75t_SL _19936_ (.A1(_11713_),
    .A2(_11714_),
    .B(_11470_),
    .Y(_11715_));
 NAND2x1_ASAP7_75t_SL _19937_ (.A(_11715_),
    .B(_11655_),
    .Y(_11716_));
 NOR2x1p5_ASAP7_75t_SL _19938_ (.A(_11489_),
    .B(_11618_),
    .Y(_11717_));
 OAI21x1_ASAP7_75t_SL _19939_ (.A1(_11678_),
    .A2(_11657_),
    .B(_11463_),
    .Y(_11718_));
 AOI21x1_ASAP7_75t_SL _19940_ (.A1(_11717_),
    .A2(_11718_),
    .B(_11549_),
    .Y(_11719_));
 OAI21x1_ASAP7_75t_SL _19941_ (.A1(_11493_),
    .A2(_11716_),
    .B(_11719_),
    .Y(_11720_));
 AO21x1_ASAP7_75t_SL _19942_ (.A1(_11626_),
    .A2(_11563_),
    .B(_11463_),
    .Y(_11721_));
 AO21x1_ASAP7_75t_SL _19943_ (.A1(_11537_),
    .A2(_11568_),
    .B(_11470_),
    .Y(_11722_));
 NAND2x1_ASAP7_75t_SL _19944_ (.A(_11721_),
    .B(_11722_),
    .Y(_11723_));
 AO21x1_ASAP7_75t_SL _19945_ (.A1(_11467_),
    .A2(_11523_),
    .B(_11470_),
    .Y(_11724_));
 AOI21x1_ASAP7_75t_SL _19947_ (.A1(_11497_),
    .A2(_11702_),
    .B(_11489_),
    .Y(_11726_));
 AOI21x1_ASAP7_75t_SL _19948_ (.A1(_11724_),
    .A2(_11726_),
    .B(_11648_),
    .Y(_11727_));
 OAI21x1_ASAP7_75t_SL _19949_ (.A1(_11493_),
    .A2(_11723_),
    .B(_11727_),
    .Y(_11728_));
 AOI21x1_ASAP7_75t_SL _19950_ (.A1(_11720_),
    .A2(_11728_),
    .B(_11512_),
    .Y(_11729_));
 OAI21x1_ASAP7_75t_SL _19951_ (.A1(_11712_),
    .A2(_11729_),
    .B(_11595_),
    .Y(_11730_));
 NAND2x1_ASAP7_75t_SL _19952_ (.A(_11698_),
    .B(_11730_),
    .Y(_00041_));
 NAND2x1_ASAP7_75t_R _19953_ (.A(_01099_),
    .B(_11463_),
    .Y(_11731_));
 AND2x2_ASAP7_75t_SL _19954_ (.A(_11583_),
    .B(_11470_),
    .Y(_11732_));
 AOI21x1_ASAP7_75t_SL _19955_ (.A1(_11530_),
    .A2(_11732_),
    .B(_11489_),
    .Y(_11733_));
 AOI21x1_ASAP7_75t_R _19957_ (.A1(_11731_),
    .A2(_11733_),
    .B(_11549_),
    .Y(_11735_));
 NAND2x1_ASAP7_75t_SL _19958_ (.A(_11523_),
    .B(_11627_),
    .Y(_11736_));
 NOR2x1_ASAP7_75t_SL _19959_ (.A(_11606_),
    .B(_11463_),
    .Y(_11737_));
 NAND2x1_ASAP7_75t_SL _19960_ (.A(_11737_),
    .B(_11526_),
    .Y(_11738_));
 AO21x1_ASAP7_75t_SL _19961_ (.A1(_11738_),
    .A2(_11736_),
    .B(_11493_),
    .Y(_11739_));
 AND2x2_ASAP7_75t_SL _19962_ (.A(_11735_),
    .B(_11739_),
    .Y(_11740_));
 NAND2x2_ASAP7_75t_SL _19963_ (.A(_11452_),
    .B(_01088_),
    .Y(_11741_));
 AO21x1_ASAP7_75t_SL _19964_ (.A1(_11552_),
    .A2(_11741_),
    .B(_11463_),
    .Y(_11742_));
 NAND3x1_ASAP7_75t_R _19965_ (.A(_11742_),
    .B(_11489_),
    .C(_11628_),
    .Y(_11743_));
 OA21x2_ASAP7_75t_R _19966_ (.A1(_01097_),
    .A2(_11470_),
    .B(_11493_),
    .Y(_11744_));
 NAND2x1_ASAP7_75t_R _19967_ (.A(_11639_),
    .B(_11557_),
    .Y(_11745_));
 AOI21x1_ASAP7_75t_R _19968_ (.A1(_11744_),
    .A2(_11745_),
    .B(_11648_),
    .Y(_11746_));
 AO21x1_ASAP7_75t_SL _19969_ (.A1(_11746_),
    .A2(_11743_),
    .B(_11512_),
    .Y(_11747_));
 NOR2x1_ASAP7_75t_SL _19970_ (.A(_11600_),
    .B(_11446_),
    .Y(_11748_));
 OA21x2_ASAP7_75t_R _19971_ (.A1(_11517_),
    .A2(_11748_),
    .B(_11470_),
    .Y(_11749_));
 OAI21x1_ASAP7_75t_R _19972_ (.A1(_11707_),
    .A2(_11708_),
    .B(_11489_),
    .Y(_11750_));
 INVx1_ASAP7_75t_SL _19973_ (.A(_01087_),
    .Y(_11751_));
 AO21x1_ASAP7_75t_R _19974_ (.A1(_11445_),
    .A2(_11439_),
    .B(_11751_),
    .Y(_11752_));
 NAND2x1p5_ASAP7_75t_SL _19975_ (.A(_11618_),
    .B(_11752_),
    .Y(_11753_));
 OA21x2_ASAP7_75t_R _19976_ (.A1(_11563_),
    .A2(_11470_),
    .B(_11493_),
    .Y(_11754_));
 AOI21x1_ASAP7_75t_SL _19977_ (.A1(_11754_),
    .A2(_11753_),
    .B(_11648_),
    .Y(_11755_));
 OAI21x1_ASAP7_75t_SL _19978_ (.A1(_11749_),
    .A2(_11750_),
    .B(_11755_),
    .Y(_11756_));
 OAI21x1_ASAP7_75t_SL _19979_ (.A1(_01082_),
    .A2(_11572_),
    .B(_11463_),
    .Y(_11757_));
 NAND2x1_ASAP7_75t_R _19980_ (.A(_01096_),
    .B(_11470_),
    .Y(_11758_));
 NAND3x1_ASAP7_75t_L _19981_ (.A(_11757_),
    .B(_11493_),
    .C(_11758_),
    .Y(_11759_));
 OA21x2_ASAP7_75t_R _19982_ (.A1(_01101_),
    .A2(_11470_),
    .B(_11489_),
    .Y(_11760_));
 NAND3x1_ASAP7_75t_SL _19983_ (.A(_11499_),
    .B(_11583_),
    .C(_11470_),
    .Y(_11761_));
 AOI21x1_ASAP7_75t_SL _19984_ (.A1(_11760_),
    .A2(_11761_),
    .B(_11549_),
    .Y(_11762_));
 AOI21x1_ASAP7_75t_R _19985_ (.A1(_11759_),
    .A2(_11762_),
    .B(_11513_),
    .Y(_11763_));
 AOI21x1_ASAP7_75t_SL _19986_ (.A1(_11763_),
    .A2(_11756_),
    .B(_11595_),
    .Y(_11764_));
 OAI21x1_ASAP7_75t_SL _19987_ (.A1(_11740_),
    .A2(_11747_),
    .B(_11764_),
    .Y(_11765_));
 NAND2x1p5_ASAP7_75t_SL _19988_ (.A(_11618_),
    .B(_11626_),
    .Y(_11766_));
 AOI21x1_ASAP7_75t_SL _19989_ (.A1(_01090_),
    .A2(_11446_),
    .B(_11470_),
    .Y(_11767_));
 NAND2x1_ASAP7_75t_SL _19990_ (.A(_11467_),
    .B(_11767_),
    .Y(_11768_));
 AOI21x1_ASAP7_75t_SL _19991_ (.A1(_11768_),
    .A2(_11766_),
    .B(_11489_),
    .Y(_11769_));
 NAND2x1_ASAP7_75t_SL _19992_ (.A(_11470_),
    .B(_11620_),
    .Y(_11770_));
 NOR2x1_ASAP7_75t_R _19993_ (.A(_11570_),
    .B(_11770_),
    .Y(_11771_));
 NAND2x1_ASAP7_75t_SL _19994_ (.A(_11463_),
    .B(_11659_),
    .Y(_11772_));
 OAI21x1_ASAP7_75t_R _19995_ (.A1(_11531_),
    .A2(_11772_),
    .B(_11489_),
    .Y(_11773_));
 NOR2x1_ASAP7_75t_R _19996_ (.A(_11771_),
    .B(_11773_),
    .Y(_11774_));
 OAI21x1_ASAP7_75t_SL _19997_ (.A1(_11774_),
    .A2(_11769_),
    .B(_11549_),
    .Y(_11775_));
 AO21x1_ASAP7_75t_R _19998_ (.A1(_11583_),
    .A2(_11611_),
    .B(_11463_),
    .Y(_11776_));
 NOR2x1_ASAP7_75t_R _19999_ (.A(_11621_),
    .B(_11612_),
    .Y(_11777_));
 NAND2x1_ASAP7_75t_R _20000_ (.A(_11776_),
    .B(_11777_),
    .Y(_11778_));
 AO21x1_ASAP7_75t_R _20001_ (.A1(_11741_),
    .A2(_11611_),
    .B(_11463_),
    .Y(_11779_));
 OAI21x1_ASAP7_75t_SL _20002_ (.A1(_11470_),
    .A2(_11659_),
    .B(_11489_),
    .Y(_11780_));
 NOR2x1_ASAP7_75t_R _20003_ (.A(_11621_),
    .B(_11780_),
    .Y(_11781_));
 AOI21x1_ASAP7_75t_R _20004_ (.A1(_11779_),
    .A2(_11781_),
    .B(_11549_),
    .Y(_11782_));
 NAND2x1_ASAP7_75t_R _20005_ (.A(_11778_),
    .B(_11782_),
    .Y(_11783_));
 AOI21x1_ASAP7_75t_SL _20006_ (.A1(_11783_),
    .A2(_11775_),
    .B(_11512_),
    .Y(_11784_));
 NAND2x1p5_ASAP7_75t_SL _20007_ (.A(_11463_),
    .B(_11519_),
    .Y(_11785_));
 NOR2x1_ASAP7_75t_R _20008_ (.A(_11570_),
    .B(_11785_),
    .Y(_11786_));
 AND3x1_ASAP7_75t_R _20009_ (.A(_11741_),
    .B(_11470_),
    .C(_11714_),
    .Y(_11787_));
 OAI21x1_ASAP7_75t_R _20010_ (.A1(_11786_),
    .A2(_11787_),
    .B(_11489_),
    .Y(_11788_));
 INVx1_ASAP7_75t_R _20011_ (.A(_11713_),
    .Y(_11789_));
 OAI21x1_ASAP7_75t_R _20012_ (.A1(_11789_),
    .A2(_11517_),
    .B(_11470_),
    .Y(_11790_));
 NAND3x1_ASAP7_75t_R _20013_ (.A(_11790_),
    .B(_11493_),
    .C(_11757_),
    .Y(_11791_));
 AOI21x1_ASAP7_75t_R _20014_ (.A1(_11788_),
    .A2(_11791_),
    .B(_11648_),
    .Y(_11792_));
 AO21x1_ASAP7_75t_R _20015_ (.A1(_11659_),
    .A2(_11653_),
    .B(_11470_),
    .Y(_11793_));
 AOI21x1_ASAP7_75t_R _20016_ (.A1(_11793_),
    .A2(_11761_),
    .B(_11493_),
    .Y(_11794_));
 AOI21x1_ASAP7_75t_R _20017_ (.A1(_11752_),
    .A2(_11639_),
    .B(_11463_),
    .Y(_11795_));
 INVx1_ASAP7_75t_SL _20018_ (.A(_11627_),
    .Y(_11796_));
 OAI21x1_ASAP7_75t_SL _20019_ (.A1(_11606_),
    .A2(_11796_),
    .B(_11493_),
    .Y(_11797_));
 OAI21x1_ASAP7_75t_SL _20020_ (.A1(_11795_),
    .A2(_11797_),
    .B(_11648_),
    .Y(_11798_));
 OAI21x1_ASAP7_75t_SL _20021_ (.A1(_11794_),
    .A2(_11798_),
    .B(_11512_),
    .Y(_11799_));
 NOR2x1_ASAP7_75t_SL _20022_ (.A(_11792_),
    .B(_11799_),
    .Y(_11800_));
 OAI21x1_ASAP7_75t_SL _20023_ (.A1(_11800_),
    .A2(_11784_),
    .B(_11595_),
    .Y(_11801_));
 NAND2x1_ASAP7_75t_SL _20024_ (.A(_11801_),
    .B(_11765_),
    .Y(_00042_));
 NAND2x1_ASAP7_75t_SL _20025_ (.A(_11600_),
    .B(_11452_),
    .Y(_11802_));
 NAND2x1_ASAP7_75t_SL _20026_ (.A(_11802_),
    .B(_11640_),
    .Y(_11803_));
 INVx1_ASAP7_75t_SL _20027_ (.A(_11803_),
    .Y(_11804_));
 NOR2x1_ASAP7_75t_SL _20028_ (.A(_11531_),
    .B(_11772_),
    .Y(_11805_));
 AOI21x1_ASAP7_75t_SL _20029_ (.A1(_11489_),
    .A2(_11805_),
    .B(_11549_),
    .Y(_11806_));
 OAI21x1_ASAP7_75t_SL _20030_ (.A1(_11709_),
    .A2(_11804_),
    .B(_11806_),
    .Y(_11807_));
 AOI21x1_ASAP7_75t_SL _20031_ (.A1(_11685_),
    .A2(_11599_),
    .B(_11489_),
    .Y(_11808_));
 AO21x1_ASAP7_75t_SL _20032_ (.A1(_11519_),
    .A2(_11659_),
    .B(_11470_),
    .Y(_11809_));
 AO21x1_ASAP7_75t_SL _20033_ (.A1(_11572_),
    .A2(_11620_),
    .B(_11463_),
    .Y(_11810_));
 AOI21x1_ASAP7_75t_SL _20034_ (.A1(_11809_),
    .A2(_11810_),
    .B(_11493_),
    .Y(_11811_));
 OAI21x1_ASAP7_75t_SL _20035_ (.A1(_11808_),
    .A2(_11811_),
    .B(_11549_),
    .Y(_11812_));
 AOI21x1_ASAP7_75t_SL _20036_ (.A1(_11807_),
    .A2(_11812_),
    .B(_11512_),
    .Y(_11813_));
 NAND2x1_ASAP7_75t_SL _20037_ (.A(_01084_),
    .B(_11683_),
    .Y(_11814_));
 NAND2x1_ASAP7_75t_SL _20038_ (.A(_11583_),
    .B(_11645_),
    .Y(_11815_));
 AOI21x1_ASAP7_75t_SL _20039_ (.A1(_11814_),
    .A2(_11815_),
    .B(_11549_),
    .Y(_11816_));
 AND2x4_ASAP7_75t_SL _20040_ (.A(_11479_),
    .B(_11463_),
    .Y(_11817_));
 INVx3_ASAP7_75t_SL _20041_ (.A(_11817_),
    .Y(_11818_));
 OAI21x1_ASAP7_75t_SL _20042_ (.A1(_11648_),
    .A2(_11818_),
    .B(_11644_),
    .Y(_11819_));
 OAI21x1_ASAP7_75t_SL _20043_ (.A1(_11819_),
    .A2(_11816_),
    .B(_11512_),
    .Y(_11820_));
 AO21x1_ASAP7_75t_SL _20044_ (.A1(_11537_),
    .A2(_11519_),
    .B(_11470_),
    .Y(_11821_));
 INVx1_ASAP7_75t_SL _20045_ (.A(_11748_),
    .Y(_11822_));
 AO21x1_ASAP7_75t_SL _20046_ (.A1(_11822_),
    .A2(_11659_),
    .B(_11463_),
    .Y(_11823_));
 AOI21x1_ASAP7_75t_SL _20047_ (.A1(_11821_),
    .A2(_11823_),
    .B(_11549_),
    .Y(_11824_));
 INVx1_ASAP7_75t_SL _20048_ (.A(_11620_),
    .Y(_11825_));
 AOI22x1_ASAP7_75t_SL _20049_ (.A1(_11470_),
    .A2(_11825_),
    .B1(_11767_),
    .B2(_11467_),
    .Y(_11826_));
 OAI21x1_ASAP7_75t_SL _20050_ (.A1(_11648_),
    .A2(_11826_),
    .B(_11493_),
    .Y(_11827_));
 NOR2x1_ASAP7_75t_SL _20051_ (.A(_11824_),
    .B(_11827_),
    .Y(_11828_));
 OAI21x1_ASAP7_75t_SL _20052_ (.A1(_11828_),
    .A2(_11820_),
    .B(_11595_),
    .Y(_11829_));
 NOR2x1_ASAP7_75t_SL _20053_ (.A(_11813_),
    .B(_11829_),
    .Y(_11830_));
 AOI21x1_ASAP7_75t_SL _20054_ (.A1(_11702_),
    .A2(_11618_),
    .B(_11489_),
    .Y(_11831_));
 NAND2x1_ASAP7_75t_SL _20055_ (.A(_11499_),
    .B(_11532_),
    .Y(_11832_));
 NAND2x1_ASAP7_75t_SL _20056_ (.A(_11832_),
    .B(_11831_),
    .Y(_11833_));
 AO21x1_ASAP7_75t_SL _20057_ (.A1(_11552_),
    .A2(_11741_),
    .B(_11470_),
    .Y(_11834_));
 AOI21x1_ASAP7_75t_SL _20058_ (.A1(_11558_),
    .A2(_11834_),
    .B(_11549_),
    .Y(_11835_));
 AOI21x1_ASAP7_75t_SL _20059_ (.A1(_11833_),
    .A2(_11835_),
    .B(_11513_),
    .Y(_11836_));
 AND2x2_ASAP7_75t_SL _20060_ (.A(_11537_),
    .B(_11526_),
    .Y(_11837_));
 AOI22x1_ASAP7_75t_SL _20061_ (.A1(_11563_),
    .A2(_11557_),
    .B1(_11837_),
    .B2(_11463_),
    .Y(_11838_));
 AO21x1_ASAP7_75t_SL _20062_ (.A1(_11713_),
    .A2(_11611_),
    .B(_11463_),
    .Y(_11839_));
 AOI21x1_ASAP7_75t_SL _20063_ (.A1(_11702_),
    .A2(_11553_),
    .B(_11489_),
    .Y(_11840_));
 AOI21x1_ASAP7_75t_SL _20064_ (.A1(_11839_),
    .A2(_11840_),
    .B(_11648_),
    .Y(_11841_));
 OAI21x1_ASAP7_75t_SL _20065_ (.A1(_11493_),
    .A2(_11838_),
    .B(_11841_),
    .Y(_11842_));
 NAND2x1_ASAP7_75t_SL _20066_ (.A(_11836_),
    .B(_11842_),
    .Y(_11843_));
 NAND2x1_ASAP7_75t_SL _20067_ (.A(_11452_),
    .B(_11470_),
    .Y(_11844_));
 AOI21x1_ASAP7_75t_SL _20068_ (.A1(_11741_),
    .A2(_11499_),
    .B(_11489_),
    .Y(_11845_));
 AOI21x1_ASAP7_75t_SL _20069_ (.A1(_11844_),
    .A2(_11845_),
    .B(_11549_),
    .Y(_11846_));
 AO21x1_ASAP7_75t_SL _20070_ (.A1(_01090_),
    .A2(_11446_),
    .B(_11785_),
    .Y(_11847_));
 NAND2x1_ASAP7_75t_SL _20071_ (.A(_11662_),
    .B(_11847_),
    .Y(_11848_));
 AOI21x1_ASAP7_75t_SL _20072_ (.A1(_11846_),
    .A2(_11848_),
    .B(_11512_),
    .Y(_11849_));
 INVx4_ASAP7_75t_SL _20073_ (.A(_11479_),
    .Y(_11850_));
 AND3x1_ASAP7_75t_SL _20074_ (.A(_11562_),
    .B(_11463_),
    .C(_11850_),
    .Y(_11851_));
 NOR2x1_ASAP7_75t_SL _20075_ (.A(_11539_),
    .B(_11851_),
    .Y(_11852_));
 NOR2x1_ASAP7_75t_SL _20076_ (.A(_11463_),
    .B(_11570_),
    .Y(_11853_));
 INVx2_ASAP7_75t_SL _20077_ (.A(_11666_),
    .Y(_11854_));
 OAI21x1_ASAP7_75t_SL _20078_ (.A1(_11854_),
    .A2(_11657_),
    .B(_11493_),
    .Y(_11855_));
 AOI21x1_ASAP7_75t_SL _20079_ (.A1(_11853_),
    .A2(_11837_),
    .B(_11855_),
    .Y(_11856_));
 OAI21x1_ASAP7_75t_SL _20080_ (.A1(_11856_),
    .A2(_11852_),
    .B(_11549_),
    .Y(_11857_));
 NAND2x1_ASAP7_75t_SL _20081_ (.A(_11857_),
    .B(_11849_),
    .Y(_11858_));
 AOI21x1_ASAP7_75t_SL _20082_ (.A1(_11843_),
    .A2(_11858_),
    .B(_11595_),
    .Y(_11859_));
 NOR2x1_ASAP7_75t_SL _20083_ (.A(_11830_),
    .B(_11859_),
    .Y(_00043_));
 NOR2x1_ASAP7_75t_SL _20084_ (.A(_11463_),
    .B(_11538_),
    .Y(_11860_));
 NOR2x1_ASAP7_75t_R _20085_ (.A(_11489_),
    .B(_11860_),
    .Y(_11861_));
 AND2x2_ASAP7_75t_SL _20086_ (.A(_11861_),
    .B(_11634_),
    .Y(_11862_));
 INVx2_ASAP7_75t_SL _20087_ (.A(_11690_),
    .Y(_11863_));
 AO21x1_ASAP7_75t_SL _20088_ (.A1(_11863_),
    .A2(_11574_),
    .B(_11470_),
    .Y(_11864_));
 AOI21x1_ASAP7_75t_R _20089_ (.A1(_11741_),
    .A2(_11640_),
    .B(_11493_),
    .Y(_11865_));
 AO21x1_ASAP7_75t_R _20090_ (.A1(_11864_),
    .A2(_11865_),
    .B(_11549_),
    .Y(_11866_));
 AO21x1_ASAP7_75t_R _20091_ (.A1(_01091_),
    .A2(_11463_),
    .B(_11489_),
    .Y(_11867_));
 OA21x2_ASAP7_75t_SL _20092_ (.A1(_11737_),
    .A2(_11867_),
    .B(_11549_),
    .Y(_11868_));
 NAND2x1_ASAP7_75t_R _20093_ (.A(_11463_),
    .B(_11602_),
    .Y(_11869_));
 AOI21x1_ASAP7_75t_SL _20094_ (.A1(_11863_),
    .A2(_11640_),
    .B(_11493_),
    .Y(_11870_));
 NAND2x1_ASAP7_75t_SL _20095_ (.A(_11869_),
    .B(_11870_),
    .Y(_11871_));
 AOI21x1_ASAP7_75t_SL _20096_ (.A1(_11871_),
    .A2(_11868_),
    .B(_11513_),
    .Y(_11872_));
 OAI21x1_ASAP7_75t_SL _20097_ (.A1(_11862_),
    .A2(_11866_),
    .B(_11872_),
    .Y(_11873_));
 NOR2x1_ASAP7_75t_R _20098_ (.A(_11489_),
    .B(_11683_),
    .Y(_11874_));
 AO21x1_ASAP7_75t_R _20099_ (.A1(_11467_),
    .A2(_11659_),
    .B(_11470_),
    .Y(_11875_));
 AOI21x1_ASAP7_75t_R _20100_ (.A1(_11874_),
    .A2(_11875_),
    .B(_11549_),
    .Y(_11876_));
 INVx2_ASAP7_75t_SL _20101_ (.A(_11563_),
    .Y(_11877_));
 AOI21x1_ASAP7_75t_R _20102_ (.A1(_11463_),
    .A2(_11877_),
    .B(_11493_),
    .Y(_11878_));
 NAND2x1_ASAP7_75t_R _20103_ (.A(_11463_),
    .B(_11570_),
    .Y(_11879_));
 NAND3x1_ASAP7_75t_L _20104_ (.A(_11878_),
    .B(_11703_),
    .C(_11879_),
    .Y(_11880_));
 AOI21x1_ASAP7_75t_R _20105_ (.A1(_11876_),
    .A2(_11880_),
    .B(_11512_),
    .Y(_11881_));
 OA21x2_ASAP7_75t_SL _20106_ (.A1(_11574_),
    .A2(_11452_),
    .B(_11470_),
    .Y(_11882_));
 AO21x1_ASAP7_75t_R _20107_ (.A1(_11446_),
    .A2(_01085_),
    .B(_11470_),
    .Y(_11883_));
 NAND2x1_ASAP7_75t_R _20108_ (.A(_11489_),
    .B(_11883_),
    .Y(_11884_));
 OA21x2_ASAP7_75t_SL _20109_ (.A1(_11882_),
    .A2(_11884_),
    .B(_11549_),
    .Y(_11885_));
 OA21x2_ASAP7_75t_SL _20110_ (.A1(_11606_),
    .A2(_11679_),
    .B(_11493_),
    .Y(_11886_));
 OAI21x1_ASAP7_75t_SL _20111_ (.A1(_11573_),
    .A2(_11576_),
    .B(_11886_),
    .Y(_11887_));
 NAND2x1_ASAP7_75t_SL _20112_ (.A(_11887_),
    .B(_11885_),
    .Y(_11888_));
 AOI21x1_ASAP7_75t_SL _20113_ (.A1(_11881_),
    .A2(_11888_),
    .B(_11596_),
    .Y(_11889_));
 NAND2x1_ASAP7_75t_SL _20114_ (.A(_11889_),
    .B(_11873_),
    .Y(_11890_));
 NAND2x1_ASAP7_75t_R _20115_ (.A(_11523_),
    .B(_11732_),
    .Y(_11891_));
 AOI21x1_ASAP7_75t_R _20116_ (.A1(_11864_),
    .A2(_11891_),
    .B(_11493_),
    .Y(_11892_));
 NAND2x1_ASAP7_75t_R _20117_ (.A(_11552_),
    .B(_11532_),
    .Y(_11893_));
 AO21x1_ASAP7_75t_R _20118_ (.A1(_11733_),
    .A2(_11893_),
    .B(_11549_),
    .Y(_11894_));
 OAI21x1_ASAP7_75t_SL _20119_ (.A1(_11689_),
    .A2(_11700_),
    .B(_11467_),
    .Y(_11895_));
 OAI21x1_ASAP7_75t_SL _20120_ (.A1(_11569_),
    .A2(_11640_),
    .B(_11489_),
    .Y(_11896_));
 OAI21x1_ASAP7_75t_R _20121_ (.A1(_11489_),
    .A2(_11895_),
    .B(_11896_),
    .Y(_11897_));
 AOI21x1_ASAP7_75t_R _20122_ (.A1(_11549_),
    .A2(_11897_),
    .B(_11512_),
    .Y(_11898_));
 OAI21x1_ASAP7_75t_R _20123_ (.A1(_11892_),
    .A2(_11894_),
    .B(_11898_),
    .Y(_11899_));
 NAND2x1_ASAP7_75t_SL _20124_ (.A(_11606_),
    .B(_11470_),
    .Y(_11900_));
 AND2x2_ASAP7_75t_SL _20125_ (.A(_11900_),
    .B(_11620_),
    .Y(_11901_));
 AOI21x1_ASAP7_75t_SL _20126_ (.A1(_11617_),
    .A2(_11901_),
    .B(_11648_),
    .Y(_11902_));
 AO21x1_ASAP7_75t_R _20127_ (.A1(_11445_),
    .A2(_11439_),
    .B(_11478_),
    .Y(_11903_));
 AND2x2_ASAP7_75t_R _20128_ (.A(_11581_),
    .B(_11463_),
    .Y(_11904_));
 AOI21x1_ASAP7_75t_R _20129_ (.A1(_11903_),
    .A2(_11904_),
    .B(_11489_),
    .Y(_11905_));
 NAND2x1_ASAP7_75t_SL _20130_ (.A(_11642_),
    .B(_11905_),
    .Y(_11906_));
 AOI21x1_ASAP7_75t_SL _20131_ (.A1(_11906_),
    .A2(_11902_),
    .B(_11513_),
    .Y(_11907_));
 INVx1_ASAP7_75t_R _20132_ (.A(_11639_),
    .Y(_11908_));
 AO21x1_ASAP7_75t_R _20133_ (.A1(_01082_),
    .A2(_11446_),
    .B(_11463_),
    .Y(_11909_));
 NOR2x1_ASAP7_75t_R _20134_ (.A(_11908_),
    .B(_11909_),
    .Y(_11910_));
 NAND2x1_ASAP7_75t_R _20135_ (.A(_11489_),
    .B(_11793_),
    .Y(_11911_));
 NAND2x1_ASAP7_75t_SL _20136_ (.A(_11563_),
    .B(_11552_),
    .Y(_11912_));
 AOI21x1_ASAP7_75t_R _20137_ (.A1(_11470_),
    .A2(_11912_),
    .B(_11489_),
    .Y(_11913_));
 AOI21x1_ASAP7_75t_SL _20138_ (.A1(_11693_),
    .A2(_11913_),
    .B(_11549_),
    .Y(_11914_));
 OAI21x1_ASAP7_75t_R _20139_ (.A1(_11910_),
    .A2(_11911_),
    .B(_11914_),
    .Y(_11915_));
 AOI21x1_ASAP7_75t_SL _20140_ (.A1(_11915_),
    .A2(_11907_),
    .B(_11595_),
    .Y(_11916_));
 NAND2x1_ASAP7_75t_SL _20141_ (.A(_11899_),
    .B(_11916_),
    .Y(_11917_));
 NAND2x1_ASAP7_75t_SL _20142_ (.A(_11890_),
    .B(_11917_),
    .Y(_00044_));
 NAND2x1_ASAP7_75t_SL _20143_ (.A(_01087_),
    .B(_11568_),
    .Y(_11918_));
 AOI22x1_ASAP7_75t_SL _20144_ (.A1(_11918_),
    .A2(_11470_),
    .B1(_11639_),
    .B2(_11767_),
    .Y(_11919_));
 NAND2x1_ASAP7_75t_SL _20145_ (.A(_11489_),
    .B(_11919_),
    .Y(_11920_));
 NAND2x1_ASAP7_75t_SL _20146_ (.A(_11476_),
    .B(_11497_),
    .Y(_11921_));
 OAI21x1_ASAP7_75t_SL _20147_ (.A1(_11407_),
    .A2(_11452_),
    .B(_11568_),
    .Y(_11922_));
 AOI21x1_ASAP7_75t_SL _20148_ (.A1(_11463_),
    .A2(_11922_),
    .B(_11489_),
    .Y(_11923_));
 AOI21x1_ASAP7_75t_SL _20149_ (.A1(_11921_),
    .A2(_11923_),
    .B(_11512_),
    .Y(_11924_));
 AOI21x1_ASAP7_75t_SL _20150_ (.A1(_11920_),
    .A2(_11924_),
    .B(_11648_),
    .Y(_11925_));
 NOR2x1_ASAP7_75t_SL _20151_ (.A(_11629_),
    .B(_11657_),
    .Y(_11926_));
 INVx1_ASAP7_75t_SL _20152_ (.A(_11574_),
    .Y(_11927_));
 OAI21x1_ASAP7_75t_SL _20153_ (.A1(_11466_),
    .A2(_11927_),
    .B(_11489_),
    .Y(_11928_));
 AOI21x1_ASAP7_75t_SL _20154_ (.A1(_11470_),
    .A2(_11926_),
    .B(_11928_),
    .Y(_11929_));
 OA21x2_ASAP7_75t_SL _20155_ (.A1(_11407_),
    .A2(_11463_),
    .B(_11493_),
    .Y(_11930_));
 AND2x2_ASAP7_75t_SL _20156_ (.A(_11864_),
    .B(_11930_),
    .Y(_11931_));
 OAI21x1_ASAP7_75t_SL _20157_ (.A1(_11929_),
    .A2(_11931_),
    .B(_11512_),
    .Y(_11932_));
 AND2x2_ASAP7_75t_SL _20158_ (.A(_11925_),
    .B(_11932_),
    .Y(_11933_));
 AOI21x1_ASAP7_75t_SL _20159_ (.A1(_11683_),
    .A2(_11499_),
    .B(_11493_),
    .Y(_11934_));
 AOI21x1_ASAP7_75t_SL _20160_ (.A1(_11679_),
    .A2(_11934_),
    .B(_11512_),
    .Y(_11935_));
 AOI21x1_ASAP7_75t_SL _20161_ (.A1(_11449_),
    .A2(_11683_),
    .B(_11489_),
    .Y(_11936_));
 INVx1_ASAP7_75t_SL _20162_ (.A(_11936_),
    .Y(_11937_));
 AO21x1_ASAP7_75t_SL _20163_ (.A1(_11818_),
    .A2(_11770_),
    .B(_11937_),
    .Y(_11938_));
 AOI21x1_ASAP7_75t_SL _20164_ (.A1(_11935_),
    .A2(_11938_),
    .B(_11549_),
    .Y(_11939_));
 NOR2x1_ASAP7_75t_SL _20165_ (.A(_01085_),
    .B(_11452_),
    .Y(_11940_));
 OAI21x1_ASAP7_75t_SL _20166_ (.A1(_11940_),
    .A2(_11690_),
    .B(_11463_),
    .Y(_11941_));
 AOI21x1_ASAP7_75t_SL _20167_ (.A1(_11900_),
    .A2(_11941_),
    .B(_11493_),
    .Y(_11942_));
 NAND2x1_ASAP7_75t_SL _20168_ (.A(_11523_),
    .B(_11618_),
    .Y(_11943_));
 AND3x1_ASAP7_75t_SL _20169_ (.A(_11943_),
    .B(_11493_),
    .C(_11772_),
    .Y(_11944_));
 OAI21x1_ASAP7_75t_SL _20170_ (.A1(_11942_),
    .A2(_11944_),
    .B(_11512_),
    .Y(_11945_));
 AO21x1_ASAP7_75t_SL _20171_ (.A1(_11945_),
    .A2(_11939_),
    .B(_11595_),
    .Y(_11946_));
 OAI21x1_ASAP7_75t_SL _20172_ (.A1(_11452_),
    .A2(_11499_),
    .B(_11618_),
    .Y(_11947_));
 NAND2x1_ASAP7_75t_SL _20173_ (.A(_11767_),
    .B(_11863_),
    .Y(_11948_));
 AND3x1_ASAP7_75t_SL _20174_ (.A(_11947_),
    .B(_11489_),
    .C(_11948_),
    .Y(_11949_));
 OA21x2_ASAP7_75t_SL _20175_ (.A1(_11449_),
    .A2(_11463_),
    .B(_11493_),
    .Y(_11950_));
 AO21x1_ASAP7_75t_SL _20176_ (.A1(_11533_),
    .A2(_11950_),
    .B(_11648_),
    .Y(_11951_));
 OAI21x1_ASAP7_75t_SL _20177_ (.A1(_11949_),
    .A2(_11951_),
    .B(_11513_),
    .Y(_11952_));
 NOR2x1_ASAP7_75t_SL _20178_ (.A(_11470_),
    .B(_11741_),
    .Y(_11953_));
 OA21x2_ASAP7_75t_SL _20179_ (.A1(_11562_),
    .A2(_11463_),
    .B(_11489_),
    .Y(_11954_));
 NOR2x1_ASAP7_75t_R _20180_ (.A(_01088_),
    .B(_11470_),
    .Y(_11955_));
 OAI21x1_ASAP7_75t_SL _20181_ (.A1(_11955_),
    .A2(_11627_),
    .B(_11476_),
    .Y(_11956_));
 AOI21x1_ASAP7_75t_SL _20182_ (.A1(_11954_),
    .A2(_11956_),
    .B(_11549_),
    .Y(_11957_));
 OA21x2_ASAP7_75t_SL _20183_ (.A1(_11614_),
    .A2(_11953_),
    .B(_11957_),
    .Y(_11958_));
 AOI21x1_ASAP7_75t_SL _20184_ (.A1(_11477_),
    .A2(_11617_),
    .B(_11648_),
    .Y(_11959_));
 AOI21x1_ASAP7_75t_SL _20185_ (.A1(_11470_),
    .A2(_11802_),
    .B(_11489_),
    .Y(_11960_));
 OAI21x1_ASAP7_75t_SL _20186_ (.A1(_11708_),
    .A2(_11757_),
    .B(_11960_),
    .Y(_11961_));
 AOI21x1_ASAP7_75t_SL _20187_ (.A1(_11959_),
    .A2(_11961_),
    .B(_11513_),
    .Y(_11962_));
 OA21x2_ASAP7_75t_SL _20188_ (.A1(_01089_),
    .A2(_11452_),
    .B(_11618_),
    .Y(_11963_));
 AO21x1_ASAP7_75t_SL _20189_ (.A1(_11463_),
    .A2(_11479_),
    .B(_11780_),
    .Y(_11964_));
 OA21x2_ASAP7_75t_SL _20190_ (.A1(_11525_),
    .A2(_11463_),
    .B(_11493_),
    .Y(_11965_));
 NOR2x1_ASAP7_75t_SL _20191_ (.A(_11955_),
    .B(_11627_),
    .Y(_11966_));
 AOI21x1_ASAP7_75t_SL _20192_ (.A1(_11965_),
    .A2(_11966_),
    .B(_11549_),
    .Y(_11967_));
 OAI21x1_ASAP7_75t_SL _20193_ (.A1(_11963_),
    .A2(_11964_),
    .B(_11967_),
    .Y(_11968_));
 AOI21x1_ASAP7_75t_SL _20194_ (.A1(_11962_),
    .A2(_11968_),
    .B(_11596_),
    .Y(_11969_));
 OAI21x1_ASAP7_75t_SL _20195_ (.A1(_11952_),
    .A2(_11958_),
    .B(_11969_),
    .Y(_11970_));
 OAI21x1_ASAP7_75t_SL _20196_ (.A1(_11933_),
    .A2(_11946_),
    .B(_11970_),
    .Y(_00045_));
 AO21x1_ASAP7_75t_SL _20197_ (.A1(_11463_),
    .A2(_11479_),
    .B(_11493_),
    .Y(_11971_));
 AO21x1_ASAP7_75t_SL _20198_ (.A1(_11757_),
    .A2(_11758_),
    .B(_11971_),
    .Y(_11972_));
 OA21x2_ASAP7_75t_R _20199_ (.A1(_11940_),
    .A2(_11479_),
    .B(_11463_),
    .Y(_11973_));
 AOI21x1_ASAP7_75t_R _20200_ (.A1(_11583_),
    .A2(_11584_),
    .B(_11463_),
    .Y(_11974_));
 OAI21x1_ASAP7_75t_R _20201_ (.A1(_11973_),
    .A2(_11974_),
    .B(_11493_),
    .Y(_11975_));
 AOI21x1_ASAP7_75t_SL _20202_ (.A1(_11975_),
    .A2(_11972_),
    .B(_11648_),
    .Y(_11976_));
 OA21x2_ASAP7_75t_R _20203_ (.A1(_11562_),
    .A2(_11470_),
    .B(_11489_),
    .Y(_11977_));
 NAND2x1_ASAP7_75t_R _20204_ (.A(_11499_),
    .B(_11689_),
    .Y(_11978_));
 AO21x1_ASAP7_75t_R _20205_ (.A1(_11977_),
    .A2(_11978_),
    .B(_11549_),
    .Y(_11979_));
 AOI211x1_ASAP7_75t_R _20206_ (.A1(_11666_),
    .A2(_11802_),
    .B(_11860_),
    .C(_11937_),
    .Y(_11980_));
 OAI21x1_ASAP7_75t_R _20207_ (.A1(_11979_),
    .A2(_11980_),
    .B(_11512_),
    .Y(_11981_));
 NOR2x1_ASAP7_75t_SL _20208_ (.A(_11981_),
    .B(_11976_),
    .Y(_11982_));
 AND2x2_ASAP7_75t_SL _20209_ (.A(_11767_),
    .B(_11581_),
    .Y(_11983_));
 OA21x2_ASAP7_75t_R _20210_ (.A1(_11517_),
    .A2(_11569_),
    .B(_11470_),
    .Y(_11984_));
 OAI21x1_ASAP7_75t_R _20211_ (.A1(_11983_),
    .A2(_11984_),
    .B(_11493_),
    .Y(_11985_));
 OR3x1_ASAP7_75t_SL _20212_ (.A(_11825_),
    .B(_11463_),
    .C(_11601_),
    .Y(_11986_));
 OA21x2_ASAP7_75t_R _20213_ (.A1(_11470_),
    .A2(_11741_),
    .B(_11607_),
    .Y(_11987_));
 AOI21x1_ASAP7_75t_R _20214_ (.A1(_11986_),
    .A2(_11987_),
    .B(_11549_),
    .Y(_11988_));
 AO21x1_ASAP7_75t_SL _20215_ (.A1(_11714_),
    .A2(_11620_),
    .B(_11463_),
    .Y(_11989_));
 NAND2x1_ASAP7_75t_R _20216_ (.A(_11878_),
    .B(_11989_),
    .Y(_11990_));
 INVx1_ASAP7_75t_R _20217_ (.A(_11499_),
    .Y(_11991_));
 AND2x2_ASAP7_75t_R _20218_ (.A(_01100_),
    .B(_01094_),
    .Y(_11992_));
 OA21x2_ASAP7_75t_R _20219_ (.A1(_11470_),
    .A2(_11992_),
    .B(_11493_),
    .Y(_11993_));
 OAI21x1_ASAP7_75t_R _20220_ (.A1(_11991_),
    .A2(_11909_),
    .B(_11993_),
    .Y(_11994_));
 AOI21x1_ASAP7_75t_R _20221_ (.A1(_11990_),
    .A2(_11994_),
    .B(_11648_),
    .Y(_11995_));
 AOI21x1_ASAP7_75t_R _20222_ (.A1(_11985_),
    .A2(_11988_),
    .B(_11995_),
    .Y(_11996_));
 OAI21x1_ASAP7_75t_SL _20223_ (.A1(_11512_),
    .A2(_11996_),
    .B(_11596_),
    .Y(_11997_));
 AOI21x1_ASAP7_75t_R _20224_ (.A1(_01095_),
    .A2(_11470_),
    .B(_11489_),
    .Y(_11998_));
 AOI21x1_ASAP7_75t_R _20225_ (.A1(_11998_),
    .A2(_11948_),
    .B(_11648_),
    .Y(_11999_));
 AO21x1_ASAP7_75t_SL _20226_ (.A1(_11850_),
    .A2(_11659_),
    .B(_11463_),
    .Y(_12000_));
 OA21x2_ASAP7_75t_R _20227_ (.A1(_11537_),
    .A2(_11470_),
    .B(_11489_),
    .Y(_12001_));
 NAND2x1_ASAP7_75t_SL _20228_ (.A(_12001_),
    .B(_12000_),
    .Y(_12002_));
 AOI21x1_ASAP7_75t_SL _20229_ (.A1(_11999_),
    .A2(_12002_),
    .B(_11513_),
    .Y(_12003_));
 NAND2x1_ASAP7_75t_R _20230_ (.A(_11493_),
    .B(_11795_),
    .Y(_12004_));
 AOI21x1_ASAP7_75t_R _20231_ (.A1(_11707_),
    .A2(_11870_),
    .B(_11549_),
    .Y(_12005_));
 NAND2x1_ASAP7_75t_SL _20232_ (.A(_12004_),
    .B(_12005_),
    .Y(_12006_));
 AOI21x1_ASAP7_75t_SL _20233_ (.A1(_12006_),
    .A2(_12003_),
    .B(_11596_),
    .Y(_12007_));
 AO21x1_ASAP7_75t_R _20234_ (.A1(_11845_),
    .A2(_11465_),
    .B(_11648_),
    .Y(_12008_));
 AO21x1_ASAP7_75t_R _20235_ (.A1(_11470_),
    .A2(_11530_),
    .B(_11904_),
    .Y(_12009_));
 AOI21x1_ASAP7_75t_R _20236_ (.A1(_11537_),
    .A2(_12009_),
    .B(_11493_),
    .Y(_12010_));
 NAND2x1_ASAP7_75t_R _20237_ (.A(_11770_),
    .B(_11785_),
    .Y(_12011_));
 AOI21x1_ASAP7_75t_R _20238_ (.A1(_11936_),
    .A2(_12011_),
    .B(_11549_),
    .Y(_12012_));
 NOR2x1_ASAP7_75t_R _20239_ (.A(_11493_),
    .B(_11689_),
    .Y(_12013_));
 NAND2x1_ASAP7_75t_SL _20240_ (.A(_12013_),
    .B(_11469_),
    .Y(_12014_));
 AOI21x1_ASAP7_75t_R _20241_ (.A1(_12012_),
    .A2(_12014_),
    .B(_11512_),
    .Y(_12015_));
 OAI21x1_ASAP7_75t_R _20242_ (.A1(_12008_),
    .A2(_12010_),
    .B(_12015_),
    .Y(_12016_));
 NAND2x1_ASAP7_75t_SL _20243_ (.A(_12016_),
    .B(_12007_),
    .Y(_12017_));
 OAI21x1_ASAP7_75t_SL _20244_ (.A1(_11997_),
    .A2(_11982_),
    .B(_12017_),
    .Y(_00046_));
 OAI21x1_ASAP7_75t_SL _20245_ (.A1(_11877_),
    .A2(_11517_),
    .B(_11463_),
    .Y(_12018_));
 AO21x1_ASAP7_75t_SL _20246_ (.A1(_11562_),
    .A2(_11850_),
    .B(_11463_),
    .Y(_12019_));
 NAND3x1_ASAP7_75t_SL _20247_ (.A(_12018_),
    .B(_12019_),
    .C(_11493_),
    .Y(_12020_));
 AND3x1_ASAP7_75t_SL _20248_ (.A(_11463_),
    .B(_11449_),
    .C(_11446_),
    .Y(_12021_));
 AO21x1_ASAP7_75t_SL _20249_ (.A1(_01082_),
    .A2(_11463_),
    .B(_11493_),
    .Y(_12022_));
 NOR2x1_ASAP7_75t_SL _20250_ (.A(_12021_),
    .B(_12022_),
    .Y(_12023_));
 AOI21x1_ASAP7_75t_SL _20251_ (.A1(_11803_),
    .A2(_12023_),
    .B(_11512_),
    .Y(_12024_));
 NAND2x1_ASAP7_75t_SL _20252_ (.A(_12024_),
    .B(_12020_),
    .Y(_12025_));
 AO21x1_ASAP7_75t_SL _20253_ (.A1(_01091_),
    .A2(_11470_),
    .B(_11489_),
    .Y(_12026_));
 NOR2x1_ASAP7_75t_SL _20254_ (.A(_11470_),
    .B(_11714_),
    .Y(_12027_));
 OA21x2_ASAP7_75t_SL _20255_ (.A1(_12026_),
    .A2(_12027_),
    .B(_11512_),
    .Y(_12028_));
 NOR2x1_ASAP7_75t_SL _20256_ (.A(_11953_),
    .B(_12022_),
    .Y(_12029_));
 NAND2x1_ASAP7_75t_SL _20257_ (.A(_11703_),
    .B(_12029_),
    .Y(_12030_));
 AOI21x1_ASAP7_75t_SL _20258_ (.A1(_12028_),
    .A2(_12030_),
    .B(_11648_),
    .Y(_12031_));
 AOI21x1_ASAP7_75t_SL _20259_ (.A1(_12031_),
    .A2(_12025_),
    .B(_11595_),
    .Y(_12032_));
 NOR2x1_ASAP7_75t_SL _20260_ (.A(_01100_),
    .B(_11463_),
    .Y(_12033_));
 AOI21x1_ASAP7_75t_SL _20261_ (.A1(_11620_),
    .A2(_11903_),
    .B(_11470_),
    .Y(_12034_));
 OAI21x1_ASAP7_75t_SL _20262_ (.A1(_12033_),
    .A2(_12034_),
    .B(_11493_),
    .Y(_12035_));
 OA21x2_ASAP7_75t_SL _20263_ (.A1(_11606_),
    .A2(_11479_),
    .B(_11470_),
    .Y(_12036_));
 NOR2x1_ASAP7_75t_SL _20264_ (.A(_11690_),
    .B(_11466_),
    .Y(_12037_));
 OAI21x1_ASAP7_75t_SL _20265_ (.A1(_12037_),
    .A2(_12036_),
    .B(_11489_),
    .Y(_12038_));
 NAND2x1_ASAP7_75t_SL _20266_ (.A(_12035_),
    .B(_12038_),
    .Y(_12039_));
 AOI21x1_ASAP7_75t_SL _20267_ (.A1(_11512_),
    .A2(_12039_),
    .B(_11549_),
    .Y(_12040_));
 NAND2x1_ASAP7_75t_SL _20268_ (.A(_11751_),
    .B(_11463_),
    .Y(_12041_));
 NAND2x1_ASAP7_75t_SL _20269_ (.A(_11499_),
    .B(_11853_),
    .Y(_12042_));
 AOI21x1_ASAP7_75t_SL _20270_ (.A1(_12041_),
    .A2(_12042_),
    .B(_11493_),
    .Y(_12043_));
 AO21x1_ASAP7_75t_SL _20271_ (.A1(_11683_),
    .A2(_01082_),
    .B(_11877_),
    .Y(_12044_));
 OA21x2_ASAP7_75t_SL _20272_ (.A1(_12044_),
    .A2(_12027_),
    .B(_11493_),
    .Y(_12045_));
 OAI21x1_ASAP7_75t_SL _20273_ (.A1(_12043_),
    .A2(_12045_),
    .B(_11513_),
    .Y(_12046_));
 NAND2x1_ASAP7_75t_SL _20274_ (.A(_12046_),
    .B(_12040_),
    .Y(_12047_));
 NAND2x1_ASAP7_75t_SL _20275_ (.A(_12047_),
    .B(_12032_),
    .Y(_12048_));
 AO21x1_ASAP7_75t_SL _20276_ (.A1(_11626_),
    .A2(_11713_),
    .B(_11463_),
    .Y(_12049_));
 NAND3x1_ASAP7_75t_SL _20277_ (.A(_11821_),
    .B(_11489_),
    .C(_12049_),
    .Y(_12050_));
 INVx1_ASAP7_75t_SL _20278_ (.A(_11983_),
    .Y(_12051_));
 AOI21x1_ASAP7_75t_SL _20279_ (.A1(_11467_),
    .A2(_11853_),
    .B(_11489_),
    .Y(_12052_));
 AOI21x1_ASAP7_75t_SL _20280_ (.A1(_12051_),
    .A2(_12052_),
    .B(_11512_),
    .Y(_12053_));
 NAND2x1_ASAP7_75t_SL _20281_ (.A(_12053_),
    .B(_12050_),
    .Y(_12054_));
 AO21x1_ASAP7_75t_SL _20282_ (.A1(_11463_),
    .A2(_11479_),
    .B(_11489_),
    .Y(_12055_));
 AO21x1_ASAP7_75t_SL _20283_ (.A1(_11470_),
    .A2(_11657_),
    .B(_12055_),
    .Y(_12056_));
 OAI21x1_ASAP7_75t_SL _20284_ (.A1(_11479_),
    .A2(_11517_),
    .B(_11463_),
    .Y(_12057_));
 AOI21x1_ASAP7_75t_SL _20285_ (.A1(_11470_),
    .A2(_11639_),
    .B(_11493_),
    .Y(_12058_));
 AOI21x1_ASAP7_75t_SL _20286_ (.A1(_12057_),
    .A2(_12058_),
    .B(_11513_),
    .Y(_12059_));
 AOI21x1_ASAP7_75t_SL _20287_ (.A1(_12059_),
    .A2(_12056_),
    .B(_11549_),
    .Y(_12060_));
 AOI21x1_ASAP7_75t_SL _20288_ (.A1(_12060_),
    .A2(_12054_),
    .B(_11596_),
    .Y(_12061_));
 AO21x1_ASAP7_75t_SL _20289_ (.A1(_11689_),
    .A2(_11467_),
    .B(_11955_),
    .Y(_12062_));
 AOI21x1_ASAP7_75t_SL _20290_ (.A1(_11489_),
    .A2(_12062_),
    .B(_11513_),
    .Y(_12063_));
 AO21x1_ASAP7_75t_SL _20291_ (.A1(_11518_),
    .A2(_11583_),
    .B(_11470_),
    .Y(_12064_));
 NAND2x1_ASAP7_75t_SL _20292_ (.A(_12064_),
    .B(_11733_),
    .Y(_12065_));
 NAND2x1_ASAP7_75t_SL _20293_ (.A(_12063_),
    .B(_12065_),
    .Y(_12066_));
 AOI21x1_ASAP7_75t_SL _20294_ (.A1(_11863_),
    .A2(_11640_),
    .B(_11904_),
    .Y(_12067_));
 AOI21x1_ASAP7_75t_SL _20295_ (.A1(_11493_),
    .A2(_12067_),
    .B(_11512_),
    .Y(_12068_));
 AO21x1_ASAP7_75t_SL _20296_ (.A1(_11518_),
    .A2(_11563_),
    .B(_11463_),
    .Y(_12069_));
 OA21x2_ASAP7_75t_SL _20297_ (.A1(_11908_),
    .A2(_11466_),
    .B(_11489_),
    .Y(_12070_));
 NAND2x1_ASAP7_75t_SL _20298_ (.A(_12069_),
    .B(_12070_),
    .Y(_12071_));
 AOI21x1_ASAP7_75t_SL _20299_ (.A1(_12068_),
    .A2(_12071_),
    .B(_11648_),
    .Y(_12072_));
 NAND2x1_ASAP7_75t_SL _20300_ (.A(_12066_),
    .B(_12072_),
    .Y(_12073_));
 NAND2x1_ASAP7_75t_SL _20301_ (.A(_12073_),
    .B(_12061_),
    .Y(_12074_));
 NAND2x1_ASAP7_75t_SL _20302_ (.A(_12074_),
    .B(_12048_),
    .Y(_00047_));
 NOR2x1_ASAP7_75t_R _20303_ (.A(_00574_),
    .B(_00450_),
    .Y(_12075_));
 XOR2x2_ASAP7_75t_SL _20304_ (.A(_00630_),
    .B(_00623_),
    .Y(_12076_));
 XOR2x2_ASAP7_75t_R _20305_ (.A(_12076_),
    .B(_00688_),
    .Y(_12077_));
 XOR2x2_ASAP7_75t_SL _20306_ (.A(_00591_),
    .B(_00598_),
    .Y(_12078_));
 XOR2x2_ASAP7_75t_SL _20307_ (.A(_00624_),
    .B(_00656_),
    .Y(_12079_));
 XOR2x2_ASAP7_75t_L _20308_ (.A(_12078_),
    .B(_12079_),
    .Y(_12080_));
 NAND2x1_ASAP7_75t_SL _20309_ (.A(_12077_),
    .B(_12080_),
    .Y(_12081_));
 INVx1_ASAP7_75t_R _20310_ (.A(_00688_),
    .Y(_12082_));
 XOR2x2_ASAP7_75t_L _20311_ (.A(_12076_),
    .B(_12082_),
    .Y(_12083_));
 XNOR2x2_ASAP7_75t_SL _20312_ (.A(_00591_),
    .B(_00598_),
    .Y(_12084_));
 XOR2x2_ASAP7_75t_L _20313_ (.A(_12084_),
    .B(_12079_),
    .Y(_12085_));
 NAND2x1_ASAP7_75t_SL _20314_ (.A(_12083_),
    .B(_12085_),
    .Y(_12086_));
 AOI21x1_ASAP7_75t_R _20315_ (.A1(_12081_),
    .A2(_12086_),
    .B(_10675_),
    .Y(_12087_));
 OAI21x1_ASAP7_75t_R _20316_ (.A1(_12075_),
    .A2(_12087_),
    .B(_00919_),
    .Y(_12088_));
 AND2x2_ASAP7_75t_R _20318_ (.A(_10675_),
    .B(_00450_),
    .Y(_12090_));
 NAND2x1_ASAP7_75t_R _20319_ (.A(_12083_),
    .B(_12080_),
    .Y(_12091_));
 NAND2x1_ASAP7_75t_R _20320_ (.A(_12077_),
    .B(_12085_),
    .Y(_12092_));
 AOI21x1_ASAP7_75t_SL _20321_ (.A1(_12091_),
    .A2(_12092_),
    .B(_10675_),
    .Y(_12093_));
 INVx1_ASAP7_75t_R _20322_ (.A(_00919_),
    .Y(_12094_));
 OAI21x1_ASAP7_75t_R _20323_ (.A1(_12090_),
    .A2(_12093_),
    .B(_12094_),
    .Y(_12095_));
 NAND2x1_ASAP7_75t_SL _20324_ (.A(_12088_),
    .B(_12095_),
    .Y(_12096_));
 INVx1_ASAP7_75t_R _20326_ (.A(_00687_),
    .Y(_12097_));
 XOR2x2_ASAP7_75t_SL _20327_ (.A(_00598_),
    .B(_00630_),
    .Y(_12098_));
 NAND2x1_ASAP7_75t_R _20328_ (.A(_12097_),
    .B(_12098_),
    .Y(_12099_));
 XNOR2x2_ASAP7_75t_SL _20329_ (.A(_00598_),
    .B(_00630_),
    .Y(_12100_));
 NAND2x1_ASAP7_75t_R _20330_ (.A(_00687_),
    .B(_12100_),
    .Y(_12101_));
 XOR2x2_ASAP7_75t_SL _20331_ (.A(_00623_),
    .B(_00655_),
    .Y(_12102_));
 INVx1_ASAP7_75t_R _20332_ (.A(_12102_),
    .Y(_12103_));
 AOI21x1_ASAP7_75t_R _20333_ (.A1(_12099_),
    .A2(_12101_),
    .B(_12103_),
    .Y(_12104_));
 NAND2x1_ASAP7_75t_R _20334_ (.A(_00687_),
    .B(_12098_),
    .Y(_12105_));
 NAND2x1_ASAP7_75t_R _20335_ (.A(_12097_),
    .B(_12100_),
    .Y(_12106_));
 AOI21x1_ASAP7_75t_R _20336_ (.A1(_12105_),
    .A2(_12106_),
    .B(_12102_),
    .Y(_12107_));
 OAI21x1_ASAP7_75t_SL _20337_ (.A1(_12104_),
    .A2(_12107_),
    .B(_00574_),
    .Y(_12108_));
 NOR2x1_ASAP7_75t_R _20338_ (.A(_00574_),
    .B(_00451_),
    .Y(_12109_));
 INVx1_ASAP7_75t_R _20339_ (.A(_12109_),
    .Y(_12110_));
 NAND3x1_ASAP7_75t_R _20340_ (.A(_12108_),
    .B(_08843_),
    .C(_12110_),
    .Y(_12111_));
 INVx1_ASAP7_75t_SL _20341_ (.A(_12108_),
    .Y(_12112_));
 OAI21x1_ASAP7_75t_R _20342_ (.A1(_12109_),
    .A2(_12112_),
    .B(_00918_),
    .Y(_12113_));
 NAND2x1_ASAP7_75t_SL _20343_ (.A(_12111_),
    .B(_12113_),
    .Y(_12114_));
 INVx1_ASAP7_75t_R _20345_ (.A(_00625_),
    .Y(_12115_));
 XOR2x2_ASAP7_75t_SL _20346_ (.A(_00592_),
    .B(_00624_),
    .Y(_12116_));
 NAND2x1_ASAP7_75t_R _20347_ (.A(_12115_),
    .B(_12116_),
    .Y(_12117_));
 XNOR2x2_ASAP7_75t_SL _20348_ (.A(_00624_),
    .B(_00592_),
    .Y(_12118_));
 NAND2x1_ASAP7_75t_R _20349_ (.A(_00625_),
    .B(_12118_),
    .Y(_12119_));
 XNOR2x1_ASAP7_75t_SL _20350_ (.B(_00689_),
    .Y(_12120_),
    .A(_00657_));
 AOI21x1_ASAP7_75t_SL _20351_ (.A1(_12117_),
    .A2(_12119_),
    .B(_12120_),
    .Y(_12121_));
 NAND2x1_ASAP7_75t_R _20352_ (.A(_00625_),
    .B(_12116_),
    .Y(_12122_));
 NAND2x1_ASAP7_75t_SL _20353_ (.A(_12115_),
    .B(_12118_),
    .Y(_12123_));
 XOR2x2_ASAP7_75t_SL _20354_ (.A(_00657_),
    .B(_00689_),
    .Y(_12124_));
 AOI21x1_ASAP7_75t_SL _20355_ (.A1(_12122_),
    .A2(_12123_),
    .B(_12124_),
    .Y(_12125_));
 OAI21x1_ASAP7_75t_SL _20356_ (.A1(_12121_),
    .A2(_12125_),
    .B(_00574_),
    .Y(_12126_));
 OR2x2_ASAP7_75t_SL _20357_ (.A(_00574_),
    .B(_00452_),
    .Y(_12127_));
 NAND3x1_ASAP7_75t_SL _20359_ (.A(_12126_),
    .B(_00920_),
    .C(_12127_),
    .Y(_12129_));
 AOI21x1_ASAP7_75t_SL _20360_ (.A1(_12127_),
    .A2(_12126_),
    .B(_00920_),
    .Y(_12130_));
 INVx3_ASAP7_75t_SL _20361_ (.A(_12130_),
    .Y(_12131_));
 NAND2x2_ASAP7_75t_SL _20362_ (.A(_12129_),
    .B(_12131_),
    .Y(_12132_));
 NAND3x1_ASAP7_75t_L _20365_ (.A(_12108_),
    .B(_00918_),
    .C(_12110_),
    .Y(_12134_));
 OAI21x1_ASAP7_75t_SL _20366_ (.A1(_12109_),
    .A2(_12112_),
    .B(_08843_),
    .Y(_12135_));
 NAND2x2_ASAP7_75t_SL _20367_ (.A(_12134_),
    .B(_12135_),
    .Y(_12136_));
 NAND3x1_ASAP7_75t_SL _20369_ (.A(_12126_),
    .B(_08848_),
    .C(_12127_),
    .Y(_12137_));
 AOI21x1_ASAP7_75t_SL _20370_ (.A1(_12127_),
    .A2(_12126_),
    .B(_08848_),
    .Y(_12138_));
 INVx2_ASAP7_75t_SL _20371_ (.A(_12138_),
    .Y(_12139_));
 NAND2x2_ASAP7_75t_SL _20372_ (.A(_12137_),
    .B(_12139_),
    .Y(_12140_));
 NAND2x1_ASAP7_75t_SL _20374_ (.A(_12114_),
    .B(_12140_),
    .Y(_12141_));
 INVx1_ASAP7_75t_SL _20376_ (.A(_01110_),
    .Y(_12143_));
 AO21x1_ASAP7_75t_R _20377_ (.A1(_12131_),
    .A2(_12129_),
    .B(_12143_),
    .Y(_12144_));
 XOR2x1_ASAP7_75t_SL _20378_ (.A(_00625_),
    .Y(_12145_),
    .B(_00630_));
 XOR2x2_ASAP7_75t_L _20379_ (.A(_00658_),
    .B(_00690_),
    .Y(_12146_));
 XOR2x2_ASAP7_75t_R _20380_ (.A(_12145_),
    .B(_12146_),
    .Y(_12147_));
 XOR2x2_ASAP7_75t_R _20381_ (.A(_00593_),
    .B(_00598_),
    .Y(_12148_));
 XOR2x2_ASAP7_75t_SL _20382_ (.A(_12148_),
    .B(_00626_),
    .Y(_12149_));
 AND2x2_ASAP7_75t_SL _20383_ (.A(_12147_),
    .B(_12149_),
    .Y(_12150_));
 OAI21x1_ASAP7_75t_R _20384_ (.A1(_12149_),
    .A2(_12147_),
    .B(_00574_),
    .Y(_12151_));
 NAND2x1_ASAP7_75t_R _20385_ (.A(_00517_),
    .B(_10675_),
    .Y(_12152_));
 OAI21x1_ASAP7_75t_SL _20386_ (.A1(_12150_),
    .A2(_12151_),
    .B(_12152_),
    .Y(_12153_));
 XOR2x2_ASAP7_75t_SL _20387_ (.A(_12153_),
    .B(_08851_),
    .Y(_12154_));
 AO21x1_ASAP7_75t_SL _20390_ (.A1(_12141_),
    .A2(_12144_),
    .B(_12154_),
    .Y(_12157_));
 XOR2x2_ASAP7_75t_L _20391_ (.A(_00626_),
    .B(_00630_),
    .Y(_12158_));
 XOR2x2_ASAP7_75t_R _20392_ (.A(_00659_),
    .B(_00691_),
    .Y(_12159_));
 XOR2x2_ASAP7_75t_SL _20393_ (.A(_12158_),
    .B(_12159_),
    .Y(_12160_));
 XOR2x2_ASAP7_75t_R _20394_ (.A(_00594_),
    .B(_00598_),
    .Y(_12161_));
 XNOR2x2_ASAP7_75t_R _20395_ (.A(_00627_),
    .B(_12161_),
    .Y(_12162_));
 XOR2x2_ASAP7_75t_SL _20396_ (.A(_12160_),
    .B(_12162_),
    .Y(_12163_));
 NOR2x1_ASAP7_75t_R _20398_ (.A(_00574_),
    .B(_00515_),
    .Y(_12165_));
 AOI21x1_ASAP7_75t_SL _20399_ (.A1(_00574_),
    .A2(_12163_),
    .B(_12165_),
    .Y(_12166_));
 XNOR2x2_ASAP7_75t_SL _20400_ (.A(_00922_),
    .B(_12166_),
    .Y(_12167_));
 INVx1_ASAP7_75t_SL _20402_ (.A(_12129_),
    .Y(_12169_));
 INVx2_ASAP7_75t_R _20404_ (.A(_01105_),
    .Y(_12171_));
 OAI21x1_ASAP7_75t_R _20405_ (.A1(_12130_),
    .A2(_12169_),
    .B(_12171_),
    .Y(_12172_));
 XOR2x2_ASAP7_75t_SL _20406_ (.A(_12153_),
    .B(_00921_),
    .Y(_12173_));
 AOI21x1_ASAP7_75t_SL _20408_ (.A1(_12140_),
    .A2(_12096_),
    .B(_12173_),
    .Y(_12175_));
 NAND2x1_ASAP7_75t_SL _20409_ (.A(_12172_),
    .B(_12175_),
    .Y(_12176_));
 AND3x1_ASAP7_75t_SL _20410_ (.A(_12157_),
    .B(_12167_),
    .C(_12176_),
    .Y(_12177_));
 AOI21x1_ASAP7_75t_SL _20415_ (.A1(_01108_),
    .A2(_12140_),
    .B(_12154_),
    .Y(_12182_));
 INVx1_ASAP7_75t_SL _20416_ (.A(_12182_),
    .Y(_12183_));
 AO21x1_ASAP7_75t_SL _20417_ (.A1(_12139_),
    .A2(_12137_),
    .B(_01106_),
    .Y(_12184_));
 INVx1_ASAP7_75t_SL _20418_ (.A(_01104_),
    .Y(_12185_));
 AO21x1_ASAP7_75t_R _20419_ (.A1(_12131_),
    .A2(_12129_),
    .B(_12185_),
    .Y(_12186_));
 AO21x1_ASAP7_75t_SL _20421_ (.A1(_12184_),
    .A2(_12186_),
    .B(_12173_),
    .Y(_12188_));
 NAND2x1_ASAP7_75t_SL _20422_ (.A(_12183_),
    .B(_12188_),
    .Y(_12189_));
 XOR2x2_ASAP7_75t_SL _20423_ (.A(_00628_),
    .B(_00660_),
    .Y(_12190_));
 XOR2x2_ASAP7_75t_R _20424_ (.A(_12190_),
    .B(_00692_),
    .Y(_12191_));
 XNOR2x2_ASAP7_75t_R _20425_ (.A(_00595_),
    .B(_00627_),
    .Y(_12192_));
 XOR2x2_ASAP7_75t_SL _20426_ (.A(_12191_),
    .B(_12192_),
    .Y(_12193_));
 NOR2x1_ASAP7_75t_R _20427_ (.A(_00574_),
    .B(_00514_),
    .Y(_12194_));
 AO21x1_ASAP7_75t_R _20428_ (.A1(_12193_),
    .A2(_00574_),
    .B(_12194_),
    .Y(_12195_));
 XOR2x2_ASAP7_75t_SL _20429_ (.A(_12195_),
    .B(_00923_),
    .Y(_12196_));
 INVx1_ASAP7_75t_SL _20430_ (.A(_12196_),
    .Y(_12197_));
 OAI21x1_ASAP7_75t_SL _20432_ (.A1(_12167_),
    .A2(_12189_),
    .B(_12197_),
    .Y(_12199_));
 AO21x1_ASAP7_75t_SL _20433_ (.A1(_12131_),
    .A2(_12129_),
    .B(_01108_),
    .Y(_12200_));
 OA21x2_ASAP7_75t_SL _20435_ (.A1(_12200_),
    .A2(_12173_),
    .B(_12167_),
    .Y(_12202_));
 NOR2x1_ASAP7_75t_SL _20436_ (.A(_12114_),
    .B(_12140_),
    .Y(_12203_));
 NOR2x1_ASAP7_75t_SL _20437_ (.A(_12154_),
    .B(_12203_),
    .Y(_12204_));
 OAI21x1_ASAP7_75t_SL _20438_ (.A1(_12075_),
    .A2(_12087_),
    .B(_12094_),
    .Y(_12205_));
 OAI21x1_ASAP7_75t_SL _20439_ (.A1(_12090_),
    .A2(_12093_),
    .B(_00919_),
    .Y(_12206_));
 NAND2x2_ASAP7_75t_SL _20440_ (.A(_12206_),
    .B(_12205_),
    .Y(_01103_));
 NOR2x1_ASAP7_75t_SL _20441_ (.A(_12136_),
    .B(_01103_),
    .Y(_12207_));
 NAND2x1_ASAP7_75t_SL _20442_ (.A(_12140_),
    .B(_12207_),
    .Y(_12208_));
 NAND2x1_ASAP7_75t_SL _20443_ (.A(_12204_),
    .B(_12208_),
    .Y(_12209_));
 NAND2x1_ASAP7_75t_SL _20444_ (.A(_12202_),
    .B(_12209_),
    .Y(_12210_));
 AOI21x1_ASAP7_75t_SL _20445_ (.A1(_12137_),
    .A2(_12139_),
    .B(_12171_),
    .Y(_12211_));
 NOR2x2_ASAP7_75t_SL _20446_ (.A(_12211_),
    .B(_12154_),
    .Y(_12212_));
 NOR2x1_ASAP7_75t_SL _20447_ (.A(_12167_),
    .B(_12212_),
    .Y(_12213_));
 NAND2x1_ASAP7_75t_SL _20448_ (.A(_12127_),
    .B(_12126_),
    .Y(_12214_));
 NOR2x1_ASAP7_75t_SL _20449_ (.A(_00920_),
    .B(_12214_),
    .Y(_12215_));
 INVx1_ASAP7_75t_SL _20450_ (.A(_01111_),
    .Y(_12216_));
 OAI21x1_ASAP7_75t_SL _20451_ (.A1(_12138_),
    .A2(_12215_),
    .B(_12216_),
    .Y(_12217_));
 AO21x1_ASAP7_75t_SL _20453_ (.A1(_12200_),
    .A2(_12217_),
    .B(_12173_),
    .Y(_12219_));
 AOI21x1_ASAP7_75t_SL _20455_ (.A1(_12213_),
    .A2(_12219_),
    .B(_12197_),
    .Y(_12221_));
 XOR2x2_ASAP7_75t_SL _20456_ (.A(_00596_),
    .B(_00628_),
    .Y(_12222_));
 XOR2x2_ASAP7_75t_SL _20457_ (.A(_00629_),
    .B(_00661_),
    .Y(_12223_));
 XOR2x2_ASAP7_75t_R _20458_ (.A(_12223_),
    .B(_00693_),
    .Y(_12224_));
 XNOR2x2_ASAP7_75t_R _20459_ (.A(_12222_),
    .B(_12224_),
    .Y(_12225_));
 NOR2x1_ASAP7_75t_SL _20460_ (.A(_00574_),
    .B(_00513_),
    .Y(_12226_));
 AO21x1_ASAP7_75t_R _20461_ (.A1(_12225_),
    .A2(_00574_),
    .B(_12226_),
    .Y(_12227_));
 XOR2x2_ASAP7_75t_SL _20462_ (.A(_12227_),
    .B(_00925_),
    .Y(_12228_));
 AOI21x1_ASAP7_75t_SL _20464_ (.A1(_12210_),
    .A2(_12221_),
    .B(_12228_),
    .Y(_12230_));
 OAI21x1_ASAP7_75t_SL _20465_ (.A1(_12177_),
    .A2(_12199_),
    .B(_12230_),
    .Y(_12231_));
 NOR2x2_ASAP7_75t_SL _20466_ (.A(_12114_),
    .B(_01103_),
    .Y(_12232_));
 NAND2x1_ASAP7_75t_SL _20467_ (.A(_12140_),
    .B(_12232_),
    .Y(_12233_));
 INVx1_ASAP7_75t_SL _20468_ (.A(_12233_),
    .Y(_12234_));
 AO21x1_ASAP7_75t_SL _20470_ (.A1(_12131_),
    .A2(_12129_),
    .B(_01110_),
    .Y(_12236_));
 NAND2x1_ASAP7_75t_SL _20471_ (.A(_12154_),
    .B(_12236_),
    .Y(_12237_));
 NOR2x1_ASAP7_75t_SL _20473_ (.A(_12154_),
    .B(_12184_),
    .Y(_12239_));
 NOR2x1_ASAP7_75t_SL _20474_ (.A(_12167_),
    .B(_12239_),
    .Y(_12240_));
 OAI21x1_ASAP7_75t_SL _20475_ (.A1(_12234_),
    .A2(_12237_),
    .B(_12240_),
    .Y(_12241_));
 OA21x2_ASAP7_75t_SL _20476_ (.A1(_12184_),
    .A2(_12173_),
    .B(_12167_),
    .Y(_12242_));
 AOI21x1_ASAP7_75t_SL _20477_ (.A1(_01111_),
    .A2(_12132_),
    .B(_12154_),
    .Y(_12243_));
 NAND2x1_ASAP7_75t_SL _20478_ (.A(_12243_),
    .B(_12233_),
    .Y(_12244_));
 AOI21x1_ASAP7_75t_SL _20480_ (.A1(_12242_),
    .A2(_12244_),
    .B(_12196_),
    .Y(_12246_));
 INVx1_ASAP7_75t_SL _20481_ (.A(_12228_),
    .Y(_12247_));
 AOI21x1_ASAP7_75t_SL _20482_ (.A1(_12241_),
    .A2(_12246_),
    .B(_12247_),
    .Y(_12248_));
 NOR2x1_ASAP7_75t_SL _20483_ (.A(_01108_),
    .B(_12140_),
    .Y(_12249_));
 AOI21x1_ASAP7_75t_SL _20484_ (.A1(_12136_),
    .A2(_12096_),
    .B(_12132_),
    .Y(_12250_));
 OAI21x1_ASAP7_75t_SL _20485_ (.A1(_12249_),
    .A2(_12250_),
    .B(_12154_),
    .Y(_12251_));
 INVx1_ASAP7_75t_SL _20486_ (.A(_12251_),
    .Y(_12252_));
 INVx1_ASAP7_75t_R _20487_ (.A(_01106_),
    .Y(_12253_));
 OAI21x1_ASAP7_75t_R _20488_ (.A1(_12130_),
    .A2(_12169_),
    .B(_12253_),
    .Y(_12254_));
 OA21x2_ASAP7_75t_SL _20489_ (.A1(_12254_),
    .A2(_12173_),
    .B(_12167_),
    .Y(_12255_));
 NAND2x2_ASAP7_75t_SL _20490_ (.A(_12114_),
    .B(_12132_),
    .Y(_12256_));
 OAI21x1_ASAP7_75t_SL _20491_ (.A1(_12138_),
    .A2(_12215_),
    .B(_01104_),
    .Y(_12257_));
 AO21x1_ASAP7_75t_SL _20493_ (.A1(_12256_),
    .A2(_12257_),
    .B(_12154_),
    .Y(_12259_));
 NAND2x1_ASAP7_75t_SL _20494_ (.A(_12255_),
    .B(_12259_),
    .Y(_12260_));
 AOI21x1_ASAP7_75t_R _20495_ (.A1(_12129_),
    .A2(_12131_),
    .B(_01105_),
    .Y(_12261_));
 AOI21x1_ASAP7_75t_R _20496_ (.A1(_12154_),
    .A2(_12261_),
    .B(_12167_),
    .Y(_12262_));
 OA21x2_ASAP7_75t_SL _20497_ (.A1(_01118_),
    .A2(_12154_),
    .B(_12262_),
    .Y(_12263_));
 NOR2x1_ASAP7_75t_SL _20498_ (.A(_12197_),
    .B(_12263_),
    .Y(_12264_));
 OAI21x1_ASAP7_75t_SL _20499_ (.A1(_12252_),
    .A2(_12260_),
    .B(_12264_),
    .Y(_12265_));
 NAND2x1_ASAP7_75t_SL _20500_ (.A(_12248_),
    .B(_12265_),
    .Y(_12266_));
 XNOR2x2_ASAP7_75t_R _20501_ (.A(_00597_),
    .B(_00629_),
    .Y(_12267_));
 INVx2_ASAP7_75t_R _20502_ (.A(_00694_),
    .Y(_12268_));
 XOR2x2_ASAP7_75t_R _20503_ (.A(_12267_),
    .B(_12268_),
    .Y(_12269_));
 XNOR2x2_ASAP7_75t_SL _20504_ (.A(_00630_),
    .B(_00662_),
    .Y(_12270_));
 XOR2x2_ASAP7_75t_SL _20505_ (.A(_12269_),
    .B(_12270_),
    .Y(_12271_));
 NOR2x1_ASAP7_75t_SL _20506_ (.A(_00574_),
    .B(_00512_),
    .Y(_12272_));
 AO21x1_ASAP7_75t_SL _20507_ (.A1(_12271_),
    .A2(_00574_),
    .B(_12272_),
    .Y(_12273_));
 XOR2x2_ASAP7_75t_SL _20508_ (.A(_12273_),
    .B(_00926_),
    .Y(_12274_));
 AOI21x1_ASAP7_75t_SL _20510_ (.A1(_12231_),
    .A2(_12266_),
    .B(_12274_),
    .Y(_12276_));
 NAND2x1_ASAP7_75t_SL _20511_ (.A(_12132_),
    .B(_12096_),
    .Y(_12277_));
 NOR2x1_ASAP7_75t_L _20512_ (.A(_12173_),
    .B(_12211_),
    .Y(_12278_));
 OAI21x1_ASAP7_75t_SL _20513_ (.A1(_12136_),
    .A2(_12277_),
    .B(_12278_),
    .Y(_12279_));
 AO21x1_ASAP7_75t_SL _20515_ (.A1(_12139_),
    .A2(_12137_),
    .B(_12143_),
    .Y(_12281_));
 NAND2x1_ASAP7_75t_SL _20516_ (.A(_12281_),
    .B(_12186_),
    .Y(_12282_));
 XOR2x2_ASAP7_75t_SL _20517_ (.A(_12166_),
    .B(_00922_),
    .Y(_12283_));
 AOI21x1_ASAP7_75t_SL _20519_ (.A1(_12173_),
    .A2(_12282_),
    .B(_12283_),
    .Y(_12285_));
 NAND2x1_ASAP7_75t_SL _20520_ (.A(_12279_),
    .B(_12285_),
    .Y(_12286_));
 AOI21x1_ASAP7_75t_R _20521_ (.A1(_12136_),
    .A2(_12096_),
    .B(_12154_),
    .Y(_12287_));
 NAND2x1_ASAP7_75t_SL _20522_ (.A(_12256_),
    .B(_12287_),
    .Y(_12288_));
 NAND2x1_ASAP7_75t_SL _20523_ (.A(_12136_),
    .B(_01103_),
    .Y(_12289_));
 AOI21x1_ASAP7_75t_SL _20524_ (.A1(_12114_),
    .A2(_12140_),
    .B(_12173_),
    .Y(_12290_));
 NAND2x1_ASAP7_75t_SL _20525_ (.A(_12289_),
    .B(_12290_),
    .Y(_12291_));
 NAND3x1_ASAP7_75t_SL _20528_ (.A(_12288_),
    .B(_12291_),
    .C(_12283_),
    .Y(_12294_));
 AOI21x1_ASAP7_75t_SL _20530_ (.A1(_12286_),
    .A2(_12294_),
    .B(_12196_),
    .Y(_12296_));
 AOI21x1_ASAP7_75t_SL _20531_ (.A1(_12137_),
    .A2(_12139_),
    .B(_01105_),
    .Y(_12297_));
 INVx1_ASAP7_75t_SL _20532_ (.A(_12297_),
    .Y(_12298_));
 AO21x1_ASAP7_75t_SL _20533_ (.A1(_12186_),
    .A2(_12298_),
    .B(_12154_),
    .Y(_12299_));
 AO21x1_ASAP7_75t_SL _20534_ (.A1(_12144_),
    .A2(_12257_),
    .B(_12173_),
    .Y(_12300_));
 AOI21x1_ASAP7_75t_SL _20535_ (.A1(_12299_),
    .A2(_12300_),
    .B(_12283_),
    .Y(_12301_));
 AOI21x1_ASAP7_75t_SL _20536_ (.A1(_01105_),
    .A2(_12132_),
    .B(_12154_),
    .Y(_12302_));
 NOR2x1_ASAP7_75t_SL _20537_ (.A(_12167_),
    .B(_12302_),
    .Y(_12303_));
 NOR2x1p5_ASAP7_75t_SL _20538_ (.A(_12173_),
    .B(_12297_),
    .Y(_12304_));
 NAND2x1_ASAP7_75t_SL _20539_ (.A(_12277_),
    .B(_12304_),
    .Y(_12305_));
 AO21x1_ASAP7_75t_SL _20540_ (.A1(_12303_),
    .A2(_12305_),
    .B(_12197_),
    .Y(_12306_));
 OAI21x1_ASAP7_75t_SL _20541_ (.A1(_12301_),
    .A2(_12306_),
    .B(_12228_),
    .Y(_12307_));
 OAI21x1_ASAP7_75t_SL _20542_ (.A1(_12296_),
    .A2(_12307_),
    .B(_12274_),
    .Y(_12308_));
 NAND2x1_ASAP7_75t_SL _20543_ (.A(_12132_),
    .B(_01103_),
    .Y(_12309_));
 AO21x1_ASAP7_75t_SL _20545_ (.A1(_12309_),
    .A2(_12184_),
    .B(_12173_),
    .Y(_12311_));
 NAND3x1_ASAP7_75t_SL _20547_ (.A(_12209_),
    .B(_12311_),
    .C(_12167_),
    .Y(_12313_));
 INVx1_ASAP7_75t_SL _20548_ (.A(_01113_),
    .Y(_12314_));
 AO21x1_ASAP7_75t_R _20549_ (.A1(_12139_),
    .A2(_12137_),
    .B(_12314_),
    .Y(_12315_));
 AOI21x1_ASAP7_75t_SL _20550_ (.A1(_12315_),
    .A2(_12204_),
    .B(_12167_),
    .Y(_12316_));
 NOR2x1_ASAP7_75t_SL _20551_ (.A(_12132_),
    .B(_01103_),
    .Y(_12317_));
 NAND2x1_ASAP7_75t_SL _20552_ (.A(_12256_),
    .B(_12309_),
    .Y(_12318_));
 OAI21x1_ASAP7_75t_SL _20553_ (.A1(_12317_),
    .A2(_12318_),
    .B(_12154_),
    .Y(_12319_));
 AOI21x1_ASAP7_75t_SL _20554_ (.A1(_12316_),
    .A2(_12319_),
    .B(_12197_),
    .Y(_12320_));
 NAND2x1_ASAP7_75t_SL _20555_ (.A(_12313_),
    .B(_12320_),
    .Y(_12321_));
 NOR2x2_ASAP7_75t_SL _20556_ (.A(_12114_),
    .B(_12132_),
    .Y(_12322_));
 NAND2x1_ASAP7_75t_SL _20557_ (.A(_12136_),
    .B(_12132_),
    .Y(_12323_));
 OAI21x1_ASAP7_75t_SL _20558_ (.A1(_01103_),
    .A2(_12323_),
    .B(_12154_),
    .Y(_12324_));
 NOR2x1_ASAP7_75t_SL _20559_ (.A(_12322_),
    .B(_12324_),
    .Y(_12325_));
 AO21x1_ASAP7_75t_R _20560_ (.A1(_12131_),
    .A2(_12129_),
    .B(_12314_),
    .Y(_12326_));
 AO21x1_ASAP7_75t_SL _20562_ (.A1(_12212_),
    .A2(_12326_),
    .B(_12167_),
    .Y(_12328_));
 NAND2x1_ASAP7_75t_R _20563_ (.A(_12132_),
    .B(_12232_),
    .Y(_12329_));
 NAND2x1_ASAP7_75t_SL _20564_ (.A(_12182_),
    .B(_12329_),
    .Y(_12330_));
 AO21x1_ASAP7_75t_SL _20565_ (.A1(_12132_),
    .A2(_12136_),
    .B(_12173_),
    .Y(_12331_));
 AND2x2_ASAP7_75t_SL _20566_ (.A(_12331_),
    .B(_12167_),
    .Y(_12332_));
 AOI21x1_ASAP7_75t_SL _20567_ (.A1(_12330_),
    .A2(_12332_),
    .B(_12196_),
    .Y(_12333_));
 OAI21x1_ASAP7_75t_SL _20568_ (.A1(_12325_),
    .A2(_12328_),
    .B(_12333_),
    .Y(_12334_));
 AOI21x1_ASAP7_75t_SL _20570_ (.A1(_12321_),
    .A2(_12334_),
    .B(_12228_),
    .Y(_12336_));
 NOR2x1_ASAP7_75t_SL _20571_ (.A(_12308_),
    .B(_12336_),
    .Y(_12337_));
 NOR2x1_ASAP7_75t_SL _20572_ (.A(_12276_),
    .B(_12337_),
    .Y(_00048_));
 INVx1_ASAP7_75t_SL _20574_ (.A(_12144_),
    .Y(_12339_));
 AOI21x1_ASAP7_75t_SL _20575_ (.A1(_12114_),
    .A2(_12096_),
    .B(_12132_),
    .Y(_12340_));
 OAI21x1_ASAP7_75t_SL _20576_ (.A1(_12339_),
    .A2(_12340_),
    .B(_12154_),
    .Y(_12341_));
 NAND2x1_ASAP7_75t_SL _20577_ (.A(_01120_),
    .B(_12173_),
    .Y(_12342_));
 AO21x1_ASAP7_75t_SL _20578_ (.A1(_12167_),
    .A2(_12342_),
    .B(_12197_),
    .Y(_12343_));
 OA21x2_ASAP7_75t_SL _20579_ (.A1(_12283_),
    .A2(_12341_),
    .B(_12343_),
    .Y(_12344_));
 OAI21x1_ASAP7_75t_SL _20581_ (.A1(_12340_),
    .A2(_12318_),
    .B(_12173_),
    .Y(_12346_));
 AO21x1_ASAP7_75t_SL _20582_ (.A1(_12141_),
    .A2(_12186_),
    .B(_12173_),
    .Y(_12347_));
 AO21x1_ASAP7_75t_SL _20583_ (.A1(_12346_),
    .A2(_12347_),
    .B(_12167_),
    .Y(_12348_));
 AO21x1_ASAP7_75t_SL _20584_ (.A1(_12182_),
    .A2(_12309_),
    .B(_12167_),
    .Y(_12349_));
 AO21x1_ASAP7_75t_SL _20585_ (.A1(_12290_),
    .A2(_12277_),
    .B(_12197_),
    .Y(_12350_));
 OAI21x1_ASAP7_75t_SL _20586_ (.A1(_12349_),
    .A2(_12350_),
    .B(_12228_),
    .Y(_12351_));
 AOI21x1_ASAP7_75t_SL _20587_ (.A1(_12344_),
    .A2(_12348_),
    .B(_12351_),
    .Y(_12352_));
 NAND2x1_ASAP7_75t_SL _20588_ (.A(_12309_),
    .B(_12182_),
    .Y(_12353_));
 NOR2x1_ASAP7_75t_SL _20589_ (.A(_12185_),
    .B(_12140_),
    .Y(_12354_));
 OAI21x1_ASAP7_75t_SL _20591_ (.A1(_12354_),
    .A2(_12322_),
    .B(_12154_),
    .Y(_12356_));
 AOI21x1_ASAP7_75t_SL _20593_ (.A1(_12353_),
    .A2(_12356_),
    .B(_12283_),
    .Y(_12358_));
 AO21x1_ASAP7_75t_SL _20594_ (.A1(_12172_),
    .A2(_12257_),
    .B(_12154_),
    .Y(_12359_));
 NOR2x1_ASAP7_75t_SL _20595_ (.A(_12136_),
    .B(_12140_),
    .Y(_12360_));
 INVx1_ASAP7_75t_SL _20596_ (.A(_12184_),
    .Y(_12361_));
 OAI21x1_ASAP7_75t_SL _20597_ (.A1(_12360_),
    .A2(_12361_),
    .B(_12154_),
    .Y(_12362_));
 AOI21x1_ASAP7_75t_SL _20598_ (.A1(_12359_),
    .A2(_12362_),
    .B(_12167_),
    .Y(_12363_));
 OAI21x1_ASAP7_75t_SL _20599_ (.A1(_12358_),
    .A2(_12363_),
    .B(_12197_),
    .Y(_12364_));
 AO21x1_ASAP7_75t_SL _20600_ (.A1(_12131_),
    .A2(_12129_),
    .B(_12253_),
    .Y(_12365_));
 AOI21x1_ASAP7_75t_SL _20601_ (.A1(_01113_),
    .A2(_12140_),
    .B(_12173_),
    .Y(_12366_));
 AOI21x1_ASAP7_75t_SL _20602_ (.A1(_12365_),
    .A2(_12366_),
    .B(_12167_),
    .Y(_12367_));
 NAND2x1_ASAP7_75t_SL _20603_ (.A(_12323_),
    .B(_12309_),
    .Y(_12368_));
 OAI21x1_ASAP7_75t_SL _20604_ (.A1(_12211_),
    .A2(_12368_),
    .B(_12173_),
    .Y(_12369_));
 NAND2x1_ASAP7_75t_SL _20605_ (.A(_12367_),
    .B(_12369_),
    .Y(_12370_));
 NOR2x1_ASAP7_75t_SL _20606_ (.A(_12283_),
    .B(_12212_),
    .Y(_12371_));
 INVx1_ASAP7_75t_SL _20607_ (.A(_12331_),
    .Y(_12372_));
 NAND2x1_ASAP7_75t_SL _20608_ (.A(_12208_),
    .B(_12372_),
    .Y(_12373_));
 AOI21x1_ASAP7_75t_SL _20610_ (.A1(_12371_),
    .A2(_12373_),
    .B(_12197_),
    .Y(_12375_));
 NAND2x1_ASAP7_75t_SL _20611_ (.A(_12370_),
    .B(_12375_),
    .Y(_12376_));
 AOI21x1_ASAP7_75t_SL _20612_ (.A1(_12364_),
    .A2(_12376_),
    .B(_12228_),
    .Y(_12377_));
 OAI21x1_ASAP7_75t_SL _20613_ (.A1(_12352_),
    .A2(_12377_),
    .B(_12274_),
    .Y(_12378_));
 NAND2x1_ASAP7_75t_SL _20614_ (.A(_12154_),
    .B(_12340_),
    .Y(_12379_));
 NAND2x1_ASAP7_75t_SL _20615_ (.A(_12140_),
    .B(_01103_),
    .Y(_12380_));
 AOI21x1_ASAP7_75t_SL _20616_ (.A1(_01113_),
    .A2(_12132_),
    .B(_12154_),
    .Y(_12381_));
 NAND2x1_ASAP7_75t_SL _20617_ (.A(_12380_),
    .B(_12381_),
    .Y(_12382_));
 NAND3x1_ASAP7_75t_SL _20618_ (.A(_12379_),
    .B(_12382_),
    .C(_12283_),
    .Y(_12383_));
 AO21x1_ASAP7_75t_SL _20619_ (.A1(_12139_),
    .A2(_12137_),
    .B(_01108_),
    .Y(_12384_));
 OA21x2_ASAP7_75t_SL _20620_ (.A1(_12384_),
    .A2(_12173_),
    .B(_12167_),
    .Y(_12385_));
 AOI21x1_ASAP7_75t_SL _20621_ (.A1(_12385_),
    .A2(_12369_),
    .B(_12228_),
    .Y(_12386_));
 NAND2x1_ASAP7_75t_SL _20622_ (.A(_12383_),
    .B(_12386_),
    .Y(_12387_));
 INVx2_ASAP7_75t_SL _20623_ (.A(_12212_),
    .Y(_12388_));
 AOI21x1_ASAP7_75t_SL _20624_ (.A1(_01108_),
    .A2(_12140_),
    .B(_12173_),
    .Y(_12389_));
 AOI21x1_ASAP7_75t_SL _20626_ (.A1(_12256_),
    .A2(_12389_),
    .B(_12167_),
    .Y(_12391_));
 OAI21x1_ASAP7_75t_SL _20627_ (.A1(_12203_),
    .A2(_12388_),
    .B(_12391_),
    .Y(_12392_));
 NAND2x1_ASAP7_75t_SL _20628_ (.A(_12289_),
    .B(_12175_),
    .Y(_12393_));
 NAND2x1_ASAP7_75t_SL _20629_ (.A(_12132_),
    .B(_12173_),
    .Y(_12394_));
 OA21x2_ASAP7_75t_SL _20630_ (.A1(_12232_),
    .A2(_12394_),
    .B(_12167_),
    .Y(_12395_));
 AOI21x1_ASAP7_75t_SL _20631_ (.A1(_12393_),
    .A2(_12395_),
    .B(_12247_),
    .Y(_12396_));
 AOI21x1_ASAP7_75t_SL _20633_ (.A1(_12392_),
    .A2(_12396_),
    .B(_12196_),
    .Y(_12398_));
 AOI21x1_ASAP7_75t_SL _20634_ (.A1(_12387_),
    .A2(_12398_),
    .B(_12274_),
    .Y(_12399_));
 NAND2x1_ASAP7_75t_SL _20635_ (.A(_12315_),
    .B(_12302_),
    .Y(_12400_));
 NAND3x1_ASAP7_75t_SL _20636_ (.A(_12251_),
    .B(_12167_),
    .C(_12400_),
    .Y(_12401_));
 AO21x1_ASAP7_75t_SL _20637_ (.A1(_12096_),
    .A2(_12132_),
    .B(_12154_),
    .Y(_12402_));
 NAND2x1_ASAP7_75t_SL _20638_ (.A(_12380_),
    .B(_12402_),
    .Y(_12403_));
 AO21x1_ASAP7_75t_SL _20639_ (.A1(_12249_),
    .A2(_12154_),
    .B(_12167_),
    .Y(_12404_));
 OA21x2_ASAP7_75t_SL _20640_ (.A1(_12403_),
    .A2(_12404_),
    .B(_12228_),
    .Y(_12405_));
 AOI21x1_ASAP7_75t_SL _20641_ (.A1(_12401_),
    .A2(_12405_),
    .B(_12197_),
    .Y(_12406_));
 NAND2x1_ASAP7_75t_SL _20642_ (.A(_12257_),
    .B(_12256_),
    .Y(_12407_));
 OAI22x1_ASAP7_75t_SL _20643_ (.A1(_12407_),
    .A2(_12173_),
    .B1(_12388_),
    .B2(_12249_),
    .Y(_12408_));
 AOI21x1_ASAP7_75t_SL _20644_ (.A1(_12283_),
    .A2(_12408_),
    .B(_12228_),
    .Y(_12409_));
 OA21x2_ASAP7_75t_SL _20645_ (.A1(_12207_),
    .A2(_12322_),
    .B(_12173_),
    .Y(_12410_));
 NAND2x1_ASAP7_75t_SL _20646_ (.A(_12154_),
    .B(_12172_),
    .Y(_12411_));
 NOR2x1_ASAP7_75t_SL _20647_ (.A(_12322_),
    .B(_12411_),
    .Y(_12412_));
 OR3x1_ASAP7_75t_SL _20648_ (.A(_12410_),
    .B(_12283_),
    .C(_12412_),
    .Y(_12413_));
 NAND2x1_ASAP7_75t_SL _20649_ (.A(_12409_),
    .B(_12413_),
    .Y(_12414_));
 NAND2x1_ASAP7_75t_SL _20650_ (.A(_12406_),
    .B(_12414_),
    .Y(_12415_));
 NAND2x1_ASAP7_75t_SL _20651_ (.A(_12399_),
    .B(_12415_),
    .Y(_12416_));
 NAND2x1_ASAP7_75t_SL _20652_ (.A(_12378_),
    .B(_12416_),
    .Y(_00049_));
 NOR2x2_ASAP7_75t_SL _20653_ (.A(_12140_),
    .B(_12154_),
    .Y(_12417_));
 NOR2x1_ASAP7_75t_R _20654_ (.A(_12154_),
    .B(_12096_),
    .Y(_12418_));
 INVx1_ASAP7_75t_SL _20655_ (.A(_12232_),
    .Y(_12419_));
 OAI21x1_ASAP7_75t_SL _20656_ (.A1(_12417_),
    .A2(_12418_),
    .B(_12419_),
    .Y(_12420_));
 NAND2x1_ASAP7_75t_SL _20657_ (.A(_12326_),
    .B(_12389_),
    .Y(_12421_));
 AO21x1_ASAP7_75t_SL _20658_ (.A1(_12420_),
    .A2(_12421_),
    .B(_12167_),
    .Y(_12422_));
 NOR2x1_ASAP7_75t_SL _20659_ (.A(_12249_),
    .B(_12250_),
    .Y(_12423_));
 AOI21x1_ASAP7_75t_SL _20660_ (.A1(_12173_),
    .A2(_12423_),
    .B(_12283_),
    .Y(_12424_));
 NAND2x1_ASAP7_75t_SL _20661_ (.A(_12176_),
    .B(_12424_),
    .Y(_12425_));
 AOI21x1_ASAP7_75t_SL _20662_ (.A1(_12422_),
    .A2(_12425_),
    .B(_12197_),
    .Y(_12426_));
 NOR2x1_ASAP7_75t_SL _20663_ (.A(_12136_),
    .B(_12132_),
    .Y(_12427_));
 NAND2x1_ASAP7_75t_R _20664_ (.A(_12173_),
    .B(_12254_),
    .Y(_12428_));
 INVx1_ASAP7_75t_R _20665_ (.A(_12304_),
    .Y(_12429_));
 INVx1_ASAP7_75t_SL _20666_ (.A(_12309_),
    .Y(_12430_));
 OA22x2_ASAP7_75t_SL _20667_ (.A1(_12427_),
    .A2(_12428_),
    .B1(_12429_),
    .B2(_12430_),
    .Y(_12431_));
 NOR2x1_ASAP7_75t_SL _20668_ (.A(_12167_),
    .B(_12431_),
    .Y(_12432_));
 NAND2x1_ASAP7_75t_SL _20669_ (.A(_12167_),
    .B(_12324_),
    .Y(_12433_));
 OA211x2_ASAP7_75t_SL _20670_ (.A1(_12277_),
    .A2(_12136_),
    .B(_12315_),
    .C(_12173_),
    .Y(_12434_));
 OAI21x1_ASAP7_75t_SL _20671_ (.A1(_12433_),
    .A2(_12434_),
    .B(_12197_),
    .Y(_12435_));
 OAI21x1_ASAP7_75t_SL _20672_ (.A1(_12432_),
    .A2(_12435_),
    .B(_12228_),
    .Y(_12436_));
 NOR2x1_ASAP7_75t_SL _20673_ (.A(_12426_),
    .B(_12436_),
    .Y(_12437_));
 AO21x1_ASAP7_75t_SL _20674_ (.A1(_12141_),
    .A2(_12200_),
    .B(_12154_),
    .Y(_12438_));
 AO21x1_ASAP7_75t_R _20675_ (.A1(_12131_),
    .A2(_12129_),
    .B(_01113_),
    .Y(_12439_));
 AO21x1_ASAP7_75t_SL _20676_ (.A1(_12439_),
    .A2(_12217_),
    .B(_12173_),
    .Y(_12440_));
 AO21x1_ASAP7_75t_SL _20677_ (.A1(_12438_),
    .A2(_12440_),
    .B(_12167_),
    .Y(_12441_));
 NAND2x1_ASAP7_75t_SL _20678_ (.A(_12140_),
    .B(_12096_),
    .Y(_12442_));
 AO21x1_ASAP7_75t_SL _20679_ (.A1(_12442_),
    .A2(_12200_),
    .B(_12154_),
    .Y(_12443_));
 AO21x1_ASAP7_75t_SL _20680_ (.A1(_12443_),
    .A2(_12219_),
    .B(_12283_),
    .Y(_12444_));
 AOI21x1_ASAP7_75t_SL _20681_ (.A1(_12441_),
    .A2(_12444_),
    .B(_12197_),
    .Y(_12445_));
 NAND2x1_ASAP7_75t_R _20683_ (.A(_12172_),
    .B(_12212_),
    .Y(_12447_));
 INVx1_ASAP7_75t_SL _20684_ (.A(_12322_),
    .Y(_12448_));
 AOI21x1_ASAP7_75t_SL _20685_ (.A1(_01111_),
    .A2(_12132_),
    .B(_12173_),
    .Y(_12449_));
 NAND2x1_ASAP7_75t_SL _20686_ (.A(_12448_),
    .B(_12449_),
    .Y(_12450_));
 AOI21x1_ASAP7_75t_SL _20687_ (.A1(_12447_),
    .A2(_12450_),
    .B(_12283_),
    .Y(_12451_));
 NAND2x1_ASAP7_75t_SL _20688_ (.A(_12173_),
    .B(_12217_),
    .Y(_12452_));
 NOR2x1_ASAP7_75t_SL _20689_ (.A(_12430_),
    .B(_12452_),
    .Y(_12453_));
 NAND2x1_ASAP7_75t_R _20690_ (.A(_12154_),
    .B(_12439_),
    .Y(_12454_));
 OAI21x1_ASAP7_75t_SL _20691_ (.A1(_12427_),
    .A2(_12454_),
    .B(_12283_),
    .Y(_12455_));
 NOR2x1_ASAP7_75t_SL _20692_ (.A(_12453_),
    .B(_12455_),
    .Y(_12456_));
 OAI21x1_ASAP7_75t_SL _20693_ (.A1(_12451_),
    .A2(_12456_),
    .B(_12197_),
    .Y(_12457_));
 NAND2x1_ASAP7_75t_SL _20694_ (.A(_12247_),
    .B(_12457_),
    .Y(_12458_));
 OAI21x1_ASAP7_75t_SL _20695_ (.A1(_12445_),
    .A2(_12458_),
    .B(_12274_),
    .Y(_12459_));
 AO21x1_ASAP7_75t_SL _20696_ (.A1(_12200_),
    .A2(_12298_),
    .B(_12154_),
    .Y(_12460_));
 OA21x2_ASAP7_75t_SL _20697_ (.A1(_12257_),
    .A2(_12173_),
    .B(_12167_),
    .Y(_12461_));
 AO21x1_ASAP7_75t_SL _20698_ (.A1(_12460_),
    .A2(_12461_),
    .B(_12196_),
    .Y(_12462_));
 AND2x2_ASAP7_75t_R _20699_ (.A(_01108_),
    .B(_01106_),
    .Y(_12463_));
 NOR2x1_ASAP7_75t_SL _20700_ (.A(_12463_),
    .B(_12132_),
    .Y(_12464_));
 OAI21x1_ASAP7_75t_SL _20701_ (.A1(_12464_),
    .A2(_12368_),
    .B(_12173_),
    .Y(_12465_));
 AND3x1_ASAP7_75t_SL _20702_ (.A(_12465_),
    .B(_12283_),
    .C(_12341_),
    .Y(_12466_));
 NAND2x1_ASAP7_75t_SL _20703_ (.A(_01117_),
    .B(_12173_),
    .Y(_12467_));
 NAND3x1_ASAP7_75t_SL _20704_ (.A(_12324_),
    .B(_12167_),
    .C(_12467_),
    .Y(_12468_));
 OA21x2_ASAP7_75t_SL _20705_ (.A1(_01122_),
    .A2(_12173_),
    .B(_12283_),
    .Y(_12469_));
 AOI21x1_ASAP7_75t_SL _20706_ (.A1(_12469_),
    .A2(_12420_),
    .B(_12197_),
    .Y(_12470_));
 AOI21x1_ASAP7_75t_SL _20707_ (.A1(_12468_),
    .A2(_12470_),
    .B(_12247_),
    .Y(_12471_));
 OAI21x1_ASAP7_75t_SL _20708_ (.A1(_12462_),
    .A2(_12466_),
    .B(_12471_),
    .Y(_12472_));
 NAND2x1_ASAP7_75t_SL _20709_ (.A(_01120_),
    .B(_12154_),
    .Y(_12473_));
 AOI21x1_ASAP7_75t_SL _20710_ (.A1(_12136_),
    .A2(_01103_),
    .B(_12154_),
    .Y(_12474_));
 AOI21x1_ASAP7_75t_SL _20711_ (.A1(_12442_),
    .A2(_12474_),
    .B(_12283_),
    .Y(_12475_));
 AOI21x1_ASAP7_75t_SL _20712_ (.A1(_12473_),
    .A2(_12475_),
    .B(_12197_),
    .Y(_12476_));
 AND2x2_ASAP7_75t_SL _20713_ (.A(_12175_),
    .B(_12186_),
    .Y(_12477_));
 AND3x1_ASAP7_75t_SL _20714_ (.A(_12281_),
    .B(_12173_),
    .C(_12172_),
    .Y(_12478_));
 OAI21x1_ASAP7_75t_SL _20715_ (.A1(_12477_),
    .A2(_12478_),
    .B(_12283_),
    .Y(_12479_));
 NAND2x1_ASAP7_75t_SL _20716_ (.A(_12476_),
    .B(_12479_),
    .Y(_12480_));
 AOI21x1_ASAP7_75t_SL _20717_ (.A1(_12132_),
    .A2(_01103_),
    .B(_12154_),
    .Y(_12481_));
 NAND2x1_ASAP7_75t_SL _20718_ (.A(_12448_),
    .B(_12481_),
    .Y(_12482_));
 NAND3x1_ASAP7_75t_SL _20719_ (.A(_12176_),
    .B(_12482_),
    .C(_12283_),
    .Y(_12483_));
 OA21x2_ASAP7_75t_SL _20720_ (.A1(_01118_),
    .A2(_12173_),
    .B(_12167_),
    .Y(_12484_));
 NAND2x1_ASAP7_75t_SL _20721_ (.A(_12302_),
    .B(_12233_),
    .Y(_12485_));
 AOI21x1_ASAP7_75t_SL _20722_ (.A1(_12484_),
    .A2(_12485_),
    .B(_12196_),
    .Y(_12486_));
 AOI21x1_ASAP7_75t_SL _20723_ (.A1(_12483_),
    .A2(_12486_),
    .B(_12228_),
    .Y(_12487_));
 AOI21x1_ASAP7_75t_SL _20724_ (.A1(_12480_),
    .A2(_12487_),
    .B(_12274_),
    .Y(_12488_));
 NAND2x1_ASAP7_75t_SL _20725_ (.A(_12472_),
    .B(_12488_),
    .Y(_12489_));
 OAI21x1_ASAP7_75t_SL _20726_ (.A1(_12437_),
    .A2(_12459_),
    .B(_12489_),
    .Y(_00050_));
 AO21x1_ASAP7_75t_SL _20727_ (.A1(_12277_),
    .A2(_12141_),
    .B(_12173_),
    .Y(_12490_));
 NAND2x1_ASAP7_75t_SL _20728_ (.A(_12303_),
    .B(_12490_),
    .Y(_12491_));
 NAND2x1_ASAP7_75t_SL _20729_ (.A(_12290_),
    .B(_12419_),
    .Y(_12492_));
 AOI21x1_ASAP7_75t_SL _20730_ (.A1(_12309_),
    .A2(_12212_),
    .B(_12283_),
    .Y(_12493_));
 AOI21x1_ASAP7_75t_SL _20731_ (.A1(_12492_),
    .A2(_12493_),
    .B(_12197_),
    .Y(_12494_));
 NAND2x1_ASAP7_75t_SL _20732_ (.A(_12491_),
    .B(_12494_),
    .Y(_12495_));
 OAI21x1_ASAP7_75t_SL _20733_ (.A1(_12138_),
    .A2(_12215_),
    .B(_12314_),
    .Y(_12496_));
 AO21x1_ASAP7_75t_SL _20734_ (.A1(_12200_),
    .A2(_12496_),
    .B(_12154_),
    .Y(_12497_));
 AOI21x1_ASAP7_75t_SL _20735_ (.A1(_12309_),
    .A2(_12304_),
    .B(_12283_),
    .Y(_12498_));
 AOI21x1_ASAP7_75t_SL _20736_ (.A1(_12497_),
    .A2(_12498_),
    .B(_12196_),
    .Y(_12499_));
 AND2x2_ASAP7_75t_SL _20737_ (.A(_12302_),
    .B(_12257_),
    .Y(_12500_));
 NAND2x1_ASAP7_75t_SL _20738_ (.A(_12281_),
    .B(_12256_),
    .Y(_12501_));
 NOR2x1_ASAP7_75t_SL _20739_ (.A(_12173_),
    .B(_12501_),
    .Y(_12502_));
 OAI21x1_ASAP7_75t_SL _20740_ (.A1(_12500_),
    .A2(_12502_),
    .B(_12283_),
    .Y(_12503_));
 NAND2x1_ASAP7_75t_SL _20741_ (.A(_12499_),
    .B(_12503_),
    .Y(_12504_));
 AOI21x1_ASAP7_75t_SL _20742_ (.A1(_12495_),
    .A2(_12504_),
    .B(_12247_),
    .Y(_12505_));
 NAND2x1_ASAP7_75t_SL _20743_ (.A(_12140_),
    .B(_12173_),
    .Y(_12506_));
 AND2x2_ASAP7_75t_SL _20744_ (.A(_12289_),
    .B(_12256_),
    .Y(_12507_));
 AOI21x1_ASAP7_75t_SL _20745_ (.A1(_12506_),
    .A2(_12507_),
    .B(_12283_),
    .Y(_12508_));
 OAI21x1_ASAP7_75t_SL _20746_ (.A1(_12216_),
    .A2(_12140_),
    .B(_12304_),
    .Y(_12509_));
 AOI21x1_ASAP7_75t_SL _20747_ (.A1(_12382_),
    .A2(_12509_),
    .B(_12167_),
    .Y(_12510_));
 OAI21x1_ASAP7_75t_SL _20748_ (.A1(_12508_),
    .A2(_12510_),
    .B(_12196_),
    .Y(_12511_));
 INVx1_ASAP7_75t_SL _20749_ (.A(_12481_),
    .Y(_12512_));
 NOR2x1_ASAP7_75t_SL _20750_ (.A(_12512_),
    .B(_12501_),
    .Y(_12513_));
 OAI21x1_ASAP7_75t_SL _20751_ (.A1(_12340_),
    .A2(_12411_),
    .B(_12167_),
    .Y(_12514_));
 NOR2x1_ASAP7_75t_SL _20752_ (.A(_12513_),
    .B(_12514_),
    .Y(_12515_));
 AOI21x1_ASAP7_75t_SL _20753_ (.A1(_12144_),
    .A2(_12278_),
    .B(_12167_),
    .Y(_12516_));
 AND2x2_ASAP7_75t_SL _20754_ (.A(_12516_),
    .B(_12288_),
    .Y(_12517_));
 OAI21x1_ASAP7_75t_SL _20755_ (.A1(_12515_),
    .A2(_12517_),
    .B(_12197_),
    .Y(_12518_));
 AOI21x1_ASAP7_75t_SL _20756_ (.A1(_12511_),
    .A2(_12518_),
    .B(_12228_),
    .Y(_12519_));
 INVx1_ASAP7_75t_SL _20757_ (.A(_12274_),
    .Y(_12520_));
 OAI21x1_ASAP7_75t_SL _20758_ (.A1(_12505_),
    .A2(_12519_),
    .B(_12520_),
    .Y(_12521_));
 NAND2x1_ASAP7_75t_SL _20759_ (.A(_01105_),
    .B(_12417_),
    .Y(_12522_));
 NAND2x1_ASAP7_75t_SL _20760_ (.A(_12236_),
    .B(_12175_),
    .Y(_12523_));
 AOI21x1_ASAP7_75t_SL _20761_ (.A1(_12522_),
    .A2(_12523_),
    .B(_12197_),
    .Y(_12524_));
 NAND2x1_ASAP7_75t_SL _20762_ (.A(_12154_),
    .B(_12211_),
    .Y(_12525_));
 OAI21x1_ASAP7_75t_SL _20763_ (.A1(_12196_),
    .A2(_12525_),
    .B(_12240_),
    .Y(_12526_));
 OAI21x1_ASAP7_75t_SL _20764_ (.A1(_12524_),
    .A2(_12526_),
    .B(_12228_),
    .Y(_12527_));
 NOR2x1_ASAP7_75t_SL _20765_ (.A(_12154_),
    .B(_12217_),
    .Y(_12528_));
 AOI21x1_ASAP7_75t_SL _20766_ (.A1(_12448_),
    .A2(_12449_),
    .B(_12528_),
    .Y(_12529_));
 OAI21x1_ASAP7_75t_SL _20767_ (.A1(_12196_),
    .A2(_12529_),
    .B(_12167_),
    .Y(_12530_));
 OAI21x1_ASAP7_75t_SL _20768_ (.A1(_12297_),
    .A2(_12360_),
    .B(_12154_),
    .Y(_12531_));
 INVx1_ASAP7_75t_SL _20769_ (.A(_12464_),
    .Y(_12532_));
 AO21x1_ASAP7_75t_SL _20770_ (.A1(_12532_),
    .A2(_12439_),
    .B(_12154_),
    .Y(_12533_));
 AOI21x1_ASAP7_75t_SL _20771_ (.A1(_12531_),
    .A2(_12533_),
    .B(_12197_),
    .Y(_12534_));
 NOR2x1_ASAP7_75t_SL _20772_ (.A(_12530_),
    .B(_12534_),
    .Y(_12535_));
 NOR2x1_ASAP7_75t_SL _20773_ (.A(_12527_),
    .B(_12535_),
    .Y(_12536_));
 NAND2x1_ASAP7_75t_SL _20774_ (.A(_12196_),
    .B(_12455_),
    .Y(_12537_));
 NAND2x1_ASAP7_75t_SL _20775_ (.A(_12463_),
    .B(_12140_),
    .Y(_12538_));
 NAND2x1_ASAP7_75t_SL _20776_ (.A(_12538_),
    .B(_12243_),
    .Y(_12539_));
 AOI21x1_ASAP7_75t_SL _20777_ (.A1(_12539_),
    .A2(_12341_),
    .B(_12283_),
    .Y(_12540_));
 OAI21x1_ASAP7_75t_SL _20778_ (.A1(_12537_),
    .A2(_12540_),
    .B(_12247_),
    .Y(_12541_));
 INVx1_ASAP7_75t_SL _20779_ (.A(_12326_),
    .Y(_12542_));
 NOR2x1_ASAP7_75t_SL _20780_ (.A(_12278_),
    .B(_12528_),
    .Y(_12543_));
 OA21x2_ASAP7_75t_SL _20781_ (.A1(_12394_),
    .A2(_12114_),
    .B(_12283_),
    .Y(_12544_));
 OAI21x1_ASAP7_75t_SL _20782_ (.A1(_12542_),
    .A2(_12543_),
    .B(_12544_),
    .Y(_12545_));
 NAND3x1_ASAP7_75t_SL _20783_ (.A(_12259_),
    .B(_12393_),
    .C(_12167_),
    .Y(_12546_));
 AOI21x1_ASAP7_75t_SL _20784_ (.A1(_12545_),
    .A2(_12546_),
    .B(_12196_),
    .Y(_12547_));
 NOR2x1_ASAP7_75t_SL _20785_ (.A(_12541_),
    .B(_12547_),
    .Y(_12548_));
 OAI21x1_ASAP7_75t_SL _20786_ (.A1(_12536_),
    .A2(_12548_),
    .B(_12274_),
    .Y(_12549_));
 NAND2x1_ASAP7_75t_SL _20787_ (.A(_12521_),
    .B(_12549_),
    .Y(_00051_));
 OAI21x1_ASAP7_75t_SL _20788_ (.A1(_12173_),
    .A2(_12257_),
    .B(_12283_),
    .Y(_12550_));
 OAI21x1_ASAP7_75t_SL _20789_ (.A1(_12173_),
    .A2(_12309_),
    .B(_12353_),
    .Y(_12551_));
 NOR2x1_ASAP7_75t_SL _20790_ (.A(_12283_),
    .B(_12417_),
    .Y(_12552_));
 NAND2x1_ASAP7_75t_SL _20791_ (.A(_12326_),
    .B(_12290_),
    .Y(_12553_));
 AOI21x1_ASAP7_75t_SL _20792_ (.A1(_12552_),
    .A2(_12553_),
    .B(_12197_),
    .Y(_12554_));
 OAI21x1_ASAP7_75t_SL _20793_ (.A1(_12550_),
    .A2(_12551_),
    .B(_12554_),
    .Y(_12555_));
 AOI21x1_ASAP7_75t_SL _20794_ (.A1(_12172_),
    .A2(_12389_),
    .B(_12283_),
    .Y(_12556_));
 NAND2x1_ASAP7_75t_SL _20795_ (.A(_12556_),
    .B(_12209_),
    .Y(_12557_));
 AOI21x1_ASAP7_75t_SL _20796_ (.A1(_12154_),
    .A2(_12365_),
    .B(_12167_),
    .Y(_12558_));
 AO21x1_ASAP7_75t_SL _20797_ (.A1(_12207_),
    .A2(_12132_),
    .B(_12154_),
    .Y(_12559_));
 AOI21x1_ASAP7_75t_SL _20798_ (.A1(_12558_),
    .A2(_12559_),
    .B(_12196_),
    .Y(_12560_));
 NAND2x1_ASAP7_75t_SL _20799_ (.A(_12557_),
    .B(_12560_),
    .Y(_12561_));
 AOI21x1_ASAP7_75t_SL _20800_ (.A1(_12555_),
    .A2(_12561_),
    .B(_12228_),
    .Y(_12562_));
 OR2x2_ASAP7_75t_SL _20801_ (.A(_12173_),
    .B(_01112_),
    .Y(_12563_));
 NAND2x1_ASAP7_75t_SL _20802_ (.A(_12173_),
    .B(_12261_),
    .Y(_12564_));
 AND3x1_ASAP7_75t_SL _20803_ (.A(_12563_),
    .B(_12167_),
    .C(_12564_),
    .Y(_12565_));
 NAND2x1_ASAP7_75t_SL _20804_ (.A(_12380_),
    .B(_12243_),
    .Y(_12566_));
 NAND2x1_ASAP7_75t_SL _20805_ (.A(_12154_),
    .B(_12250_),
    .Y(_12567_));
 AOI21x1_ASAP7_75t_SL _20806_ (.A1(_12566_),
    .A2(_12567_),
    .B(_12167_),
    .Y(_12568_));
 OAI21x1_ASAP7_75t_SL _20807_ (.A1(_12565_),
    .A2(_12568_),
    .B(_12197_),
    .Y(_12569_));
 NAND2x1_ASAP7_75t_SL _20808_ (.A(_12141_),
    .B(_12243_),
    .Y(_12570_));
 NOR2x2_ASAP7_75t_SL _20809_ (.A(_12132_),
    .B(_12096_),
    .Y(_12571_));
 OAI21x1_ASAP7_75t_SL _20810_ (.A1(_12207_),
    .A2(_12571_),
    .B(_12154_),
    .Y(_12572_));
 AOI21x1_ASAP7_75t_SL _20811_ (.A1(_12570_),
    .A2(_12572_),
    .B(_12167_),
    .Y(_12573_));
 AOI21x1_ASAP7_75t_SL _20812_ (.A1(_12288_),
    .A2(_12188_),
    .B(_12283_),
    .Y(_12574_));
 OAI21x1_ASAP7_75t_SL _20813_ (.A1(_12573_),
    .A2(_12574_),
    .B(_12196_),
    .Y(_12575_));
 AOI21x1_ASAP7_75t_SL _20814_ (.A1(_12569_),
    .A2(_12575_),
    .B(_12247_),
    .Y(_12576_));
 OAI21x1_ASAP7_75t_SL _20815_ (.A1(_12562_),
    .A2(_12576_),
    .B(_12274_),
    .Y(_12577_));
 AO21x1_ASAP7_75t_SL _20816_ (.A1(_12309_),
    .A2(_12141_),
    .B(_12154_),
    .Y(_12578_));
 NAND2x1_ASAP7_75t_SL _20817_ (.A(_12347_),
    .B(_12578_),
    .Y(_12579_));
 NOR2x1_ASAP7_75t_SL _20818_ (.A(_12361_),
    .B(_12243_),
    .Y(_12580_));
 AOI21x1_ASAP7_75t_SL _20819_ (.A1(_12283_),
    .A2(_12580_),
    .B(_12196_),
    .Y(_12581_));
 OAI21x1_ASAP7_75t_SL _20820_ (.A1(_12283_),
    .A2(_12579_),
    .B(_12581_),
    .Y(_12582_));
 NAND2x1_ASAP7_75t_SL _20821_ (.A(_12277_),
    .B(_12290_),
    .Y(_12583_));
 NAND2x1_ASAP7_75t_SL _20822_ (.A(_12442_),
    .B(_12474_),
    .Y(_12584_));
 AOI21x1_ASAP7_75t_SL _20823_ (.A1(_12583_),
    .A2(_12584_),
    .B(_12283_),
    .Y(_12585_));
 OAI21x1_ASAP7_75t_SL _20824_ (.A1(_12354_),
    .A2(_12317_),
    .B(_12173_),
    .Y(_12586_));
 OAI21x1_ASAP7_75t_SL _20825_ (.A1(_12232_),
    .A2(_12430_),
    .B(_12154_),
    .Y(_12587_));
 AOI21x1_ASAP7_75t_SL _20826_ (.A1(_12586_),
    .A2(_12587_),
    .B(_12167_),
    .Y(_12588_));
 OAI21x1_ASAP7_75t_SL _20827_ (.A1(_12585_),
    .A2(_12588_),
    .B(_12196_),
    .Y(_12589_));
 AOI21x1_ASAP7_75t_SL _20828_ (.A1(_12582_),
    .A2(_12589_),
    .B(_12228_),
    .Y(_12590_));
 AO21x1_ASAP7_75t_SL _20829_ (.A1(_12131_),
    .A2(_12129_),
    .B(_12171_),
    .Y(_12591_));
 AND2x2_ASAP7_75t_SL _20830_ (.A(_12366_),
    .B(_12591_),
    .Y(_12592_));
 AO21x1_ASAP7_75t_SL _20831_ (.A1(_12233_),
    .A2(_12243_),
    .B(_12283_),
    .Y(_12593_));
 AND2x2_ASAP7_75t_SL _20832_ (.A(_12564_),
    .B(_12217_),
    .Y(_12594_));
 OA21x2_ASAP7_75t_SL _20833_ (.A1(_12200_),
    .A2(_12173_),
    .B(_12283_),
    .Y(_12595_));
 AOI21x1_ASAP7_75t_SL _20834_ (.A1(_12594_),
    .A2(_12595_),
    .B(_12196_),
    .Y(_12596_));
 OAI21x1_ASAP7_75t_SL _20835_ (.A1(_12592_),
    .A2(_12593_),
    .B(_12596_),
    .Y(_12597_));
 NAND2x1_ASAP7_75t_SL _20836_ (.A(_12167_),
    .B(_12251_),
    .Y(_12598_));
 AOI21x1_ASAP7_75t_SL _20837_ (.A1(_12257_),
    .A2(_12277_),
    .B(_12154_),
    .Y(_12599_));
 AOI21x1_ASAP7_75t_SL _20838_ (.A1(_12326_),
    .A2(_12389_),
    .B(_12167_),
    .Y(_12600_));
 NAND2x1_ASAP7_75t_SL _20839_ (.A(_12481_),
    .B(_12233_),
    .Y(_12601_));
 AOI21x1_ASAP7_75t_SL _20840_ (.A1(_12600_),
    .A2(_12601_),
    .B(_12197_),
    .Y(_12602_));
 OAI21x1_ASAP7_75t_SL _20841_ (.A1(_12598_),
    .A2(_12599_),
    .B(_12602_),
    .Y(_12603_));
 AOI21x1_ASAP7_75t_SL _20842_ (.A1(_12597_),
    .A2(_12603_),
    .B(_12247_),
    .Y(_12604_));
 OAI21x1_ASAP7_75t_SL _20843_ (.A1(_12590_),
    .A2(_12604_),
    .B(_12520_),
    .Y(_12605_));
 NAND2x1_ASAP7_75t_SL _20844_ (.A(_12577_),
    .B(_12605_),
    .Y(_00052_));
 AO21x1_ASAP7_75t_SL _20845_ (.A1(_01110_),
    .A2(_12173_),
    .B(_12283_),
    .Y(_12606_));
 AO21x1_ASAP7_75t_SL _20846_ (.A1(_12208_),
    .A2(_12154_),
    .B(_12606_),
    .Y(_12607_));
 AND2x2_ASAP7_75t_SL _20847_ (.A(_12607_),
    .B(_12196_),
    .Y(_12608_));
 AO221x1_ASAP7_75t_SL _20848_ (.A1(_12326_),
    .A2(_12304_),
    .B1(_12212_),
    .B2(_12236_),
    .C(_12167_),
    .Y(_12609_));
 AND2x2_ASAP7_75t_SL _20849_ (.A(_12608_),
    .B(_12609_),
    .Y(_12610_));
 OA21x2_ASAP7_75t_SL _20850_ (.A1(_12404_),
    .A2(_12381_),
    .B(_12197_),
    .Y(_12611_));
 NOR2x1_ASAP7_75t_R _20851_ (.A(_12173_),
    .B(_12096_),
    .Y(_12612_));
 INVx1_ASAP7_75t_SL _20852_ (.A(_12612_),
    .Y(_12613_));
 NAND2x1_ASAP7_75t_SL _20853_ (.A(_12613_),
    .B(_12331_),
    .Y(_12614_));
 AO21x1_ASAP7_75t_SL _20854_ (.A1(_12538_),
    .A2(_12173_),
    .B(_12283_),
    .Y(_12615_));
 AO21x1_ASAP7_75t_SL _20855_ (.A1(_12614_),
    .A2(_12208_),
    .B(_12615_),
    .Y(_12616_));
 AO21x1_ASAP7_75t_SL _20856_ (.A1(_12611_),
    .A2(_12616_),
    .B(_12247_),
    .Y(_12617_));
 OA21x2_ASAP7_75t_SL _20857_ (.A1(_12136_),
    .A2(_12154_),
    .B(_12167_),
    .Y(_12618_));
 AOI21x1_ASAP7_75t_SL _20858_ (.A1(_12618_),
    .A2(_12291_),
    .B(_12196_),
    .Y(_12619_));
 AOI21x1_ASAP7_75t_SL _20859_ (.A1(_12380_),
    .A2(_12449_),
    .B(_12167_),
    .Y(_12620_));
 NAND2x1_ASAP7_75t_SL _20860_ (.A(_12212_),
    .B(_12329_),
    .Y(_12621_));
 NAND2x1_ASAP7_75t_SL _20861_ (.A(_12620_),
    .B(_12621_),
    .Y(_12622_));
 AOI21x1_ASAP7_75t_SL _20862_ (.A1(_12619_),
    .A2(_12622_),
    .B(_12228_),
    .Y(_12623_));
 NAND2x1_ASAP7_75t_SL _20863_ (.A(_12154_),
    .B(_12427_),
    .Y(_12624_));
 INVx1_ASAP7_75t_SL _20864_ (.A(_12624_),
    .Y(_12625_));
 OA21x2_ASAP7_75t_SL _20865_ (.A1(_12144_),
    .A2(_12154_),
    .B(_12283_),
    .Y(_12626_));
 NOR2x1_ASAP7_75t_R _20866_ (.A(_12114_),
    .B(_12173_),
    .Y(_12627_));
 OAI21x1_ASAP7_75t_SL _20867_ (.A1(_12627_),
    .A2(_12175_),
    .B(_12326_),
    .Y(_12628_));
 AOI21x1_ASAP7_75t_SL _20868_ (.A1(_12626_),
    .A2(_12628_),
    .B(_12197_),
    .Y(_12629_));
 OAI21x1_ASAP7_75t_SL _20869_ (.A1(_12210_),
    .A2(_12625_),
    .B(_12629_),
    .Y(_12630_));
 AOI21x1_ASAP7_75t_SL _20870_ (.A1(_12623_),
    .A2(_12630_),
    .B(_12520_),
    .Y(_12631_));
 OAI21x1_ASAP7_75t_SL _20871_ (.A1(_12610_),
    .A2(_12617_),
    .B(_12631_),
    .Y(_12632_));
 AND2x2_ASAP7_75t_SL _20872_ (.A(_12212_),
    .B(_12186_),
    .Y(_12633_));
 AO21x1_ASAP7_75t_SL _20873_ (.A1(_12439_),
    .A2(_12154_),
    .B(_12283_),
    .Y(_12634_));
 OAI21x1_ASAP7_75t_SL _20874_ (.A1(_12633_),
    .A2(_12634_),
    .B(_12196_),
    .Y(_12635_));
 AO21x1_ASAP7_75t_SL _20875_ (.A1(_12380_),
    .A2(_12254_),
    .B(_12173_),
    .Y(_12636_));
 AOI21x1_ASAP7_75t_SL _20876_ (.A1(_12564_),
    .A2(_12636_),
    .B(_12167_),
    .Y(_12637_));
 OAI21x1_ASAP7_75t_SL _20877_ (.A1(_12635_),
    .A2(_12637_),
    .B(_12228_),
    .Y(_12638_));
 OR3x1_ASAP7_75t_SL _20878_ (.A(_12340_),
    .B(_12154_),
    .C(_12339_),
    .Y(_12639_));
 OA21x2_ASAP7_75t_SL _20879_ (.A1(_12331_),
    .A2(_12207_),
    .B(_12283_),
    .Y(_12640_));
 NOR2x1_ASAP7_75t_SL _20880_ (.A(_12283_),
    .B(_12418_),
    .Y(_12641_));
 AO21x1_ASAP7_75t_SL _20881_ (.A1(_12572_),
    .A2(_12641_),
    .B(_12196_),
    .Y(_12642_));
 AOI21x1_ASAP7_75t_SL _20882_ (.A1(_12639_),
    .A2(_12640_),
    .B(_12642_),
    .Y(_12643_));
 NOR2x1_ASAP7_75t_SL _20883_ (.A(_12638_),
    .B(_12643_),
    .Y(_12644_));
 AO21x1_ASAP7_75t_SL _20884_ (.A1(_12419_),
    .A2(_12417_),
    .B(_12389_),
    .Y(_12645_));
 AOI21x1_ASAP7_75t_SL _20885_ (.A1(_12136_),
    .A2(_12417_),
    .B(_12283_),
    .Y(_12646_));
 AOI21x1_ASAP7_75t_SL _20886_ (.A1(_12646_),
    .A2(_12543_),
    .B(_12197_),
    .Y(_12647_));
 OAI21x1_ASAP7_75t_SL _20887_ (.A1(_12167_),
    .A2(_12645_),
    .B(_12647_),
    .Y(_12648_));
 NAND2x1_ASAP7_75t_SL _20888_ (.A(_12449_),
    .B(_12233_),
    .Y(_12649_));
 NAND2x1_ASAP7_75t_SL _20889_ (.A(_01108_),
    .B(_12184_),
    .Y(_12650_));
 AOI21x1_ASAP7_75t_SL _20890_ (.A1(_12173_),
    .A2(_12650_),
    .B(_12167_),
    .Y(_12651_));
 AOI21x1_ASAP7_75t_SL _20891_ (.A1(_12649_),
    .A2(_12651_),
    .B(_12196_),
    .Y(_12652_));
 NAND2x1_ASAP7_75t_SL _20892_ (.A(_12326_),
    .B(_12182_),
    .Y(_12653_));
 NAND3x1_ASAP7_75t_SL _20893_ (.A(_12311_),
    .B(_12167_),
    .C(_12653_),
    .Y(_12654_));
 NAND2x1_ASAP7_75t_SL _20894_ (.A(_12652_),
    .B(_12654_),
    .Y(_12655_));
 AOI21x1_ASAP7_75t_SL _20895_ (.A1(_12648_),
    .A2(_12655_),
    .B(_12228_),
    .Y(_12656_));
 OAI21x1_ASAP7_75t_SL _20896_ (.A1(_12644_),
    .A2(_12656_),
    .B(_12520_),
    .Y(_12657_));
 NAND2x1_ASAP7_75t_SL _20897_ (.A(_12632_),
    .B(_12657_),
    .Y(_00053_));
 AND2x2_ASAP7_75t_SL _20898_ (.A(_12525_),
    .B(_12283_),
    .Y(_12658_));
 NAND2x1_ASAP7_75t_SL _20899_ (.A(_12467_),
    .B(_12324_),
    .Y(_12659_));
 AOI21x1_ASAP7_75t_SL _20900_ (.A1(_12658_),
    .A2(_12659_),
    .B(_12196_),
    .Y(_12660_));
 OAI21x1_ASAP7_75t_SL _20901_ (.A1(_12317_),
    .A2(_12318_),
    .B(_12173_),
    .Y(_12661_));
 NAND2x1_ASAP7_75t_SL _20902_ (.A(_12365_),
    .B(_12304_),
    .Y(_12662_));
 AO21x1_ASAP7_75t_SL _20903_ (.A1(_12661_),
    .A2(_12662_),
    .B(_12283_),
    .Y(_12663_));
 NAND2x1_ASAP7_75t_SL _20904_ (.A(_12660_),
    .B(_12663_),
    .Y(_12664_));
 AND3x1_ASAP7_75t_SL _20905_ (.A(_12538_),
    .B(_12154_),
    .C(_12172_),
    .Y(_12665_));
 NAND2x1_ASAP7_75t_SL _20906_ (.A(_12646_),
    .B(_12288_),
    .Y(_12666_));
 AOI21x1_ASAP7_75t_SL _20907_ (.A1(_12154_),
    .A2(_12339_),
    .B(_12167_),
    .Y(_12667_));
 OAI21x1_ASAP7_75t_SL _20908_ (.A1(_12232_),
    .A2(_12402_),
    .B(_12667_),
    .Y(_12668_));
 OAI21x1_ASAP7_75t_SL _20909_ (.A1(_12665_),
    .A2(_12666_),
    .B(_12668_),
    .Y(_12669_));
 AOI21x1_ASAP7_75t_SL _20910_ (.A1(_12196_),
    .A2(_12669_),
    .B(_12247_),
    .Y(_12670_));
 NAND2x1_ASAP7_75t_R _20911_ (.A(_12217_),
    .B(_12200_),
    .Y(_12671_));
 NOR2x1_ASAP7_75t_SL _20912_ (.A(_12428_),
    .B(_12671_),
    .Y(_12672_));
 NAND2x1_ASAP7_75t_SL _20913_ (.A(_12262_),
    .B(_12624_),
    .Y(_12673_));
 OAI21x1_ASAP7_75t_SL _20914_ (.A1(_12672_),
    .A2(_12673_),
    .B(_12196_),
    .Y(_12674_));
 INVx1_ASAP7_75t_SL _20915_ (.A(_12207_),
    .Y(_12675_));
 NAND2x1_ASAP7_75t_SL _20916_ (.A(_12417_),
    .B(_12675_),
    .Y(_12676_));
 OAI21x1_ASAP7_75t_R _20917_ (.A1(_12130_),
    .A2(_12169_),
    .B(_12216_),
    .Y(_12677_));
 AOI21x1_ASAP7_75t_SL _20918_ (.A1(_12496_),
    .A2(_12677_),
    .B(_12173_),
    .Y(_12678_));
 NOR2x1_ASAP7_75t_SL _20919_ (.A(_12239_),
    .B(_12678_),
    .Y(_12679_));
 AOI21x1_ASAP7_75t_SL _20920_ (.A1(_12676_),
    .A2(_12679_),
    .B(_12283_),
    .Y(_12680_));
 NOR2x1_ASAP7_75t_SL _20921_ (.A(_12674_),
    .B(_12680_),
    .Y(_12681_));
 AOI21x1_ASAP7_75t_SL _20922_ (.A1(_12217_),
    .A2(_12254_),
    .B(_12154_),
    .Y(_12682_));
 NOR2x1_ASAP7_75t_SL _20923_ (.A(_12550_),
    .B(_12682_),
    .Y(_12683_));
 AND2x2_ASAP7_75t_R _20924_ (.A(_01121_),
    .B(_01115_),
    .Y(_12684_));
 OAI21x1_ASAP7_75t_SL _20925_ (.A1(_12684_),
    .A2(_12173_),
    .B(_12167_),
    .Y(_12685_));
 AOI21x1_ASAP7_75t_SL _20926_ (.A1(_12419_),
    .A2(_12481_),
    .B(_12685_),
    .Y(_12686_));
 OAI21x1_ASAP7_75t_SL _20927_ (.A1(_12683_),
    .A2(_12686_),
    .B(_12197_),
    .Y(_12687_));
 NAND2x1_ASAP7_75t_SL _20928_ (.A(_12247_),
    .B(_12687_),
    .Y(_12688_));
 NOR2x1_ASAP7_75t_SL _20929_ (.A(_12681_),
    .B(_12688_),
    .Y(_12689_));
 AOI21x1_ASAP7_75t_SL _20930_ (.A1(_12664_),
    .A2(_12670_),
    .B(_12689_),
    .Y(_12690_));
 NOR2x1_ASAP7_75t_SL _20931_ (.A(_12366_),
    .B(_12474_),
    .Y(_12691_));
 OAI21x1_ASAP7_75t_SL _20932_ (.A1(_12360_),
    .A2(_12691_),
    .B(_12283_),
    .Y(_12692_));
 OAI21x1_ASAP7_75t_SL _20933_ (.A1(_12096_),
    .A2(_12114_),
    .B(_12167_),
    .Y(_12693_));
 NOR2x1_ASAP7_75t_SL _20934_ (.A(_12360_),
    .B(_12693_),
    .Y(_12694_));
 AOI21x1_ASAP7_75t_SL _20935_ (.A1(_12613_),
    .A2(_12694_),
    .B(_12196_),
    .Y(_12695_));
 NAND2x1_ASAP7_75t_SL _20936_ (.A(_12692_),
    .B(_12695_),
    .Y(_12696_));
 AOI21x1_ASAP7_75t_SL _20937_ (.A1(_12173_),
    .A2(_12277_),
    .B(_12167_),
    .Y(_12697_));
 OAI21x1_ASAP7_75t_SL _20938_ (.A1(_12322_),
    .A2(_12324_),
    .B(_12697_),
    .Y(_12698_));
 NAND2x1_ASAP7_75t_SL _20939_ (.A(_12452_),
    .B(_12429_),
    .Y(_12699_));
 AOI21x1_ASAP7_75t_SL _20940_ (.A1(_12646_),
    .A2(_12699_),
    .B(_12197_),
    .Y(_12700_));
 NAND2x1_ASAP7_75t_SL _20941_ (.A(_12698_),
    .B(_12700_),
    .Y(_12701_));
 AOI21x1_ASAP7_75t_SL _20942_ (.A1(_12696_),
    .A2(_12701_),
    .B(_12228_),
    .Y(_12702_));
 AOI21x1_ASAP7_75t_SL _20943_ (.A1(_12154_),
    .A2(_12360_),
    .B(_12167_),
    .Y(_12703_));
 NAND2x1_ASAP7_75t_SL _20944_ (.A(_12298_),
    .B(_12381_),
    .Y(_12704_));
 NAND2x1_ASAP7_75t_SL _20945_ (.A(_12703_),
    .B(_12704_),
    .Y(_12705_));
 AOI21x1_ASAP7_75t_SL _20946_ (.A1(_01116_),
    .A2(_12173_),
    .B(_12283_),
    .Y(_12706_));
 NAND2x1_ASAP7_75t_SL _20947_ (.A(_12380_),
    .B(_12449_),
    .Y(_12707_));
 NAND2x1_ASAP7_75t_SL _20948_ (.A(_12706_),
    .B(_12707_),
    .Y(_12708_));
 NAND3x1_ASAP7_75t_SL _20949_ (.A(_12705_),
    .B(_12708_),
    .C(_12197_),
    .Y(_12709_));
 AOI21x1_ASAP7_75t_SL _20950_ (.A1(_12237_),
    .A2(_12566_),
    .B(_12167_),
    .Y(_12710_));
 OAI21x1_ASAP7_75t_SL _20951_ (.A1(_12710_),
    .A2(_12424_),
    .B(_12196_),
    .Y(_12711_));
 AOI21x1_ASAP7_75t_SL _20952_ (.A1(_12709_),
    .A2(_12711_),
    .B(_12247_),
    .Y(_12712_));
 OAI21x1_ASAP7_75t_SL _20953_ (.A1(_12702_),
    .A2(_12712_),
    .B(_12274_),
    .Y(_12713_));
 OAI21x1_ASAP7_75t_SL _20954_ (.A1(_12274_),
    .A2(_12690_),
    .B(_12713_),
    .Y(_00054_));
 OA21x2_ASAP7_75t_SL _20955_ (.A1(_01108_),
    .A2(_12173_),
    .B(_12283_),
    .Y(_12714_));
 NAND2x1_ASAP7_75t_SL _20956_ (.A(_12481_),
    .B(_12419_),
    .Y(_12715_));
 AOI21x1_ASAP7_75t_SL _20957_ (.A1(_12714_),
    .A2(_12715_),
    .B(_12197_),
    .Y(_12716_));
 OA21x2_ASAP7_75t_SL _20958_ (.A1(_12309_),
    .A2(_12154_),
    .B(_12257_),
    .Y(_12717_));
 NAND2x1_ASAP7_75t_SL _20959_ (.A(_12255_),
    .B(_12717_),
    .Y(_12718_));
 AOI21x1_ASAP7_75t_SL _20960_ (.A1(_12716_),
    .A2(_12718_),
    .B(_12228_),
    .Y(_12719_));
 AO21x1_ASAP7_75t_SL _20961_ (.A1(_12323_),
    .A2(_12096_),
    .B(_12173_),
    .Y(_12720_));
 AOI21x1_ASAP7_75t_SL _20962_ (.A1(_12539_),
    .A2(_12720_),
    .B(_12167_),
    .Y(_12721_));
 AND2x2_ASAP7_75t_SL _20963_ (.A(_12212_),
    .B(_12144_),
    .Y(_12722_));
 NAND2x1_ASAP7_75t_SL _20964_ (.A(_12257_),
    .B(_12309_),
    .Y(_12723_));
 OAI21x1_ASAP7_75t_SL _20965_ (.A1(_12331_),
    .A2(_12723_),
    .B(_12167_),
    .Y(_12724_));
 NOR2x1_ASAP7_75t_SL _20966_ (.A(_12722_),
    .B(_12724_),
    .Y(_12725_));
 OAI21x1_ASAP7_75t_SL _20967_ (.A1(_12721_),
    .A2(_12725_),
    .B(_12197_),
    .Y(_12726_));
 AOI21x1_ASAP7_75t_SL _20968_ (.A1(_12719_),
    .A2(_12726_),
    .B(_12274_),
    .Y(_12727_));
 AOI21x1_ASAP7_75t_SL _20969_ (.A1(_12217_),
    .A2(_12591_),
    .B(_12173_),
    .Y(_12728_));
 NOR2x1_ASAP7_75t_SL _20970_ (.A(_01121_),
    .B(_12154_),
    .Y(_12729_));
 OA21x2_ASAP7_75t_SL _20971_ (.A1(_12728_),
    .A2(_12729_),
    .B(_12167_),
    .Y(_12730_));
 NAND2x1_ASAP7_75t_SL _20972_ (.A(_12298_),
    .B(_12302_),
    .Y(_12731_));
 AO21x1_ASAP7_75t_SL _20973_ (.A1(_12442_),
    .A2(_12256_),
    .B(_12173_),
    .Y(_12732_));
 AOI21x1_ASAP7_75t_SL _20974_ (.A1(_12731_),
    .A2(_12732_),
    .B(_12167_),
    .Y(_12733_));
 OAI21x1_ASAP7_75t_SL _20975_ (.A1(_12730_),
    .A2(_12733_),
    .B(_12196_),
    .Y(_12734_));
 AO21x1_ASAP7_75t_SL _20976_ (.A1(_12427_),
    .A2(_12154_),
    .B(_12612_),
    .Y(_12735_));
 NAND2x1_ASAP7_75t_SL _20977_ (.A(_01112_),
    .B(_12173_),
    .Y(_12736_));
 AOI21x1_ASAP7_75t_SL _20978_ (.A1(_12736_),
    .A2(_12255_),
    .B(_12196_),
    .Y(_12737_));
 OAI21x1_ASAP7_75t_SL _20979_ (.A1(_12349_),
    .A2(_12735_),
    .B(_12737_),
    .Y(_12738_));
 NAND3x1_ASAP7_75t_SL _20980_ (.A(_12734_),
    .B(_12228_),
    .C(_12738_),
    .Y(_12739_));
 NAND2x1_ASAP7_75t_SL _20981_ (.A(_12727_),
    .B(_12739_),
    .Y(_12740_));
 AOI21x1_ASAP7_75t_SL _20982_ (.A1(_12531_),
    .A2(_12400_),
    .B(_12167_),
    .Y(_12741_));
 INVx1_ASAP7_75t_SL _20983_ (.A(_12678_),
    .Y(_12742_));
 AOI21x1_ASAP7_75t_SL _20984_ (.A1(_12742_),
    .A2(_12482_),
    .B(_12283_),
    .Y(_12743_));
 OAI21x1_ASAP7_75t_SL _20985_ (.A1(_12741_),
    .A2(_12743_),
    .B(_12196_),
    .Y(_12744_));
 OA21x2_ASAP7_75t_SL _20986_ (.A1(_12723_),
    .A2(_12203_),
    .B(_12173_),
    .Y(_12745_));
 AO21x1_ASAP7_75t_SL _20987_ (.A1(_12372_),
    .A2(_12233_),
    .B(_12167_),
    .Y(_12746_));
 AOI21x1_ASAP7_75t_SL _20988_ (.A1(_12380_),
    .A2(_12243_),
    .B(_12366_),
    .Y(_12747_));
 AOI21x1_ASAP7_75t_SL _20989_ (.A1(_12167_),
    .A2(_12747_),
    .B(_12196_),
    .Y(_12748_));
 OAI21x1_ASAP7_75t_SL _20990_ (.A1(_12745_),
    .A2(_12746_),
    .B(_12748_),
    .Y(_12749_));
 AOI21x1_ASAP7_75t_SL _20991_ (.A1(_12744_),
    .A2(_12749_),
    .B(_12228_),
    .Y(_12750_));
 OA21x2_ASAP7_75t_SL _20992_ (.A1(_12207_),
    .A2(_12506_),
    .B(_12167_),
    .Y(_12751_));
 NAND2x1_ASAP7_75t_SL _20993_ (.A(_12525_),
    .B(_12751_),
    .Y(_12752_));
 OAI21x1_ASAP7_75t_SL _20994_ (.A1(_12136_),
    .A2(_12277_),
    .B(_12304_),
    .Y(_12753_));
 NOR3x1_ASAP7_75t_SL _20995_ (.A(_12287_),
    .B(_12167_),
    .C(_12417_),
    .Y(_12754_));
 AOI21x1_ASAP7_75t_SL _20996_ (.A1(_12753_),
    .A2(_12754_),
    .B(_12197_),
    .Y(_12755_));
 NAND2x1_ASAP7_75t_SL _20997_ (.A(_12752_),
    .B(_12755_),
    .Y(_12756_));
 AO21x1_ASAP7_75t_SL _20998_ (.A1(_12207_),
    .A2(_12132_),
    .B(_12173_),
    .Y(_12757_));
 OAI21x1_ASAP7_75t_SL _20999_ (.A1(_12571_),
    .A2(_12757_),
    .B(_12475_),
    .Y(_12758_));
 INVx1_ASAP7_75t_SL _21000_ (.A(_12627_),
    .Y(_12759_));
 OAI21x1_ASAP7_75t_SL _21001_ (.A1(_12322_),
    .A2(_12402_),
    .B(_12759_),
    .Y(_12760_));
 AOI21x1_ASAP7_75t_SL _21002_ (.A1(_12283_),
    .A2(_12760_),
    .B(_12196_),
    .Y(_12761_));
 NAND2x1_ASAP7_75t_SL _21003_ (.A(_12758_),
    .B(_12761_),
    .Y(_12762_));
 AOI21x1_ASAP7_75t_SL _21004_ (.A1(_12756_),
    .A2(_12762_),
    .B(_12247_),
    .Y(_12763_));
 OAI21x1_ASAP7_75t_SL _21005_ (.A1(_12750_),
    .A2(_12763_),
    .B(_12274_),
    .Y(_12764_));
 NAND2x1_ASAP7_75t_SL _21006_ (.A(_12740_),
    .B(_12764_),
    .Y(_00055_));
 NOR2x1_ASAP7_75t_R _21007_ (.A(_00574_),
    .B(_00453_),
    .Y(_12765_));
 XOR2x2_ASAP7_75t_SL _21008_ (.A(_00638_),
    .B(_00631_),
    .Y(_12766_));
 XOR2x2_ASAP7_75t_L _21009_ (.A(_12766_),
    .B(_00696_),
    .Y(_12767_));
 XOR2x2_ASAP7_75t_SL _21010_ (.A(_00599_),
    .B(_00606_),
    .Y(_12768_));
 XOR2x2_ASAP7_75t_SL _21011_ (.A(_00632_),
    .B(_00664_),
    .Y(_12769_));
 XOR2x2_ASAP7_75t_L _21012_ (.A(_12768_),
    .B(_12769_),
    .Y(_12770_));
 NAND2x1_ASAP7_75t_SL _21013_ (.A(_12767_),
    .B(_12770_),
    .Y(_12771_));
 INVx1_ASAP7_75t_R _21014_ (.A(_00696_),
    .Y(_12772_));
 XOR2x2_ASAP7_75t_L _21015_ (.A(_12766_),
    .B(_12772_),
    .Y(_12773_));
 XNOR2x2_ASAP7_75t_SL _21016_ (.A(_00599_),
    .B(_00606_),
    .Y(_12774_));
 XOR2x2_ASAP7_75t_L _21017_ (.A(_12774_),
    .B(_12769_),
    .Y(_12775_));
 NAND2x1_ASAP7_75t_SL _21018_ (.A(_12773_),
    .B(_12775_),
    .Y(_12776_));
 AOI21x1_ASAP7_75t_R _21019_ (.A1(_12771_),
    .A2(_12776_),
    .B(_10675_),
    .Y(_12777_));
 OAI21x1_ASAP7_75t_SL _21020_ (.A1(_12777_),
    .A2(_12765_),
    .B(_00951_),
    .Y(_12778_));
 AND2x2_ASAP7_75t_R _21021_ (.A(_10675_),
    .B(_00453_),
    .Y(_12779_));
 NAND2x1_ASAP7_75t_R _21022_ (.A(_12773_),
    .B(_12770_),
    .Y(_12780_));
 NAND2x1_ASAP7_75t_R _21023_ (.A(_12767_),
    .B(_12775_),
    .Y(_12781_));
 AOI21x1_ASAP7_75t_R _21024_ (.A1(_12780_),
    .A2(_12781_),
    .B(_10675_),
    .Y(_12782_));
 INVx1_ASAP7_75t_R _21025_ (.A(_00951_),
    .Y(_12783_));
 OAI21x1_ASAP7_75t_SL _21026_ (.A1(_12782_),
    .A2(_12779_),
    .B(_12783_),
    .Y(_12784_));
 NAND2x2_ASAP7_75t_SL _21027_ (.A(_12784_),
    .B(_12778_),
    .Y(_12785_));
 INVx1_ASAP7_75t_R _21029_ (.A(_00695_),
    .Y(_12786_));
 XOR2x2_ASAP7_75t_SL _21030_ (.A(_00638_),
    .B(_00606_),
    .Y(_12787_));
 NAND2x1_ASAP7_75t_L _21031_ (.A(_12786_),
    .B(_12787_),
    .Y(_12788_));
 XNOR2x2_ASAP7_75t_SL _21032_ (.A(_00606_),
    .B(_00638_),
    .Y(_12789_));
 NAND2x1_ASAP7_75t_L _21033_ (.A(_00695_),
    .B(_12789_),
    .Y(_12790_));
 XOR2x2_ASAP7_75t_SL _21034_ (.A(_00631_),
    .B(_00663_),
    .Y(_12791_));
 INVx1_ASAP7_75t_R _21035_ (.A(_12791_),
    .Y(_12792_));
 AOI21x1_ASAP7_75t_SL _21036_ (.A1(_12790_),
    .A2(_12788_),
    .B(_12792_),
    .Y(_12793_));
 NAND2x1_ASAP7_75t_L _21037_ (.A(_00695_),
    .B(_12787_),
    .Y(_12794_));
 NAND2x1p5_ASAP7_75t_L _21038_ (.A(_12786_),
    .B(_12789_),
    .Y(_12795_));
 AOI21x1_ASAP7_75t_SL _21039_ (.A1(_12795_),
    .A2(_12794_),
    .B(_12791_),
    .Y(_12796_));
 OAI21x1_ASAP7_75t_SL _21040_ (.A1(_12796_),
    .A2(_12793_),
    .B(_00574_),
    .Y(_12797_));
 INVx1_ASAP7_75t_SL _21041_ (.A(_00950_),
    .Y(_12798_));
 NOR2x1_ASAP7_75t_R _21042_ (.A(_00574_),
    .B(_00454_),
    .Y(_12799_));
 INVx1_ASAP7_75t_SL _21043_ (.A(_12799_),
    .Y(_12800_));
 NAND3x1_ASAP7_75t_SL _21044_ (.A(_12797_),
    .B(_12798_),
    .C(_12800_),
    .Y(_12801_));
 AO21x1_ASAP7_75t_SL _21045_ (.A1(_12800_),
    .A2(_12797_),
    .B(_12798_),
    .Y(_12802_));
 NAND2x2_ASAP7_75t_SL _21046_ (.A(_12802_),
    .B(_12801_),
    .Y(_12803_));
 INVx1_ASAP7_75t_R _21048_ (.A(_00633_),
    .Y(_12804_));
 XOR2x2_ASAP7_75t_SL _21049_ (.A(_00600_),
    .B(_00632_),
    .Y(_12805_));
 NAND2x1_ASAP7_75t_R _21050_ (.A(_12804_),
    .B(_12805_),
    .Y(_12806_));
 XNOR2x2_ASAP7_75t_SL _21051_ (.A(_00600_),
    .B(_00632_),
    .Y(_12807_));
 NAND2x1_ASAP7_75t_R _21052_ (.A(_00633_),
    .B(_12807_),
    .Y(_12808_));
 XNOR2x2_ASAP7_75t_SL _21053_ (.A(_00665_),
    .B(_00697_),
    .Y(_12809_));
 AOI21x1_ASAP7_75t_R _21054_ (.A1(_12806_),
    .A2(_12808_),
    .B(_12809_),
    .Y(_12810_));
 NAND2x1_ASAP7_75t_R _21055_ (.A(_00633_),
    .B(_12805_),
    .Y(_12811_));
 NAND2x1_ASAP7_75t_R _21056_ (.A(_12804_),
    .B(_12807_),
    .Y(_12812_));
 XOR2x2_ASAP7_75t_SL _21057_ (.A(_00665_),
    .B(_00697_),
    .Y(_12813_));
 AOI21x1_ASAP7_75t_R _21058_ (.A1(_12811_),
    .A2(_12812_),
    .B(_12813_),
    .Y(_12814_));
 OAI21x1_ASAP7_75t_SL _21059_ (.A1(_12810_),
    .A2(_12814_),
    .B(_00574_),
    .Y(_12815_));
 NOR2x1_ASAP7_75t_R _21060_ (.A(_00574_),
    .B(_00455_),
    .Y(_12816_));
 INVx1_ASAP7_75t_R _21061_ (.A(_12816_),
    .Y(_12817_));
 NAND3x1_ASAP7_75t_SL _21062_ (.A(_12815_),
    .B(_00952_),
    .C(_12817_),
    .Y(_12818_));
 AOI21x1_ASAP7_75t_R _21063_ (.A1(_12817_),
    .A2(_12815_),
    .B(_00952_),
    .Y(_12819_));
 INVx1_ASAP7_75t_SL _21064_ (.A(_12819_),
    .Y(_12820_));
 NAND2x2_ASAP7_75t_SL _21065_ (.A(_12818_),
    .B(_12820_),
    .Y(_12821_));
 INVx5_ASAP7_75t_SL _21067_ (.A(_12803_),
    .Y(_01123_));
 INVx1_ASAP7_75t_R _21068_ (.A(_00952_),
    .Y(_12822_));
 NAND3x1_ASAP7_75t_SL _21069_ (.A(_12815_),
    .B(_12822_),
    .C(_12817_),
    .Y(_12823_));
 INVx1_ASAP7_75t_SL _21070_ (.A(_12815_),
    .Y(_12824_));
 OAI21x1_ASAP7_75t_SL _21071_ (.A1(_12816_),
    .A2(_12824_),
    .B(_00952_),
    .Y(_12825_));
 NAND2x2_ASAP7_75t_SL _21072_ (.A(_12823_),
    .B(_12825_),
    .Y(_12826_));
 NOR2x1_ASAP7_75t_SL _21074_ (.A(_01134_),
    .B(_12821_),
    .Y(_12827_));
 NAND2x1_ASAP7_75t_SL _21075_ (.A(_12821_),
    .B(_12803_),
    .Y(_12828_));
 INVx1_ASAP7_75t_SL _21076_ (.A(_12828_),
    .Y(_12829_));
 XNOR2x2_ASAP7_75t_R _21077_ (.A(_00666_),
    .B(_00698_),
    .Y(_12830_));
 XOR2x2_ASAP7_75t_SL _21078_ (.A(_00633_),
    .B(_00638_),
    .Y(_12831_));
 XOR2x2_ASAP7_75t_SL _21079_ (.A(_12830_),
    .B(_12831_),
    .Y(_12832_));
 XOR2x2_ASAP7_75t_L _21080_ (.A(_00601_),
    .B(_00606_),
    .Y(_12833_));
 XOR2x2_ASAP7_75t_SL _21081_ (.A(_12833_),
    .B(_00634_),
    .Y(_12834_));
 XOR2x2_ASAP7_75t_SL _21082_ (.A(_12832_),
    .B(_12834_),
    .Y(_12835_));
 NOR2x1_ASAP7_75t_R _21083_ (.A(_00574_),
    .B(_00539_),
    .Y(_12836_));
 AOI21x1_ASAP7_75t_SL _21084_ (.A1(_00574_),
    .A2(_12835_),
    .B(_12836_),
    .Y(_12837_));
 XOR2x2_ASAP7_75t_SL _21085_ (.A(_12837_),
    .B(_00953_),
    .Y(_12838_));
 OAI21x1_ASAP7_75t_R _21088_ (.A1(_12827_),
    .A2(_12829_),
    .B(_12838_),
    .Y(_12841_));
 NOR2x1_ASAP7_75t_SL _21089_ (.A(_12821_),
    .B(_12785_),
    .Y(_12842_));
 NOR2x1_ASAP7_75t_SL _21090_ (.A(_12838_),
    .B(_12842_),
    .Y(_12843_));
 NAND2x1_ASAP7_75t_SL _21091_ (.A(_12821_),
    .B(_12785_),
    .Y(_12844_));
 NOR2x1_ASAP7_75t_SL _21092_ (.A(_12803_),
    .B(_12844_),
    .Y(_12845_));
 INVx1_ASAP7_75t_SL _21093_ (.A(_12845_),
    .Y(_12846_));
 XNOR2x2_ASAP7_75t_SL _21094_ (.A(_00634_),
    .B(_00638_),
    .Y(_12847_));
 XOR2x2_ASAP7_75t_L _21095_ (.A(_00667_),
    .B(_00699_),
    .Y(_12848_));
 XOR2x2_ASAP7_75t_R _21096_ (.A(_12847_),
    .B(_12848_),
    .Y(_12849_));
 XOR2x2_ASAP7_75t_R _21097_ (.A(_00602_),
    .B(_00606_),
    .Y(_12850_));
 XOR2x2_ASAP7_75t_SL _21098_ (.A(_12850_),
    .B(_00635_),
    .Y(_12851_));
 XOR2x2_ASAP7_75t_SL _21099_ (.A(_12849_),
    .B(_12851_),
    .Y(_12852_));
 NOR2x1_ASAP7_75t_R _21100_ (.A(_00574_),
    .B(_00538_),
    .Y(_12853_));
 AOI21x1_ASAP7_75t_SL _21101_ (.A1(_00574_),
    .A2(_12852_),
    .B(_12853_),
    .Y(_12854_));
 XNOR2x2_ASAP7_75t_SL _21102_ (.A(_00954_),
    .B(_12854_),
    .Y(_12855_));
 AOI21x1_ASAP7_75t_R _21104_ (.A1(_12843_),
    .A2(_12846_),
    .B(_12855_),
    .Y(_12857_));
 NAND2x1_ASAP7_75t_R _21105_ (.A(_12841_),
    .B(_12857_),
    .Y(_12858_));
 AOI21x1_ASAP7_75t_SL _21106_ (.A1(_12803_),
    .A2(_12785_),
    .B(_12821_),
    .Y(_12859_));
 OAI21x1_ASAP7_75t_SL _21108_ (.A1(_12829_),
    .A2(_12859_),
    .B(_12838_),
    .Y(_12861_));
 AO21x1_ASAP7_75t_R _21109_ (.A1(_12825_),
    .A2(_12823_),
    .B(_01127_),
    .Y(_12862_));
 OAI21x1_ASAP7_75t_R _21110_ (.A1(_12838_),
    .A2(_12862_),
    .B(_12855_),
    .Y(_12863_));
 XNOR2x2_ASAP7_75t_SL _21111_ (.A(_00953_),
    .B(_12837_),
    .Y(_12864_));
 NOR2x2_ASAP7_75t_SL _21113_ (.A(_12826_),
    .B(_12785_),
    .Y(_12866_));
 NAND2x1_ASAP7_75t_SL _21114_ (.A(_12864_),
    .B(_12866_),
    .Y(_12867_));
 INVx1_ASAP7_75t_SL _21115_ (.A(_12867_),
    .Y(_12868_));
 NOR2x1_ASAP7_75t_SL _21116_ (.A(_12863_),
    .B(_12868_),
    .Y(_12869_));
 XOR2x2_ASAP7_75t_SL _21117_ (.A(_00636_),
    .B(_00668_),
    .Y(_12870_));
 XOR2x2_ASAP7_75t_R _21118_ (.A(_12870_),
    .B(_00700_),
    .Y(_12871_));
 XNOR2x2_ASAP7_75t_R _21119_ (.A(_00603_),
    .B(_00635_),
    .Y(_12872_));
 XOR2x2_ASAP7_75t_SL _21120_ (.A(_12871_),
    .B(_12872_),
    .Y(_12873_));
 NOR2x1_ASAP7_75t_SL _21121_ (.A(_00574_),
    .B(_00537_),
    .Y(_12874_));
 AO21x1_ASAP7_75t_R _21122_ (.A1(_12873_),
    .A2(_00574_),
    .B(_12874_),
    .Y(_12875_));
 NOR2x1_ASAP7_75t_R _21123_ (.A(_00955_),
    .B(_12875_),
    .Y(_12876_));
 AND2x2_ASAP7_75t_SL _21124_ (.A(_12875_),
    .B(_00955_),
    .Y(_12877_));
 NOR2x2_ASAP7_75t_SL _21125_ (.A(_12876_),
    .B(_12877_),
    .Y(_12878_));
 INVx1_ASAP7_75t_SL _21126_ (.A(_12878_),
    .Y(_12879_));
 AOI21x1_ASAP7_75t_R _21128_ (.A1(_12861_),
    .A2(_12869_),
    .B(_12879_),
    .Y(_12881_));
 NAND2x1_ASAP7_75t_SL _21129_ (.A(_12858_),
    .B(_12881_),
    .Y(_12882_));
 OAI21x1_ASAP7_75t_R _21131_ (.A1(_12785_),
    .A2(_12826_),
    .B(_01123_),
    .Y(_12884_));
 NAND2x1_ASAP7_75t_SL _21132_ (.A(_12864_),
    .B(_12884_),
    .Y(_12885_));
 INVx1_ASAP7_75t_SL _21135_ (.A(_01134_),
    .Y(_12888_));
 AOI21x1_ASAP7_75t_SL _21136_ (.A1(_12818_),
    .A2(_12820_),
    .B(_12888_),
    .Y(_12889_));
 INVx2_ASAP7_75t_L _21137_ (.A(_12889_),
    .Y(_12890_));
 INVx1_ASAP7_75t_SL _21138_ (.A(_01126_),
    .Y(_12891_));
 AOI21x1_ASAP7_75t_SL _21139_ (.A1(_12823_),
    .A2(_12825_),
    .B(_12891_),
    .Y(_12892_));
 NOR2x2_ASAP7_75t_SL _21140_ (.A(_12864_),
    .B(_12892_),
    .Y(_12893_));
 AOI21x1_ASAP7_75t_SL _21142_ (.A1(_12893_),
    .A2(_12890_),
    .B(_12855_),
    .Y(_12895_));
 AOI21x1_ASAP7_75t_SL _21144_ (.A1(_12885_),
    .A2(_12895_),
    .B(_12878_),
    .Y(_12897_));
 INVx1_ASAP7_75t_R _21146_ (.A(_01129_),
    .Y(_12899_));
 OA21x2_ASAP7_75t_SL _21147_ (.A1(_12899_),
    .A2(_12821_),
    .B(_12838_),
    .Y(_12900_));
 OAI21x1_ASAP7_75t_R _21149_ (.A1(_12803_),
    .A2(_12826_),
    .B(_12864_),
    .Y(_12902_));
 NAND2x1_ASAP7_75t_SL _21150_ (.A(_12855_),
    .B(_12902_),
    .Y(_12903_));
 AO21x1_ASAP7_75t_R _21151_ (.A1(_12900_),
    .A2(_12846_),
    .B(_12903_),
    .Y(_12904_));
 XOR2x2_ASAP7_75t_SL _21152_ (.A(_00604_),
    .B(_00636_),
    .Y(_12905_));
 XOR2x2_ASAP7_75t_R _21153_ (.A(_00637_),
    .B(_00669_),
    .Y(_12906_));
 XOR2x2_ASAP7_75t_R _21154_ (.A(_12906_),
    .B(_00701_),
    .Y(_12907_));
 XNOR2x2_ASAP7_75t_R _21155_ (.A(_12905_),
    .B(_12907_),
    .Y(_12908_));
 NOR2x1_ASAP7_75t_R _21156_ (.A(_00574_),
    .B(_00536_),
    .Y(_12909_));
 AO21x1_ASAP7_75t_R _21157_ (.A1(_12908_),
    .A2(_00574_),
    .B(_12909_),
    .Y(_12910_));
 XOR2x2_ASAP7_75t_SL _21158_ (.A(_12910_),
    .B(_00957_),
    .Y(_12911_));
 AOI21x1_ASAP7_75t_SL _21160_ (.A1(_12904_),
    .A2(_12897_),
    .B(_12911_),
    .Y(_12913_));
 XNOR2x2_ASAP7_75t_R _21161_ (.A(_00638_),
    .B(_00670_),
    .Y(_12914_));
 XOR2x2_ASAP7_75t_R _21162_ (.A(_12914_),
    .B(_00569_),
    .Y(_12915_));
 XOR2x2_ASAP7_75t_R _21163_ (.A(_00605_),
    .B(_00637_),
    .Y(_12916_));
 XOR2x2_ASAP7_75t_SL _21164_ (.A(_12915_),
    .B(_12916_),
    .Y(_12917_));
 NOR2x1_ASAP7_75t_SL _21165_ (.A(_00574_),
    .B(_00535_),
    .Y(_12918_));
 AO21x1_ASAP7_75t_SL _21166_ (.A1(_12917_),
    .A2(_00574_),
    .B(_12918_),
    .Y(_12919_));
 XOR2x2_ASAP7_75t_SL _21167_ (.A(_12919_),
    .B(_00958_),
    .Y(_12920_));
 INVx2_ASAP7_75t_SL _21168_ (.A(_12920_),
    .Y(_12921_));
 AOI21x1_ASAP7_75t_SL _21169_ (.A1(_12913_),
    .A2(_12882_),
    .B(_12921_),
    .Y(_12922_));
 AOI21x1_ASAP7_75t_R _21171_ (.A1(_12785_),
    .A2(_01123_),
    .B(_12864_),
    .Y(_12924_));
 AOI21x1_ASAP7_75t_R _21172_ (.A1(_12828_),
    .A2(_12924_),
    .B(_12855_),
    .Y(_12925_));
 NAND2x1_ASAP7_75t_SL _21173_ (.A(_12785_),
    .B(_01123_),
    .Y(_12926_));
 AO21x1_ASAP7_75t_R _21175_ (.A1(_12926_),
    .A2(_12828_),
    .B(_12838_),
    .Y(_12928_));
 NAND2x1_ASAP7_75t_R _21176_ (.A(_12925_),
    .B(_12928_),
    .Y(_12929_));
 NAND2x1_ASAP7_75t_SL _21177_ (.A(_12803_),
    .B(_12785_),
    .Y(_12930_));
 NOR2x1p5_ASAP7_75t_SL _21178_ (.A(_12838_),
    .B(_12892_),
    .Y(_12931_));
 OAI21x1_ASAP7_75t_SL _21179_ (.A1(_12826_),
    .A2(_12930_),
    .B(_12931_),
    .Y(_12932_));
 INVx2_ASAP7_75t_R _21180_ (.A(_01131_),
    .Y(_12933_));
 AO21x1_ASAP7_75t_R _21181_ (.A1(_12825_),
    .A2(_12823_),
    .B(_12933_),
    .Y(_12934_));
 INVx1_ASAP7_75t_SL _21182_ (.A(_01125_),
    .Y(_12935_));
 AO21x1_ASAP7_75t_SL _21183_ (.A1(_12820_),
    .A2(_12818_),
    .B(_12935_),
    .Y(_12936_));
 NAND2x1_ASAP7_75t_R _21184_ (.A(_12934_),
    .B(_12936_),
    .Y(_12937_));
 XOR2x2_ASAP7_75t_L _21185_ (.A(_12854_),
    .B(_00954_),
    .Y(_12938_));
 AOI21x1_ASAP7_75t_R _21187_ (.A1(_12838_),
    .A2(_12937_),
    .B(_12938_),
    .Y(_12940_));
 AOI21x1_ASAP7_75t_R _21188_ (.A1(_12932_),
    .A2(_12940_),
    .B(_12878_),
    .Y(_12941_));
 NAND2x1_ASAP7_75t_SL _21189_ (.A(_12929_),
    .B(_12941_),
    .Y(_12942_));
 AO21x1_ASAP7_75t_SL _21190_ (.A1(_12820_),
    .A2(_12818_),
    .B(_01125_),
    .Y(_12943_));
 NAND2x1p5_ASAP7_75t_L _21191_ (.A(_12893_),
    .B(_12943_),
    .Y(_12944_));
 NOR2x2_ASAP7_75t_L _21193_ (.A(_12933_),
    .B(_12826_),
    .Y(_12946_));
 AO21x1_ASAP7_75t_SL _21194_ (.A1(_12825_),
    .A2(_12823_),
    .B(_12935_),
    .Y(_12947_));
 INVx1_ASAP7_75t_R _21195_ (.A(_12947_),
    .Y(_12948_));
 OAI21x1_ASAP7_75t_R _21197_ (.A1(_12946_),
    .A2(_12948_),
    .B(_12864_),
    .Y(_12950_));
 AOI21x1_ASAP7_75t_SL _21199_ (.A1(_12950_),
    .A2(_12944_),
    .B(_12938_),
    .Y(_12952_));
 AO21x1_ASAP7_75t_R _21200_ (.A1(_12820_),
    .A2(_12818_),
    .B(_12891_),
    .Y(_12953_));
 AO21x1_ASAP7_75t_R _21202_ (.A1(_12953_),
    .A2(_12838_),
    .B(_12855_),
    .Y(_12955_));
 AND2x2_ASAP7_75t_SL _21203_ (.A(_12892_),
    .B(_12864_),
    .Y(_12956_));
 INVx2_ASAP7_75t_SL _21204_ (.A(_12956_),
    .Y(_12957_));
 NAND2x1_ASAP7_75t_L _21205_ (.A(_12867_),
    .B(_12957_),
    .Y(_12958_));
 NOR2x1_ASAP7_75t_SL _21206_ (.A(_12955_),
    .B(_12958_),
    .Y(_12959_));
 OAI21x1_ASAP7_75t_SL _21208_ (.A1(_12959_),
    .A2(_12952_),
    .B(_12878_),
    .Y(_12961_));
 NAND3x1_ASAP7_75t_SL _21210_ (.A(_12961_),
    .B(_12942_),
    .C(_12911_),
    .Y(_12963_));
 NAND2x1_ASAP7_75t_SL _21211_ (.A(_12922_),
    .B(_12963_),
    .Y(_12964_));
 INVx1_ASAP7_75t_R _21212_ (.A(_12900_),
    .Y(_12965_));
 AO21x1_ASAP7_75t_R _21213_ (.A1(_12936_),
    .A2(_12862_),
    .B(_12838_),
    .Y(_12966_));
 AOI21x1_ASAP7_75t_R _21215_ (.A1(_12965_),
    .A2(_12966_),
    .B(_12855_),
    .Y(_12968_));
 NAND2x2_ASAP7_75t_SL _21216_ (.A(_12826_),
    .B(_12803_),
    .Y(_12969_));
 INVx1_ASAP7_75t_SL _21217_ (.A(_12969_),
    .Y(_12970_));
 OAI21x1_ASAP7_75t_R _21219_ (.A1(_12946_),
    .A2(_12970_),
    .B(_12838_),
    .Y(_12972_));
 AO21x1_ASAP7_75t_R _21220_ (.A1(_12820_),
    .A2(_12818_),
    .B(_01126_),
    .Y(_12973_));
 AOI21x1_ASAP7_75t_SL _21222_ (.A1(_12785_),
    .A2(_12826_),
    .B(_12838_),
    .Y(_12975_));
 NAND2x1_ASAP7_75t_R _21223_ (.A(_12973_),
    .B(_12975_),
    .Y(_12976_));
 AOI21x1_ASAP7_75t_SL _21224_ (.A1(_12972_),
    .A2(_12976_),
    .B(_12938_),
    .Y(_12977_));
 INVx1_ASAP7_75t_SL _21225_ (.A(_12911_),
    .Y(_12978_));
 OAI21x1_ASAP7_75t_R _21226_ (.A1(_12968_),
    .A2(_12977_),
    .B(_12978_),
    .Y(_12979_));
 NAND2x2_ASAP7_75t_SL _21227_ (.A(_12826_),
    .B(_12785_),
    .Y(_12980_));
 INVx1_ASAP7_75t_SL _21228_ (.A(_12980_),
    .Y(_12981_));
 NAND2x1_ASAP7_75t_SL _21229_ (.A(_01123_),
    .B(_12981_),
    .Y(_12982_));
 INVx1_ASAP7_75t_R _21230_ (.A(_01132_),
    .Y(_12983_));
 NOR2x1_ASAP7_75t_SL _21231_ (.A(_12983_),
    .B(_12826_),
    .Y(_12984_));
 NOR2x1_ASAP7_75t_SL _21232_ (.A(_12864_),
    .B(_12984_),
    .Y(_12985_));
 AO21x1_ASAP7_75t_R _21233_ (.A1(_12982_),
    .A2(_12985_),
    .B(_12863_),
    .Y(_12986_));
 OA21x2_ASAP7_75t_R _21235_ (.A1(_12862_),
    .A2(_12864_),
    .B(_12938_),
    .Y(_12988_));
 NOR2x2_ASAP7_75t_SL _21236_ (.A(_01131_),
    .B(_12826_),
    .Y(_12989_));
 NOR2x1_ASAP7_75t_SL _21237_ (.A(_12838_),
    .B(_12989_),
    .Y(_12990_));
 NAND2x1_ASAP7_75t_SL _21238_ (.A(_12990_),
    .B(_12982_),
    .Y(_12991_));
 AOI21x1_ASAP7_75t_R _21239_ (.A1(_12988_),
    .A2(_12991_),
    .B(_12978_),
    .Y(_12992_));
 AOI21x1_ASAP7_75t_R _21240_ (.A1(_12986_),
    .A2(_12992_),
    .B(_12878_),
    .Y(_12993_));
 NAND2x1_ASAP7_75t_R _21241_ (.A(_12979_),
    .B(_12993_),
    .Y(_12994_));
 NOR2x2_ASAP7_75t_SL _21243_ (.A(_01129_),
    .B(_12826_),
    .Y(_12996_));
 AOI21x1_ASAP7_75t_SL _21244_ (.A1(_12864_),
    .A2(_12996_),
    .B(_12938_),
    .Y(_12997_));
 NAND2x1_ASAP7_75t_SL _21245_ (.A(_12997_),
    .B(_12861_),
    .Y(_12998_));
 AOI21x1_ASAP7_75t_SL _21246_ (.A1(_12864_),
    .A2(_12996_),
    .B(_12855_),
    .Y(_12999_));
 AO21x1_ASAP7_75t_R _21247_ (.A1(_12825_),
    .A2(_12823_),
    .B(_01132_),
    .Y(_13000_));
 NOR2x1_ASAP7_75t_R _21249_ (.A(_12838_),
    .B(_13000_),
    .Y(_13002_));
 NOR2x1p5_ASAP7_75t_SL _21250_ (.A(_13002_),
    .B(_12893_),
    .Y(_13003_));
 AOI21x1_ASAP7_75t_SL _21251_ (.A1(_12999_),
    .A2(_13003_),
    .B(_12911_),
    .Y(_13004_));
 NAND2x1_ASAP7_75t_L _21252_ (.A(_12998_),
    .B(_13004_),
    .Y(_13005_));
 OR2x2_ASAP7_75t_R _21253_ (.A(_12864_),
    .B(_01139_),
    .Y(_13006_));
 OA21x2_ASAP7_75t_R _21254_ (.A1(_12973_),
    .A2(_12838_),
    .B(_12938_),
    .Y(_13007_));
 AOI21x1_ASAP7_75t_R _21255_ (.A1(_13006_),
    .A2(_13007_),
    .B(_12978_),
    .Y(_13008_));
 AOI21x1_ASAP7_75t_SL _21256_ (.A1(_12785_),
    .A2(_01123_),
    .B(_12821_),
    .Y(_13009_));
 OAI21x1_ASAP7_75t_SL _21257_ (.A1(_12996_),
    .A2(_13009_),
    .B(_12864_),
    .Y(_13010_));
 NAND2x1_ASAP7_75t_SL _21258_ (.A(_12947_),
    .B(_12828_),
    .Y(_13011_));
 AO21x1_ASAP7_75t_R _21259_ (.A1(_12820_),
    .A2(_12818_),
    .B(_01127_),
    .Y(_13012_));
 OAI21x1_ASAP7_75t_R _21260_ (.A1(_12838_),
    .A2(_13012_),
    .B(_12855_),
    .Y(_13013_));
 AOI21x1_ASAP7_75t_R _21261_ (.A1(_12838_),
    .A2(_13011_),
    .B(_13013_),
    .Y(_13014_));
 NAND2x1_ASAP7_75t_SL _21262_ (.A(_13010_),
    .B(_13014_),
    .Y(_13015_));
 AOI21x1_ASAP7_75t_R _21264_ (.A1(_13008_),
    .A2(_13015_),
    .B(_12879_),
    .Y(_13017_));
 AOI21x1_ASAP7_75t_SL _21266_ (.A1(_13017_),
    .A2(_13005_),
    .B(_12920_),
    .Y(_13019_));
 NAND2x1_ASAP7_75t_SL _21267_ (.A(_12994_),
    .B(_13019_),
    .Y(_13020_));
 NAND2x1_ASAP7_75t_SL _21268_ (.A(_13020_),
    .B(_12964_),
    .Y(_00056_));
 OAI21x1_ASAP7_75t_SL _21269_ (.A1(_12866_),
    .A2(_12829_),
    .B(_12838_),
    .Y(_13021_));
 NOR2x1_ASAP7_75t_SL _21270_ (.A(_12803_),
    .B(_12785_),
    .Y(_13022_));
 INVx1_ASAP7_75t_SL _21271_ (.A(_13022_),
    .Y(_13023_));
 NAND2x1_ASAP7_75t_SL _21272_ (.A(_13023_),
    .B(_12975_),
    .Y(_13024_));
 AOI21x1_ASAP7_75t_SL _21273_ (.A1(_13021_),
    .A2(_13024_),
    .B(_12938_),
    .Y(_13025_));
 AOI21x1_ASAP7_75t_SL _21274_ (.A1(_01129_),
    .A2(_12826_),
    .B(_12838_),
    .Y(_13026_));
 NAND2x1_ASAP7_75t_SL _21275_ (.A(_12828_),
    .B(_13026_),
    .Y(_13027_));
 AOI21x1_ASAP7_75t_R _21276_ (.A1(_12823_),
    .A2(_12825_),
    .B(_01126_),
    .Y(_13028_));
 INVx2_ASAP7_75t_SL _21277_ (.A(_13028_),
    .Y(_13029_));
 AO21x1_ASAP7_75t_SL _21278_ (.A1(_12828_),
    .A2(_13029_),
    .B(_12864_),
    .Y(_13030_));
 AOI21x1_ASAP7_75t_SL _21279_ (.A1(_13027_),
    .A2(_13030_),
    .B(_12855_),
    .Y(_13031_));
 OAI21x1_ASAP7_75t_SL _21280_ (.A1(_13025_),
    .A2(_13031_),
    .B(_12879_),
    .Y(_13032_));
 AOI21x1_ASAP7_75t_SL _21281_ (.A1(_12785_),
    .A2(_12821_),
    .B(_12864_),
    .Y(_13033_));
 NOR2x1_ASAP7_75t_SL _21282_ (.A(_12842_),
    .B(_13033_),
    .Y(_13034_));
 AOI21x1_ASAP7_75t_SL _21283_ (.A1(_12999_),
    .A2(_13034_),
    .B(_12879_),
    .Y(_13035_));
 AO21x1_ASAP7_75t_R _21284_ (.A1(_12825_),
    .A2(_12823_),
    .B(_12888_),
    .Y(_13036_));
 NOR2x2_ASAP7_75t_SL _21285_ (.A(_12891_),
    .B(_12826_),
    .Y(_13037_));
 NOR2x2_ASAP7_75t_SL _21286_ (.A(_12864_),
    .B(_13037_),
    .Y(_13038_));
 AOI21x1_ASAP7_75t_SL _21288_ (.A1(_13036_),
    .A2(_13038_),
    .B(_12938_),
    .Y(_13040_));
 NAND2x1_ASAP7_75t_SL _21289_ (.A(_13010_),
    .B(_13040_),
    .Y(_13041_));
 AOI21x1_ASAP7_75t_SL _21290_ (.A1(_13035_),
    .A2(_13041_),
    .B(_12920_),
    .Y(_13042_));
 AOI21x1_ASAP7_75t_SL _21292_ (.A1(_13032_),
    .A2(_13042_),
    .B(_12978_),
    .Y(_13044_));
 AND3x1_ASAP7_75t_SL _21293_ (.A(_12878_),
    .B(_01141_),
    .C(_12838_),
    .Y(_13045_));
 NAND3x2_ASAP7_75t_SL _21294_ (.B(_12803_),
    .C(_12826_),
    .Y(_13046_),
    .A(_12785_));
 AO21x1_ASAP7_75t_SL _21295_ (.A1(_12990_),
    .A2(_13046_),
    .B(_12938_),
    .Y(_13047_));
 NOR2x1_ASAP7_75t_SL _21296_ (.A(_13045_),
    .B(_13047_),
    .Y(_13048_));
 AND2x2_ASAP7_75t_SL _21297_ (.A(_12969_),
    .B(_12864_),
    .Y(_13049_));
 NAND2x1_ASAP7_75t_SL _21298_ (.A(_12844_),
    .B(_13049_),
    .Y(_13050_));
 INVx1_ASAP7_75t_SL _21299_ (.A(_12866_),
    .Y(_13051_));
 AOI21x1_ASAP7_75t_SL _21300_ (.A1(_13051_),
    .A2(_12900_),
    .B(_12879_),
    .Y(_13052_));
 NAND2x1_ASAP7_75t_SL _21301_ (.A(_13050_),
    .B(_13052_),
    .Y(_13053_));
 NAND2x1_ASAP7_75t_SL _21302_ (.A(_12838_),
    .B(_13046_),
    .Y(_13054_));
 NAND2x1_ASAP7_75t_L _21304_ (.A(_12936_),
    .B(_12969_),
    .Y(_13056_));
 AOI21x1_ASAP7_75t_SL _21305_ (.A1(_12864_),
    .A2(_13056_),
    .B(_12878_),
    .Y(_13057_));
 OAI21x1_ASAP7_75t_SL _21306_ (.A1(_13054_),
    .A2(_12845_),
    .B(_13057_),
    .Y(_13058_));
 AOI21x1_ASAP7_75t_SL _21308_ (.A1(_13053_),
    .A2(_13058_),
    .B(_12855_),
    .Y(_13060_));
 OAI21x1_ASAP7_75t_SL _21309_ (.A1(_13048_),
    .A2(_13060_),
    .B(_12920_),
    .Y(_13061_));
 NAND2x1_ASAP7_75t_SL _21310_ (.A(_13044_),
    .B(_13061_),
    .Y(_13062_));
 OA21x2_ASAP7_75t_SL _21312_ (.A1(_12996_),
    .A2(_12892_),
    .B(_12838_),
    .Y(_13064_));
 AOI211x1_ASAP7_75t_SL _21313_ (.A1(_12864_),
    .A2(_13011_),
    .B(_13064_),
    .C(_12855_),
    .Y(_13065_));
 NAND2x1_ASAP7_75t_SL _21314_ (.A(_12864_),
    .B(_12973_),
    .Y(_13066_));
 NAND2x2_ASAP7_75t_SL _21315_ (.A(_12826_),
    .B(_01123_),
    .Y(_13067_));
 INVx1_ASAP7_75t_SL _21316_ (.A(_13067_),
    .Y(_13068_));
 OA21x2_ASAP7_75t_SL _21317_ (.A1(_13066_),
    .A2(_13068_),
    .B(_12855_),
    .Y(_13069_));
 AO21x1_ASAP7_75t_SL _21318_ (.A1(_13067_),
    .A2(_12930_),
    .B(_12864_),
    .Y(_13070_));
 AO21x1_ASAP7_75t_SL _21320_ (.A1(_13069_),
    .A2(_13070_),
    .B(_12879_),
    .Y(_13072_));
 INVx1_ASAP7_75t_SL _21322_ (.A(_12859_),
    .Y(_13074_));
 AND2x4_ASAP7_75t_SL _21323_ (.A(_12784_),
    .B(_12778_),
    .Y(_01124_));
 NAND2x2_ASAP7_75t_SL _21324_ (.A(_12826_),
    .B(_01124_),
    .Y(_13075_));
 NOR2x1_ASAP7_75t_SL _21325_ (.A(_12889_),
    .B(_12864_),
    .Y(_13076_));
 AOI21x1_ASAP7_75t_SL _21326_ (.A1(_13075_),
    .A2(_13076_),
    .B(_12855_),
    .Y(_13077_));
 OAI21x1_ASAP7_75t_SL _21327_ (.A1(_12838_),
    .A2(_13074_),
    .B(_13077_),
    .Y(_13078_));
 NOR2x1_ASAP7_75t_SL _21328_ (.A(_01129_),
    .B(_12821_),
    .Y(_13079_));
 AOI21x1_ASAP7_75t_SL _21329_ (.A1(_12864_),
    .A2(_13079_),
    .B(_12938_),
    .Y(_13080_));
 AOI21x1_ASAP7_75t_SL _21330_ (.A1(_12803_),
    .A2(_12785_),
    .B(_12826_),
    .Y(_13081_));
 OAI21x1_ASAP7_75t_SL _21331_ (.A1(_12892_),
    .A2(_13081_),
    .B(_12838_),
    .Y(_13082_));
 AOI21x1_ASAP7_75t_SL _21332_ (.A1(_13080_),
    .A2(_13082_),
    .B(_12878_),
    .Y(_13083_));
 AOI21x1_ASAP7_75t_SL _21333_ (.A1(_13078_),
    .A2(_13083_),
    .B(_12920_),
    .Y(_13084_));
 OAI21x1_ASAP7_75t_SL _21334_ (.A1(_13065_),
    .A2(_13072_),
    .B(_13084_),
    .Y(_13085_));
 NOR2x1_ASAP7_75t_SL _21335_ (.A(_12938_),
    .B(_12893_),
    .Y(_13086_));
 OAI21x1_ASAP7_75t_SL _21336_ (.A1(_12829_),
    .A2(_12859_),
    .B(_12864_),
    .Y(_13087_));
 AOI21x1_ASAP7_75t_SL _21337_ (.A1(_13086_),
    .A2(_13087_),
    .B(_12879_),
    .Y(_13088_));
 NAND2x1_ASAP7_75t_R _21338_ (.A(_01127_),
    .B(_12821_),
    .Y(_13089_));
 AND2x2_ASAP7_75t_R _21339_ (.A(_13036_),
    .B(_12864_),
    .Y(_13090_));
 AOI21x1_ASAP7_75t_SL _21340_ (.A1(_13089_),
    .A2(_13090_),
    .B(_12855_),
    .Y(_13091_));
 NAND2x1_ASAP7_75t_SL _21341_ (.A(_13082_),
    .B(_13091_),
    .Y(_13092_));
 AOI21x1_ASAP7_75t_SL _21342_ (.A1(_13088_),
    .A2(_13092_),
    .B(_12921_),
    .Y(_13093_));
 AO21x1_ASAP7_75t_SL _21343_ (.A1(_12973_),
    .A2(_12947_),
    .B(_12864_),
    .Y(_13094_));
 AO21x1_ASAP7_75t_SL _21345_ (.A1(_12828_),
    .A2(_12862_),
    .B(_12838_),
    .Y(_13096_));
 AOI21x1_ASAP7_75t_SL _21346_ (.A1(_13094_),
    .A2(_13096_),
    .B(_12855_),
    .Y(_13097_));
 NAND2x1_ASAP7_75t_SL _21347_ (.A(_13051_),
    .B(_12900_),
    .Y(_13098_));
 AO21x1_ASAP7_75t_SL _21348_ (.A1(_13067_),
    .A2(_12936_),
    .B(_12838_),
    .Y(_13099_));
 AOI21x1_ASAP7_75t_SL _21350_ (.A1(_13098_),
    .A2(_13099_),
    .B(_12938_),
    .Y(_13101_));
 OAI21x1_ASAP7_75t_SL _21351_ (.A1(_13097_),
    .A2(_13101_),
    .B(_12879_),
    .Y(_13102_));
 AOI21x1_ASAP7_75t_SL _21352_ (.A1(_13093_),
    .A2(_13102_),
    .B(_12911_),
    .Y(_13103_));
 NAND2x1_ASAP7_75t_SL _21353_ (.A(_13085_),
    .B(_13103_),
    .Y(_13104_));
 NAND2x1_ASAP7_75t_SL _21354_ (.A(_13062_),
    .B(_13104_),
    .Y(_00057_));
 OA21x2_ASAP7_75t_SL _21355_ (.A1(_13081_),
    .A2(_12827_),
    .B(_12838_),
    .Y(_13105_));
 NOR2x2_ASAP7_75t_SL _21357_ (.A(_12826_),
    .B(_12803_),
    .Y(_13107_));
 AO21x2_ASAP7_75t_SL _21358_ (.A1(_13107_),
    .A2(_12785_),
    .B(_12838_),
    .Y(_13108_));
 NAND2x1_ASAP7_75t_SL _21359_ (.A(_12855_),
    .B(_13108_),
    .Y(_13109_));
 OAI21x1_ASAP7_75t_SL _21360_ (.A1(_13105_),
    .A2(_13109_),
    .B(_12911_),
    .Y(_13110_));
 AO21x1_ASAP7_75t_SL _21361_ (.A1(_13051_),
    .A2(_13029_),
    .B(_12838_),
    .Y(_13111_));
 AO21x1_ASAP7_75t_SL _21362_ (.A1(_12969_),
    .A2(_13012_),
    .B(_12864_),
    .Y(_13112_));
 AND3x1_ASAP7_75t_SL _21363_ (.A(_13111_),
    .B(_12938_),
    .C(_13112_),
    .Y(_13113_));
 NOR2x1_ASAP7_75t_SL _21364_ (.A(_13110_),
    .B(_13113_),
    .Y(_13114_));
 NAND2x1_ASAP7_75t_SL _21365_ (.A(_12973_),
    .B(_12893_),
    .Y(_13115_));
 AO21x1_ASAP7_75t_R _21366_ (.A1(_12820_),
    .A2(_12818_),
    .B(_01132_),
    .Y(_13116_));
 AO21x1_ASAP7_75t_SL _21367_ (.A1(_12969_),
    .A2(_13116_),
    .B(_12838_),
    .Y(_13117_));
 AOI21x1_ASAP7_75t_SL _21368_ (.A1(_13115_),
    .A2(_13117_),
    .B(_12938_),
    .Y(_13118_));
 NOR2x1_ASAP7_75t_SL _21369_ (.A(_12864_),
    .B(_12866_),
    .Y(_13119_));
 OAI21x1_ASAP7_75t_R _21370_ (.A1(_01134_),
    .A2(_12826_),
    .B(_12864_),
    .Y(_13120_));
 OAI21x1_ASAP7_75t_SL _21371_ (.A1(_12970_),
    .A2(_13120_),
    .B(_12938_),
    .Y(_13121_));
 AOI21x1_ASAP7_75t_SL _21372_ (.A1(_13000_),
    .A2(_13119_),
    .B(_13121_),
    .Y(_13122_));
 OAI21x1_ASAP7_75t_SL _21373_ (.A1(_13118_),
    .A2(_13122_),
    .B(_12978_),
    .Y(_13123_));
 NAND2x1_ASAP7_75t_SL _21374_ (.A(_12879_),
    .B(_13123_),
    .Y(_13124_));
 NOR2x1_ASAP7_75t_SL _21375_ (.A(_13114_),
    .B(_13124_),
    .Y(_13125_));
 INVx1_ASAP7_75t_R _21376_ (.A(_13000_),
    .Y(_13126_));
 NOR2x1_ASAP7_75t_SL _21377_ (.A(_01134_),
    .B(_12826_),
    .Y(_13127_));
 OA21x2_ASAP7_75t_SL _21378_ (.A1(_13126_),
    .A2(_13127_),
    .B(_12864_),
    .Y(_13128_));
 AO21x1_ASAP7_75t_SL _21379_ (.A1(_12820_),
    .A2(_12818_),
    .B(_12899_),
    .Y(_13129_));
 AND3x1_ASAP7_75t_SL _21380_ (.A(_13067_),
    .B(_13129_),
    .C(_12838_),
    .Y(_13130_));
 NOR2x1_ASAP7_75t_SL _21381_ (.A(_13128_),
    .B(_13130_),
    .Y(_13131_));
 AND3x1_ASAP7_75t_SL _21382_ (.A(_13075_),
    .B(_13129_),
    .C(_12838_),
    .Y(_13132_));
 OAI21x1_ASAP7_75t_SL _21383_ (.A1(_12838_),
    .A2(_13000_),
    .B(_12997_),
    .Y(_13133_));
 OAI21x1_ASAP7_75t_SL _21384_ (.A1(_13132_),
    .A2(_13133_),
    .B(_12978_),
    .Y(_13134_));
 AOI21x1_ASAP7_75t_SL _21385_ (.A1(_12938_),
    .A2(_13131_),
    .B(_13134_),
    .Y(_13135_));
 OAI21x1_ASAP7_75t_R _21386_ (.A1(_01129_),
    .A2(_12826_),
    .B(_12838_),
    .Y(_13136_));
 NOR2x1_ASAP7_75t_SL _21387_ (.A(_13136_),
    .B(_13009_),
    .Y(_13137_));
 INVx2_ASAP7_75t_R _21388_ (.A(_12973_),
    .Y(_13138_));
 OAI21x1_ASAP7_75t_R _21389_ (.A1(_12821_),
    .A2(_01124_),
    .B(_12864_),
    .Y(_13139_));
 OAI21x1_ASAP7_75t_SL _21390_ (.A1(_13138_),
    .A2(_13139_),
    .B(_12855_),
    .Y(_13140_));
 NOR2x1_ASAP7_75t_SL _21391_ (.A(_13137_),
    .B(_13140_),
    .Y(_13141_));
 NAND2x1_ASAP7_75t_SL _21392_ (.A(_12890_),
    .B(_13026_),
    .Y(_13142_));
 NAND2x1_ASAP7_75t_SL _21393_ (.A(_12980_),
    .B(_12924_),
    .Y(_13143_));
 AOI21x1_ASAP7_75t_SL _21394_ (.A1(_13142_),
    .A2(_13143_),
    .B(_12855_),
    .Y(_13144_));
 OAI21x1_ASAP7_75t_SL _21395_ (.A1(_13141_),
    .A2(_13144_),
    .B(_12911_),
    .Y(_13145_));
 NAND2x1_ASAP7_75t_SL _21396_ (.A(_12878_),
    .B(_13145_),
    .Y(_13146_));
 OAI21x1_ASAP7_75t_SL _21397_ (.A1(_13135_),
    .A2(_13146_),
    .B(_12920_),
    .Y(_13147_));
 INVx1_ASAP7_75t_R _21398_ (.A(_12936_),
    .Y(_13148_));
 NOR2x1_ASAP7_75t_SL _21399_ (.A(_13148_),
    .B(_13139_),
    .Y(_13149_));
 AND3x1_ASAP7_75t_SL _21400_ (.A(_12973_),
    .B(_12934_),
    .C(_12838_),
    .Y(_13150_));
 OAI21x1_ASAP7_75t_SL _21401_ (.A1(_13149_),
    .A2(_13150_),
    .B(_12938_),
    .Y(_13151_));
 NAND2x1_ASAP7_75t_SL _21402_ (.A(_01141_),
    .B(_12864_),
    .Y(_13152_));
 NOR2x1_ASAP7_75t_SL _21403_ (.A(_12864_),
    .B(_13022_),
    .Y(_13153_));
 AOI21x1_ASAP7_75t_SL _21404_ (.A1(_12980_),
    .A2(_13153_),
    .B(_12938_),
    .Y(_13154_));
 AOI21x1_ASAP7_75t_SL _21405_ (.A1(_13152_),
    .A2(_13154_),
    .B(_12911_),
    .Y(_13155_));
 NAND2x1_ASAP7_75t_SL _21406_ (.A(_13151_),
    .B(_13155_),
    .Y(_13156_));
 OA21x2_ASAP7_75t_SL _21407_ (.A1(_12838_),
    .A2(_01143_),
    .B(_12938_),
    .Y(_13157_));
 AOI21x1_ASAP7_75t_SL _21408_ (.A1(_13157_),
    .A2(_13143_),
    .B(_12978_),
    .Y(_13158_));
 NAND2x1_ASAP7_75t_SL _21409_ (.A(_01138_),
    .B(_12838_),
    .Y(_13159_));
 NAND3x1_ASAP7_75t_SL _21410_ (.A(_13108_),
    .B(_12855_),
    .C(_13159_),
    .Y(_13160_));
 AOI21x1_ASAP7_75t_SL _21411_ (.A1(_13158_),
    .A2(_13160_),
    .B(_12879_),
    .Y(_13161_));
 NAND2x1_ASAP7_75t_SL _21412_ (.A(_13156_),
    .B(_13161_),
    .Y(_13162_));
 OA21x2_ASAP7_75t_SL _21413_ (.A1(_12838_),
    .A2(_01139_),
    .B(_12855_),
    .Y(_13163_));
 OAI21x1_ASAP7_75t_SL _21414_ (.A1(_13138_),
    .A2(_13009_),
    .B(_12838_),
    .Y(_13164_));
 AOI21x1_ASAP7_75t_SL _21415_ (.A1(_13163_),
    .A2(_13164_),
    .B(_12911_),
    .Y(_13165_));
 AO21x1_ASAP7_75t_SL _21416_ (.A1(_01124_),
    .A2(_12821_),
    .B(_12864_),
    .Y(_13166_));
 AOI21x1_ASAP7_75t_SL _21417_ (.A1(_12973_),
    .A2(_12975_),
    .B(_12855_),
    .Y(_13167_));
 OAI21x1_ASAP7_75t_SL _21418_ (.A1(_13068_),
    .A2(_13166_),
    .B(_13167_),
    .Y(_13168_));
 NAND2x1_ASAP7_75t_SL _21419_ (.A(_13165_),
    .B(_13168_),
    .Y(_13169_));
 NAND2x1_ASAP7_75t_SL _21420_ (.A(_13129_),
    .B(_12893_),
    .Y(_13170_));
 NOR2x1_ASAP7_75t_SL _21421_ (.A(_12838_),
    .B(_12947_),
    .Y(_13171_));
 NOR2x1_ASAP7_75t_SL _21422_ (.A(_12938_),
    .B(_13171_),
    .Y(_13172_));
 AOI21x1_ASAP7_75t_SL _21423_ (.A1(_13170_),
    .A2(_13172_),
    .B(_12978_),
    .Y(_13173_));
 AND2x4_ASAP7_75t_SL _21424_ (.A(_01129_),
    .B(_01127_),
    .Y(_13174_));
 NOR2x1_ASAP7_75t_L _21425_ (.A(_13174_),
    .B(_12821_),
    .Y(_13175_));
 OAI21x1_ASAP7_75t_SL _21426_ (.A1(_13175_),
    .A2(_13081_),
    .B(_12838_),
    .Y(_13176_));
 AOI21x1_ASAP7_75t_SL _21427_ (.A1(_13046_),
    .A2(_12990_),
    .B(_12855_),
    .Y(_13177_));
 NAND2x1_ASAP7_75t_SL _21428_ (.A(_13176_),
    .B(_13177_),
    .Y(_13178_));
 AOI21x1_ASAP7_75t_SL _21429_ (.A1(_13173_),
    .A2(_13178_),
    .B(_12878_),
    .Y(_13179_));
 AOI21x1_ASAP7_75t_SL _21430_ (.A1(_13169_),
    .A2(_13179_),
    .B(_12920_),
    .Y(_13180_));
 NAND2x1_ASAP7_75t_SL _21431_ (.A(_13162_),
    .B(_13180_),
    .Y(_13181_));
 OAI21x1_ASAP7_75t_SL _21432_ (.A1(_13125_),
    .A2(_13147_),
    .B(_13181_),
    .Y(_00058_));
 INVx1_ASAP7_75t_SL _21433_ (.A(_13175_),
    .Y(_13182_));
 AO21x1_ASAP7_75t_SL _21434_ (.A1(_13116_),
    .A2(_13182_),
    .B(_12864_),
    .Y(_13183_));
 INVx1_ASAP7_75t_R _21435_ (.A(_13183_),
    .Y(_13184_));
 NOR2x1_ASAP7_75t_R _21436_ (.A(_12970_),
    .B(_13120_),
    .Y(_13185_));
 AOI21x1_ASAP7_75t_R _21437_ (.A1(_12938_),
    .A2(_13185_),
    .B(_12879_),
    .Y(_13186_));
 OAI21x1_ASAP7_75t_SL _21438_ (.A1(_13047_),
    .A2(_13184_),
    .B(_13186_),
    .Y(_13187_));
 NAND2x1p5_ASAP7_75t_L _21439_ (.A(_12890_),
    .B(_12931_),
    .Y(_13188_));
 OAI21x1_ASAP7_75t_SL _21440_ (.A1(_13107_),
    .A2(_13126_),
    .B(_12838_),
    .Y(_13189_));
 AOI21x1_ASAP7_75t_R _21441_ (.A1(_13188_),
    .A2(_13189_),
    .B(_12855_),
    .Y(_13190_));
 AO21x1_ASAP7_75t_R _21442_ (.A1(_12828_),
    .A2(_12947_),
    .B(_12864_),
    .Y(_13191_));
 AOI21x1_ASAP7_75t_R _21443_ (.A1(_13024_),
    .A2(_13191_),
    .B(_12938_),
    .Y(_13192_));
 OAI21x1_ASAP7_75t_R _21444_ (.A1(_13190_),
    .A2(_13192_),
    .B(_12879_),
    .Y(_13193_));
 AOI21x1_ASAP7_75t_SL _21445_ (.A1(_13193_),
    .A2(_13187_),
    .B(_12911_),
    .Y(_13194_));
 NOR2x1_ASAP7_75t_SL _21446_ (.A(_12838_),
    .B(_12984_),
    .Y(_13195_));
 NOR2x1_ASAP7_75t_R _21447_ (.A(_12864_),
    .B(_13000_),
    .Y(_13196_));
 AOI21x1_ASAP7_75t_SL _21448_ (.A1(_13067_),
    .A2(_13195_),
    .B(_13196_),
    .Y(_13197_));
 OAI21x1_ASAP7_75t_R _21449_ (.A1(_12878_),
    .A2(_13197_),
    .B(_12855_),
    .Y(_13198_));
 AO21x1_ASAP7_75t_R _21450_ (.A1(_12828_),
    .A2(_13029_),
    .B(_12838_),
    .Y(_13199_));
 AND3x1_ASAP7_75t_L _21451_ (.A(_12820_),
    .B(_12818_),
    .C(_13174_),
    .Y(_13200_));
 OR3x1_ASAP7_75t_L _21452_ (.A(_13200_),
    .B(_12864_),
    .C(_12889_),
    .Y(_13201_));
 AOI21x1_ASAP7_75t_R _21453_ (.A1(_13199_),
    .A2(_13201_),
    .B(_12879_),
    .Y(_13202_));
 NOR2x1_ASAP7_75t_L _21454_ (.A(_13198_),
    .B(_13202_),
    .Y(_13203_));
 OAI21x1_ASAP7_75t_R _21455_ (.A1(_12878_),
    .A2(_12957_),
    .B(_12988_),
    .Y(_13204_));
 AO21x1_ASAP7_75t_R _21456_ (.A1(_12820_),
    .A2(_12818_),
    .B(_01131_),
    .Y(_13205_));
 NAND2x1_ASAP7_75t_R _21457_ (.A(_13205_),
    .B(_12980_),
    .Y(_13206_));
 AOI211x1_ASAP7_75t_R _21458_ (.A1(_13206_),
    .A2(_12864_),
    .B(_12879_),
    .C(_13038_),
    .Y(_13207_));
 OAI21x1_ASAP7_75t_SL _21459_ (.A1(_13207_),
    .A2(_13204_),
    .B(_12911_),
    .Y(_13208_));
 OAI21x1_ASAP7_75t_SL _21460_ (.A1(_13208_),
    .A2(_13203_),
    .B(_12920_),
    .Y(_13209_));
 NOR2x1_ASAP7_75t_SL _21461_ (.A(_13194_),
    .B(_13209_),
    .Y(_13210_));
 OAI21x1_ASAP7_75t_R _21462_ (.A1(_12996_),
    .A2(_12827_),
    .B(_12838_),
    .Y(_13211_));
 NOR2x1_ASAP7_75t_R _21463_ (.A(_13028_),
    .B(_12838_),
    .Y(_13212_));
 AOI21x1_ASAP7_75t_SL _21464_ (.A1(_13212_),
    .A2(_13051_),
    .B(_12938_),
    .Y(_13213_));
 AOI21x1_ASAP7_75t_R _21465_ (.A1(_13211_),
    .A2(_13213_),
    .B(_12878_),
    .Y(_13214_));
 NAND2x1_ASAP7_75t_L _21466_ (.A(_12934_),
    .B(_12828_),
    .Y(_13215_));
 NOR2x1_ASAP7_75t_R _21467_ (.A(_12838_),
    .B(_13215_),
    .Y(_13216_));
 AOI21x1_ASAP7_75t_R _21468_ (.A1(_12838_),
    .A2(_12948_),
    .B(_12855_),
    .Y(_13217_));
 OAI21x1_ASAP7_75t_R _21469_ (.A1(_13038_),
    .A2(_13216_),
    .B(_13217_),
    .Y(_13218_));
 NAND2x1_ASAP7_75t_R _21470_ (.A(_13214_),
    .B(_13218_),
    .Y(_13219_));
 AOI21x1_ASAP7_75t_SL _21471_ (.A1(_13051_),
    .A2(_12893_),
    .B(_12938_),
    .Y(_13220_));
 NAND2x1_ASAP7_75t_R _21472_ (.A(_12926_),
    .B(_13049_),
    .Y(_13221_));
 NAND2x1_ASAP7_75t_SL _21473_ (.A(_13221_),
    .B(_13220_),
    .Y(_13222_));
 AO21x1_ASAP7_75t_R _21474_ (.A1(_12844_),
    .A2(_12969_),
    .B(_12838_),
    .Y(_13223_));
 INVx1_ASAP7_75t_R _21475_ (.A(_12955_),
    .Y(_13224_));
 AOI21x1_ASAP7_75t_R _21476_ (.A1(_13223_),
    .A2(_13224_),
    .B(_12879_),
    .Y(_13225_));
 AOI21x1_ASAP7_75t_SL _21477_ (.A1(_13222_),
    .A2(_13225_),
    .B(_12978_),
    .Y(_13226_));
 NAND2x1_ASAP7_75t_SL _21478_ (.A(_13226_),
    .B(_13219_),
    .Y(_13227_));
 OAI21x1_ASAP7_75t_R _21479_ (.A1(_12859_),
    .A2(_13066_),
    .B(_12855_),
    .Y(_13228_));
 NOR2x1_ASAP7_75t_R _21480_ (.A(_13215_),
    .B(_13166_),
    .Y(_13229_));
 NOR2x1_ASAP7_75t_SL _21481_ (.A(_13228_),
    .B(_13229_),
    .Y(_13230_));
 AOI21x1_ASAP7_75t_R _21482_ (.A1(_12969_),
    .A2(_13023_),
    .B(_12864_),
    .Y(_13231_));
 INVx2_ASAP7_75t_SL _21483_ (.A(_12931_),
    .Y(_13232_));
 OAI21x1_ASAP7_75t_R _21484_ (.A1(_12946_),
    .A2(_13232_),
    .B(_12938_),
    .Y(_13233_));
 OAI21x1_ASAP7_75t_SL _21485_ (.A1(_13233_),
    .A2(_13231_),
    .B(_12879_),
    .Y(_13234_));
 NOR2x1_ASAP7_75t_SL _21486_ (.A(_13230_),
    .B(_13234_),
    .Y(_13235_));
 OAI21x1_ASAP7_75t_R _21487_ (.A1(_12826_),
    .A2(_01123_),
    .B(_12855_),
    .Y(_13236_));
 NOR2x1_ASAP7_75t_SL _21488_ (.A(_13022_),
    .B(_13236_),
    .Y(_13237_));
 OAI21x1_ASAP7_75t_R _21489_ (.A1(_12821_),
    .A2(_12864_),
    .B(_13237_),
    .Y(_13238_));
 INVx1_ASAP7_75t_R _21490_ (.A(_13212_),
    .Y(_13239_));
 OAI21x1_ASAP7_75t_R _21491_ (.A1(_12984_),
    .A2(_13239_),
    .B(_13077_),
    .Y(_13240_));
 AOI21x1_ASAP7_75t_R _21492_ (.A1(_13238_),
    .A2(_13240_),
    .B(_12879_),
    .Y(_13241_));
 OAI21x1_ASAP7_75t_SL _21493_ (.A1(_13241_),
    .A2(_13235_),
    .B(_12978_),
    .Y(_13242_));
 AOI21x1_ASAP7_75t_SL _21494_ (.A1(_13227_),
    .A2(_13242_),
    .B(_12920_),
    .Y(_13243_));
 NOR2x1_ASAP7_75t_SL _21495_ (.A(_13210_),
    .B(_13243_),
    .Y(_00059_));
 AO21x1_ASAP7_75t_SL _21496_ (.A1(_13154_),
    .A2(_13050_),
    .B(_12879_),
    .Y(_13244_));
 AND3x1_ASAP7_75t_SL _21497_ (.A(_13075_),
    .B(_12943_),
    .C(_12838_),
    .Y(_13245_));
 AOI211x1_ASAP7_75t_SL _21498_ (.A1(_12930_),
    .A2(_12843_),
    .B(_13245_),
    .C(_12855_),
    .Y(_13246_));
 NAND2x1_ASAP7_75t_SL _21499_ (.A(_12938_),
    .B(_12862_),
    .Y(_13247_));
 OA21x2_ASAP7_75t_SL _21500_ (.A1(_12985_),
    .A2(_13247_),
    .B(_12879_),
    .Y(_13248_));
 NAND2x1_ASAP7_75t_SL _21501_ (.A(_13067_),
    .B(_13033_),
    .Y(_13249_));
 AOI21x1_ASAP7_75t_SL _21502_ (.A1(_12864_),
    .A2(_13056_),
    .B(_12938_),
    .Y(_13250_));
 NAND2x1_ASAP7_75t_SL _21503_ (.A(_13249_),
    .B(_13250_),
    .Y(_13251_));
 AOI21x1_ASAP7_75t_SL _21504_ (.A1(_13248_),
    .A2(_13251_),
    .B(_12911_),
    .Y(_13252_));
 OAI21x1_ASAP7_75t_SL _21505_ (.A1(_13244_),
    .A2(_13246_),
    .B(_13252_),
    .Y(_13253_));
 OA21x2_ASAP7_75t_SL _21506_ (.A1(_12973_),
    .A2(_12864_),
    .B(_13000_),
    .Y(_13254_));
 AOI21x1_ASAP7_75t_SL _21507_ (.A1(_12999_),
    .A2(_13254_),
    .B(_12878_),
    .Y(_13255_));
 NAND2x1_ASAP7_75t_SL _21508_ (.A(_12985_),
    .B(_12982_),
    .Y(_13256_));
 AOI21x1_ASAP7_75t_SL _21509_ (.A1(_12953_),
    .A2(_13090_),
    .B(_12938_),
    .Y(_13257_));
 NAND2x1_ASAP7_75t_SL _21510_ (.A(_13256_),
    .B(_13257_),
    .Y(_13258_));
 AOI21x1_ASAP7_75t_SL _21511_ (.A1(_13255_),
    .A2(_13258_),
    .B(_12978_),
    .Y(_13259_));
 INVx1_ASAP7_75t_R _21512_ (.A(_12844_),
    .Y(_13260_));
 OAI21x1_ASAP7_75t_SL _21513_ (.A1(_13260_),
    .A2(_13009_),
    .B(_12838_),
    .Y(_13261_));
 AOI21x1_ASAP7_75t_SL _21514_ (.A1(_13142_),
    .A2(_13261_),
    .B(_12855_),
    .Y(_13262_));
 AO21x1_ASAP7_75t_SL _21515_ (.A1(_12844_),
    .A2(_12947_),
    .B(_12864_),
    .Y(_13263_));
 AOI21x1_ASAP7_75t_SL _21516_ (.A1(_13263_),
    .A2(_13010_),
    .B(_12938_),
    .Y(_13264_));
 OAI21x1_ASAP7_75t_SL _21517_ (.A1(_13262_),
    .A2(_13264_),
    .B(_12878_),
    .Y(_13265_));
 AOI21x1_ASAP7_75t_SL _21518_ (.A1(_13259_),
    .A2(_13265_),
    .B(_12920_),
    .Y(_13266_));
 NAND2x1_ASAP7_75t_SL _21519_ (.A(_13253_),
    .B(_13266_),
    .Y(_13267_));
 NAND2x1_ASAP7_75t_R _21520_ (.A(_12821_),
    .B(_12838_),
    .Y(_13268_));
 AND2x2_ASAP7_75t_SL _21521_ (.A(_13268_),
    .B(_12855_),
    .Y(_13269_));
 NAND2x1_ASAP7_75t_SL _21522_ (.A(_12890_),
    .B(_13049_),
    .Y(_13270_));
 AOI21x1_ASAP7_75t_SL _21523_ (.A1(_13269_),
    .A2(_13270_),
    .B(_12879_),
    .Y(_13271_));
 NOR2x1_ASAP7_75t_SL _21524_ (.A(_12855_),
    .B(_13171_),
    .Y(_13272_));
 NAND3x1_ASAP7_75t_SL _21525_ (.A(_13098_),
    .B(_12867_),
    .C(_13272_),
    .Y(_13273_));
 AOI21x1_ASAP7_75t_SL _21526_ (.A1(_13271_),
    .A2(_13273_),
    .B(_12911_),
    .Y(_13274_));
 AND2x2_ASAP7_75t_SL _21527_ (.A(_13026_),
    .B(_12973_),
    .Y(_13275_));
 NOR2x1_ASAP7_75t_SL _21528_ (.A(_12938_),
    .B(_13275_),
    .Y(_13276_));
 AO21x1_ASAP7_75t_SL _21529_ (.A1(_13089_),
    .A2(_12864_),
    .B(_12855_),
    .Y(_13277_));
 NOR2x1_ASAP7_75t_R _21530_ (.A(_01123_),
    .B(_12844_),
    .Y(_13278_));
 NOR2x1_ASAP7_75t_SL _21531_ (.A(_12864_),
    .B(_13278_),
    .Y(_13279_));
 OAI21x1_ASAP7_75t_SL _21532_ (.A1(_13277_),
    .A2(_13279_),
    .B(_12879_),
    .Y(_13280_));
 AO21x1_ASAP7_75t_SL _21533_ (.A1(_12861_),
    .A2(_13276_),
    .B(_13280_),
    .Y(_13281_));
 NAND2x1_ASAP7_75t_SL _21534_ (.A(_13274_),
    .B(_13281_),
    .Y(_13282_));
 NAND2x1_ASAP7_75t_SL _21535_ (.A(_12864_),
    .B(_13009_),
    .Y(_13283_));
 AOI21x1_ASAP7_75t_SL _21536_ (.A1(_13075_),
    .A2(_12985_),
    .B(_12855_),
    .Y(_13284_));
 NAND2x1_ASAP7_75t_SL _21537_ (.A(_13283_),
    .B(_13284_),
    .Y(_13285_));
 NOR2x1_ASAP7_75t_R _21538_ (.A(_01133_),
    .B(_12838_),
    .Y(_13286_));
 AO21x1_ASAP7_75t_SL _21539_ (.A1(_13138_),
    .A2(_12838_),
    .B(_13286_),
    .Y(_13287_));
 AOI21x1_ASAP7_75t_SL _21540_ (.A1(_12855_),
    .A2(_13287_),
    .B(_12878_),
    .Y(_13288_));
 AOI21x1_ASAP7_75t_SL _21541_ (.A1(_13285_),
    .A2(_13288_),
    .B(_12978_),
    .Y(_13289_));
 NAND2x1_ASAP7_75t_SL _21542_ (.A(_12930_),
    .B(_12843_),
    .Y(_13290_));
 AO21x1_ASAP7_75t_R _21543_ (.A1(_12820_),
    .A2(_12818_),
    .B(_12983_),
    .Y(_13291_));
 AO21x1_ASAP7_75t_SL _21544_ (.A1(_12969_),
    .A2(_13291_),
    .B(_12864_),
    .Y(_13292_));
 AO21x1_ASAP7_75t_SL _21545_ (.A1(_13290_),
    .A2(_13292_),
    .B(_12855_),
    .Y(_13293_));
 INVx1_ASAP7_75t_SL _21546_ (.A(_13231_),
    .Y(_13294_));
 AOI21x1_ASAP7_75t_SL _21547_ (.A1(_12864_),
    .A2(_13148_),
    .B(_12863_),
    .Y(_13295_));
 AOI21x1_ASAP7_75t_SL _21548_ (.A1(_13294_),
    .A2(_13295_),
    .B(_12879_),
    .Y(_13296_));
 NAND2x1_ASAP7_75t_SL _21549_ (.A(_13293_),
    .B(_13296_),
    .Y(_13297_));
 AOI21x1_ASAP7_75t_SL _21550_ (.A1(_13289_),
    .A2(_13297_),
    .B(_12921_),
    .Y(_13298_));
 NAND2x1_ASAP7_75t_SL _21551_ (.A(_13282_),
    .B(_13298_),
    .Y(_13299_));
 NAND2x1_ASAP7_75t_SL _21552_ (.A(_13267_),
    .B(_13299_),
    .Y(_00060_));
 AND2x2_ASAP7_75t_L _21553_ (.A(_12893_),
    .B(_13205_),
    .Y(_13300_));
 AO21x1_ASAP7_75t_R _21554_ (.A1(_13212_),
    .A2(_12890_),
    .B(_12855_),
    .Y(_13301_));
 OA21x2_ASAP7_75t_R _21555_ (.A1(_12864_),
    .A2(_12933_),
    .B(_12855_),
    .Y(_13302_));
 NAND2x1_ASAP7_75t_SL _21556_ (.A(_12864_),
    .B(_13046_),
    .Y(_13303_));
 AOI21x1_ASAP7_75t_R _21557_ (.A1(_13302_),
    .A2(_13303_),
    .B(_12879_),
    .Y(_13304_));
 OAI21x1_ASAP7_75t_R _21558_ (.A1(_13300_),
    .A2(_13301_),
    .B(_13304_),
    .Y(_13305_));
 INVx1_ASAP7_75t_R _21559_ (.A(_13076_),
    .Y(_13306_));
 AOI21x1_ASAP7_75t_R _21560_ (.A1(_13306_),
    .A2(_12999_),
    .B(_12878_),
    .Y(_13307_));
 INVx1_ASAP7_75t_R _21561_ (.A(_13046_),
    .Y(_13308_));
 OA21x2_ASAP7_75t_R _21562_ (.A1(_13200_),
    .A2(_12864_),
    .B(_12855_),
    .Y(_13309_));
 OAI21x1_ASAP7_75t_R _21563_ (.A1(_13308_),
    .A2(_13108_),
    .B(_13309_),
    .Y(_13310_));
 AOI21x1_ASAP7_75t_R _21564_ (.A1(_13307_),
    .A2(_13310_),
    .B(_12978_),
    .Y(_13311_));
 AOI21x1_ASAP7_75t_R _21565_ (.A1(_13305_),
    .A2(_13311_),
    .B(_12921_),
    .Y(_13312_));
 NOR2x1_ASAP7_75t_L _21566_ (.A(_12838_),
    .B(_12969_),
    .Y(_13313_));
 NOR2x1_ASAP7_75t_R _21567_ (.A(_13313_),
    .B(_12998_),
    .Y(_13314_));
 AO21x1_ASAP7_75t_R _21568_ (.A1(_12946_),
    .A2(_12838_),
    .B(_12855_),
    .Y(_13315_));
 NOR2x1_ASAP7_75t_R _21569_ (.A(_12889_),
    .B(_13303_),
    .Y(_13316_));
 OAI21x1_ASAP7_75t_R _21570_ (.A1(_13315_),
    .A2(_13316_),
    .B(_12878_),
    .Y(_13317_));
 INVx2_ASAP7_75t_R _21571_ (.A(_12893_),
    .Y(_13318_));
 AOI21x1_ASAP7_75t_R _21572_ (.A1(_13075_),
    .A2(_13195_),
    .B(_12855_),
    .Y(_13319_));
 OAI21x1_ASAP7_75t_R _21573_ (.A1(_13318_),
    .A2(_12845_),
    .B(_13319_),
    .Y(_13320_));
 OA21x2_ASAP7_75t_R _21574_ (.A1(_01123_),
    .A2(_12864_),
    .B(_12855_),
    .Y(_13321_));
 AOI21x1_ASAP7_75t_R _21575_ (.A1(_13321_),
    .A2(_12928_),
    .B(_12878_),
    .Y(_13322_));
 AOI21x1_ASAP7_75t_R _21576_ (.A1(_13320_),
    .A2(_13322_),
    .B(_12911_),
    .Y(_13323_));
 OAI21x1_ASAP7_75t_R _21577_ (.A1(_13314_),
    .A2(_13317_),
    .B(_13323_),
    .Y(_13324_));
 NAND2x1_ASAP7_75t_SL _21578_ (.A(_13312_),
    .B(_13324_),
    .Y(_13325_));
 NAND2x1_ASAP7_75t_R _21579_ (.A(_12785_),
    .B(_12838_),
    .Y(_13326_));
 AOI21x1_ASAP7_75t_R _21580_ (.A1(_13326_),
    .A2(_13290_),
    .B(_12938_),
    .Y(_13327_));
 INVx1_ASAP7_75t_L _21581_ (.A(_12930_),
    .Y(_13328_));
 OAI21x1_ASAP7_75t_R _21582_ (.A1(_13328_),
    .A2(_12902_),
    .B(_12938_),
    .Y(_13329_));
 AOI21x1_ASAP7_75t_R _21583_ (.A1(_13205_),
    .A2(_13046_),
    .B(_12864_),
    .Y(_13330_));
 OAI21x1_ASAP7_75t_R _21584_ (.A1(_13329_),
    .A2(_13330_),
    .B(_12879_),
    .Y(_13331_));
 NOR2x1_ASAP7_75t_SL _21585_ (.A(_13327_),
    .B(_13331_),
    .Y(_13332_));
 NAND2x1_ASAP7_75t_R _21586_ (.A(_12838_),
    .B(_13138_),
    .Y(_13333_));
 AO21x1_ASAP7_75t_R _21587_ (.A1(_13075_),
    .A2(_13012_),
    .B(_12838_),
    .Y(_13334_));
 AOI21x1_ASAP7_75t_R _21588_ (.A1(_13333_),
    .A2(_13334_),
    .B(_12855_),
    .Y(_13335_));
 AND2x2_ASAP7_75t_SL _21589_ (.A(_13120_),
    .B(_12855_),
    .Y(_13336_));
 NAND2x1p5_ASAP7_75t_L _21590_ (.A(_12936_),
    .B(_12893_),
    .Y(_13337_));
 AO21x1_ASAP7_75t_R _21591_ (.A1(_13337_),
    .A2(_13336_),
    .B(_12879_),
    .Y(_13338_));
 NOR2x1_ASAP7_75t_L _21592_ (.A(_13335_),
    .B(_13338_),
    .Y(_13339_));
 OAI21x1_ASAP7_75t_R _21593_ (.A1(_13332_),
    .A2(_13339_),
    .B(_12911_),
    .Y(_13340_));
 AOI21x1_ASAP7_75t_R _21594_ (.A1(_13232_),
    .A2(_13189_),
    .B(_12938_),
    .Y(_13341_));
 INVx1_ASAP7_75t_R _21595_ (.A(_13026_),
    .Y(_13342_));
 AOI21x1_ASAP7_75t_R _21596_ (.A1(_13342_),
    .A2(_13021_),
    .B(_12855_),
    .Y(_13343_));
 OAI21x1_ASAP7_75t_R _21597_ (.A1(_13341_),
    .A2(_13343_),
    .B(_12878_),
    .Y(_13344_));
 OAI21x1_ASAP7_75t_R _21598_ (.A1(_13127_),
    .A2(_13079_),
    .B(_12838_),
    .Y(_13345_));
 NAND2x1_ASAP7_75t_SL _21599_ (.A(_13345_),
    .B(_12869_),
    .Y(_13346_));
 NOR2x1_ASAP7_75t_R _21600_ (.A(_13174_),
    .B(_12864_),
    .Y(_13347_));
 AOI21x1_ASAP7_75t_R _21601_ (.A1(_13129_),
    .A2(_13347_),
    .B(_12855_),
    .Y(_13348_));
 NAND2x1_ASAP7_75t_SL _21602_ (.A(_13195_),
    .B(_12982_),
    .Y(_13349_));
 AOI21x1_ASAP7_75t_SL _21603_ (.A1(_13348_),
    .A2(_13349_),
    .B(_12878_),
    .Y(_13350_));
 AOI21x1_ASAP7_75t_R _21604_ (.A1(_13346_),
    .A2(_13350_),
    .B(_12911_),
    .Y(_13351_));
 AOI21x1_ASAP7_75t_R _21605_ (.A1(_13344_),
    .A2(_13351_),
    .B(_12920_),
    .Y(_13352_));
 NAND2x1_ASAP7_75t_SL _21606_ (.A(_13340_),
    .B(_13352_),
    .Y(_13353_));
 NAND2x1_ASAP7_75t_SL _21607_ (.A(_13325_),
    .B(_13353_),
    .Y(_00061_));
 AO21x1_ASAP7_75t_SL _21608_ (.A1(_13108_),
    .A2(_13159_),
    .B(_12956_),
    .Y(_13354_));
 AO21x1_ASAP7_75t_R _21609_ (.A1(_01124_),
    .A2(_12826_),
    .B(_12864_),
    .Y(_13355_));
 NOR2x1_ASAP7_75t_SL _21610_ (.A(_12845_),
    .B(_13355_),
    .Y(_13356_));
 AO21x1_ASAP7_75t_SL _21611_ (.A1(_13212_),
    .A2(_13089_),
    .B(_12938_),
    .Y(_13357_));
 OAI21x1_ASAP7_75t_SL _21612_ (.A1(_13356_),
    .A2(_13357_),
    .B(_12879_),
    .Y(_13358_));
 AOI21x1_ASAP7_75t_SL _21613_ (.A1(_12938_),
    .A2(_13354_),
    .B(_13358_),
    .Y(_13359_));
 AO21x1_ASAP7_75t_SL _21614_ (.A1(_12946_),
    .A2(_12864_),
    .B(_12855_),
    .Y(_13360_));
 AND2x2_ASAP7_75t_SL _21615_ (.A(_13033_),
    .B(_12926_),
    .Y(_13361_));
 OAI21x1_ASAP7_75t_SL _21616_ (.A1(_13360_),
    .A2(_13361_),
    .B(_12878_),
    .Y(_13362_));
 NOR2x1_ASAP7_75t_SL _21617_ (.A(_12803_),
    .B(_12980_),
    .Y(_13363_));
 NOR2x1_ASAP7_75t_SL _21618_ (.A(_12864_),
    .B(_13363_),
    .Y(_13364_));
 AOI21x1_ASAP7_75t_R _21619_ (.A1(_12864_),
    .A2(_13037_),
    .B(_12938_),
    .Y(_13365_));
 OAI21x1_ASAP7_75t_SL _21620_ (.A1(_12838_),
    .A2(_13182_),
    .B(_13365_),
    .Y(_13366_));
 AOI21x1_ASAP7_75t_SL _21621_ (.A1(_12828_),
    .A2(_13364_),
    .B(_13366_),
    .Y(_13367_));
 OAI21x1_ASAP7_75t_SL _21622_ (.A1(_13362_),
    .A2(_13367_),
    .B(_12911_),
    .Y(_13368_));
 OAI21x1_ASAP7_75t_SL _21623_ (.A1(_13359_),
    .A2(_13368_),
    .B(_12921_),
    .Y(_13369_));
 NAND2x1_ASAP7_75t_SL _21624_ (.A(_12926_),
    .B(_13119_),
    .Y(_13370_));
 AO21x1_ASAP7_75t_R _21625_ (.A1(_01142_),
    .A2(_01136_),
    .B(_12838_),
    .Y(_13371_));
 AND2x2_ASAP7_75t_SL _21626_ (.A(_13371_),
    .B(_12855_),
    .Y(_13372_));
 NAND2x1_ASAP7_75t_SL _21627_ (.A(_13370_),
    .B(_13372_),
    .Y(_13373_));
 AO21x1_ASAP7_75t_SL _21628_ (.A1(_13012_),
    .A2(_13000_),
    .B(_12864_),
    .Y(_13374_));
 NAND2x1_ASAP7_75t_SL _21629_ (.A(_13374_),
    .B(_13272_),
    .Y(_13375_));
 AO21x1_ASAP7_75t_SL _21630_ (.A1(_13373_),
    .A2(_13375_),
    .B(_12878_),
    .Y(_13376_));
 AND3x1_ASAP7_75t_SL _21631_ (.A(_13291_),
    .B(_13036_),
    .C(_12864_),
    .Y(_13377_));
 OAI22x1_ASAP7_75t_SL _21632_ (.A1(_13328_),
    .A2(_13268_),
    .B1(_12864_),
    .B2(_12862_),
    .Y(_13378_));
 OAI21x1_ASAP7_75t_SL _21633_ (.A1(_13377_),
    .A2(_13378_),
    .B(_12855_),
    .Y(_13379_));
 NOR2x1_ASAP7_75t_SL _21634_ (.A(_01127_),
    .B(_12826_),
    .Y(_13380_));
 OR3x1_ASAP7_75t_SL _21635_ (.A(_13136_),
    .B(_13126_),
    .C(_13380_),
    .Y(_13381_));
 AOI211x1_ASAP7_75t_SL _21636_ (.A1(_13138_),
    .A2(_12864_),
    .B(_13313_),
    .C(_12855_),
    .Y(_13382_));
 AOI21x1_ASAP7_75t_SL _21637_ (.A1(_13381_),
    .A2(_13382_),
    .B(_12879_),
    .Y(_13383_));
 NAND2x1_ASAP7_75t_SL _21638_ (.A(_13379_),
    .B(_13383_),
    .Y(_13384_));
 AOI21x1_ASAP7_75t_SL _21639_ (.A1(_13376_),
    .A2(_13384_),
    .B(_12911_),
    .Y(_13385_));
 AO21x1_ASAP7_75t_SL _21640_ (.A1(_12829_),
    .A2(_12864_),
    .B(_12855_),
    .Y(_13386_));
 AND2x2_ASAP7_75t_SL _21641_ (.A(_13076_),
    .B(_13029_),
    .Y(_13387_));
 AOI21x1_ASAP7_75t_SL _21642_ (.A1(_01137_),
    .A2(_12838_),
    .B(_12938_),
    .Y(_13388_));
 NAND2x1_ASAP7_75t_SL _21643_ (.A(_13075_),
    .B(_13195_),
    .Y(_13389_));
 AOI21x1_ASAP7_75t_SL _21644_ (.A1(_13388_),
    .A2(_13389_),
    .B(_12878_),
    .Y(_13390_));
 OAI21x1_ASAP7_75t_SL _21645_ (.A1(_13386_),
    .A2(_13387_),
    .B(_13390_),
    .Y(_13391_));
 AOI21x1_ASAP7_75t_SL _21646_ (.A1(_12855_),
    .A2(_13137_),
    .B(_12879_),
    .Y(_13392_));
 OAI21x1_ASAP7_75t_SL _21647_ (.A1(_12838_),
    .A2(_12989_),
    .B(_13284_),
    .Y(_13393_));
 AOI21x1_ASAP7_75t_SL _21648_ (.A1(_13392_),
    .A2(_13393_),
    .B(_12978_),
    .Y(_13394_));
 NAND2x1_ASAP7_75t_SL _21649_ (.A(_13391_),
    .B(_13394_),
    .Y(_13395_));
 NOR2x1_ASAP7_75t_SL _21650_ (.A(_12855_),
    .B(_13033_),
    .Y(_13396_));
 NAND2x1_ASAP7_75t_SL _21651_ (.A(_12885_),
    .B(_13396_),
    .Y(_13397_));
 OA21x2_ASAP7_75t_SL _21652_ (.A1(_13029_),
    .A2(_12838_),
    .B(_12855_),
    .Y(_13398_));
 AOI21x1_ASAP7_75t_SL _21653_ (.A1(_13189_),
    .A2(_13398_),
    .B(_12879_),
    .Y(_13399_));
 AOI21x1_ASAP7_75t_SL _21654_ (.A1(_13397_),
    .A2(_13399_),
    .B(_12911_),
    .Y(_13400_));
 OA21x2_ASAP7_75t_SL _21655_ (.A1(_13090_),
    .A2(_13153_),
    .B(_12828_),
    .Y(_13401_));
 NAND2x1_ASAP7_75t_SL _21656_ (.A(_12864_),
    .B(_01124_),
    .Y(_13402_));
 AOI21x1_ASAP7_75t_SL _21657_ (.A1(_13402_),
    .A2(_13237_),
    .B(_12878_),
    .Y(_13403_));
 OAI21x1_ASAP7_75t_SL _21658_ (.A1(_12855_),
    .A2(_13401_),
    .B(_13403_),
    .Y(_13404_));
 AOI21x1_ASAP7_75t_SL _21659_ (.A1(_13400_),
    .A2(_13404_),
    .B(_12921_),
    .Y(_13405_));
 NAND2x1_ASAP7_75t_SL _21660_ (.A(_13395_),
    .B(_13405_),
    .Y(_13406_));
 OAI21x1_ASAP7_75t_SL _21661_ (.A1(_13369_),
    .A2(_13385_),
    .B(_13406_),
    .Y(_00062_));
 NOR2x1_ASAP7_75t_R _21662_ (.A(_12803_),
    .B(_12838_),
    .Y(_13407_));
 AOI21x1_ASAP7_75t_R _21663_ (.A1(_13067_),
    .A2(_13033_),
    .B(_13407_),
    .Y(_13408_));
 OAI21x1_ASAP7_75t_R _21664_ (.A1(_12855_),
    .A2(_13408_),
    .B(_12879_),
    .Y(_13409_));
 OA21x2_ASAP7_75t_R _21665_ (.A1(_13081_),
    .A2(_12981_),
    .B(_12864_),
    .Y(_13410_));
 INVx1_ASAP7_75t_R _21666_ (.A(_13154_),
    .Y(_13411_));
 NOR2x1_ASAP7_75t_SL _21667_ (.A(_13410_),
    .B(_13411_),
    .Y(_13412_));
 NOR2x1_ASAP7_75t_R _21668_ (.A(_13239_),
    .B(_13278_),
    .Y(_13413_));
 OAI21x1_ASAP7_75t_R _21669_ (.A1(_12864_),
    .A2(_13363_),
    .B(_12938_),
    .Y(_13414_));
 AOI21x1_ASAP7_75t_R _21670_ (.A1(_12864_),
    .A2(_12892_),
    .B(_12938_),
    .Y(_13415_));
 NAND2x1_ASAP7_75t_R _21671_ (.A(_12838_),
    .B(_12859_),
    .Y(_13416_));
 AOI21x1_ASAP7_75t_R _21672_ (.A1(_13415_),
    .A2(_13416_),
    .B(_12879_),
    .Y(_13417_));
 OAI21x1_ASAP7_75t_SL _21673_ (.A1(_13413_),
    .A2(_13414_),
    .B(_13417_),
    .Y(_13418_));
 OAI21x1_ASAP7_75t_R _21674_ (.A1(_13409_),
    .A2(_13412_),
    .B(_13418_),
    .Y(_13419_));
 OAI21x1_ASAP7_75t_R _21675_ (.A1(_12978_),
    .A2(_13419_),
    .B(_12920_),
    .Y(_13420_));
 NAND2x1_ASAP7_75t_R _21676_ (.A(_13036_),
    .B(_13038_),
    .Y(_13421_));
 AND3x1_ASAP7_75t_SL _21677_ (.A(_13421_),
    .B(_13199_),
    .C(_12938_),
    .Y(_13422_));
 OAI21x1_ASAP7_75t_R _21678_ (.A1(_13068_),
    .A2(_13166_),
    .B(_12855_),
    .Y(_13423_));
 OAI21x1_ASAP7_75t_R _21679_ (.A1(_13377_),
    .A2(_13423_),
    .B(_12878_),
    .Y(_13424_));
 NOR2x1_ASAP7_75t_R _21680_ (.A(_13422_),
    .B(_13424_),
    .Y(_13425_));
 AO21x1_ASAP7_75t_R _21681_ (.A1(_13036_),
    .A2(_12864_),
    .B(_12938_),
    .Y(_13426_));
 AND2x2_ASAP7_75t_R _21682_ (.A(_12985_),
    .B(_13075_),
    .Y(_13427_));
 OAI21x1_ASAP7_75t_R _21683_ (.A1(_13426_),
    .A2(_13427_),
    .B(_12879_),
    .Y(_13428_));
 NOR2x1_ASAP7_75t_R _21684_ (.A(_12902_),
    .B(_13363_),
    .Y(_13429_));
 OAI21x1_ASAP7_75t_R _21685_ (.A1(_13268_),
    .A2(_13328_),
    .B(_13217_),
    .Y(_13430_));
 NOR2x1_ASAP7_75t_SL _21686_ (.A(_13429_),
    .B(_13430_),
    .Y(_13431_));
 NOR2x1_ASAP7_75t_L _21687_ (.A(_13428_),
    .B(_13431_),
    .Y(_13432_));
 NOR3x1_ASAP7_75t_SL _21688_ (.A(_13425_),
    .B(_12911_),
    .C(_13432_),
    .Y(_13433_));
 NOR2x1_ASAP7_75t_R _21689_ (.A(_01142_),
    .B(_12864_),
    .Y(_13434_));
 NOR2x1_ASAP7_75t_R _21690_ (.A(_13434_),
    .B(_13002_),
    .Y(_13435_));
 AOI21x1_ASAP7_75t_R _21691_ (.A1(_13365_),
    .A2(_13435_),
    .B(_12879_),
    .Y(_13436_));
 AO21x1_ASAP7_75t_R _21692_ (.A1(_12980_),
    .A2(_12828_),
    .B(_12838_),
    .Y(_13437_));
 AOI21x1_ASAP7_75t_SL _21693_ (.A1(_13029_),
    .A2(_13038_),
    .B(_12855_),
    .Y(_13438_));
 NAND2x1_ASAP7_75t_R _21694_ (.A(_13437_),
    .B(_13438_),
    .Y(_13439_));
 NAND2x1_ASAP7_75t_SL _21695_ (.A(_13436_),
    .B(_13439_),
    .Y(_13440_));
 INVx1_ASAP7_75t_R _21696_ (.A(_13098_),
    .Y(_13441_));
 OAI21x1_ASAP7_75t_R _21697_ (.A1(_12785_),
    .A2(_12838_),
    .B(_12938_),
    .Y(_13442_));
 AO21x1_ASAP7_75t_R _21698_ (.A1(_12864_),
    .A2(_12970_),
    .B(_13442_),
    .Y(_13443_));
 NAND2x1_ASAP7_75t_R _21699_ (.A(_01133_),
    .B(_12838_),
    .Y(_13444_));
 AOI21x1_ASAP7_75t_R _21700_ (.A1(_12864_),
    .A2(_13380_),
    .B(_12938_),
    .Y(_13445_));
 AOI21x1_ASAP7_75t_R _21701_ (.A1(_13444_),
    .A2(_13445_),
    .B(_12878_),
    .Y(_13446_));
 OAI21x1_ASAP7_75t_SL _21702_ (.A1(_13441_),
    .A2(_13443_),
    .B(_13446_),
    .Y(_13447_));
 NAND3x1_ASAP7_75t_R _21703_ (.A(_13440_),
    .B(_12911_),
    .C(_13447_),
    .Y(_13448_));
 AOI21x1_ASAP7_75t_R _21704_ (.A1(_12838_),
    .A2(_12866_),
    .B(_12948_),
    .Y(_13449_));
 AOI21x1_ASAP7_75t_R _21705_ (.A1(_13445_),
    .A2(_13449_),
    .B(_12879_),
    .Y(_13450_));
 AO21x1_ASAP7_75t_R _21706_ (.A1(_12864_),
    .A2(_12899_),
    .B(_12855_),
    .Y(_13451_));
 AO21x1_ASAP7_75t_SL _21707_ (.A1(_12926_),
    .A2(_13119_),
    .B(_13451_),
    .Y(_13452_));
 AOI21x1_ASAP7_75t_R _21708_ (.A1(_13450_),
    .A2(_13452_),
    .B(_12911_),
    .Y(_13453_));
 NOR2x1_ASAP7_75t_R _21709_ (.A(_13028_),
    .B(_12864_),
    .Y(_13454_));
 AOI21x1_ASAP7_75t_R _21710_ (.A1(_13205_),
    .A2(_13454_),
    .B(_12938_),
    .Y(_13455_));
 OAI21x1_ASAP7_75t_R _21711_ (.A1(_12948_),
    .A2(_13081_),
    .B(_12864_),
    .Y(_13456_));
 NAND2x1_ASAP7_75t_SL _21712_ (.A(_13455_),
    .B(_13456_),
    .Y(_13457_));
 AOI21x1_ASAP7_75t_R _21713_ (.A1(_12821_),
    .A2(_13407_),
    .B(_13442_),
    .Y(_13458_));
 AOI21x1_ASAP7_75t_R _21714_ (.A1(_13183_),
    .A2(_13458_),
    .B(_12878_),
    .Y(_13459_));
 NAND2x1_ASAP7_75t_R _21715_ (.A(_13457_),
    .B(_13459_),
    .Y(_13460_));
 AOI21x1_ASAP7_75t_R _21716_ (.A1(_13453_),
    .A2(_13460_),
    .B(_12920_),
    .Y(_13461_));
 NAND2x1_ASAP7_75t_SL _21717_ (.A(_13448_),
    .B(_13461_),
    .Y(_13462_));
 OAI21x1_ASAP7_75t_SL _21718_ (.A1(_13420_),
    .A2(_13433_),
    .B(_13462_),
    .Y(_00063_));
 XOR2x2_ASAP7_75t_SL _21719_ (.A(_00646_),
    .B(_00639_),
    .Y(_13463_));
 XOR2x1_ASAP7_75t_SL _21720_ (.A(_00640_),
    .Y(_13464_),
    .B(_00672_));
 XOR2x2_ASAP7_75t_SL _21721_ (.A(_13464_),
    .B(_13463_),
    .Y(_13465_));
 XOR2x2_ASAP7_75t_SL _21722_ (.A(_00576_),
    .B(_10669_),
    .Y(_13466_));
 AND2x2_ASAP7_75t_SL _21723_ (.A(_13466_),
    .B(_13465_),
    .Y(_13467_));
 OAI21x1_ASAP7_75t_SL _21724_ (.A1(_13465_),
    .A2(_13466_),
    .B(_00574_),
    .Y(_13468_));
 NAND2x1_ASAP7_75t_R _21725_ (.A(_00456_),
    .B(_10675_),
    .Y(_13469_));
 OAI21x1_ASAP7_75t_SL _21726_ (.A1(_13468_),
    .A2(_13467_),
    .B(_13469_),
    .Y(_13470_));
 XOR2x2_ASAP7_75t_SL _21727_ (.A(_13470_),
    .B(_00846_),
    .Y(_13471_));
 NOR2x1_ASAP7_75t_L _21729_ (.A(_00574_),
    .B(_00457_),
    .Y(_13472_));
 XOR2x2_ASAP7_75t_SL _21730_ (.A(_00614_),
    .B(_00575_),
    .Y(_13473_));
 INVx2_ASAP7_75t_L _21731_ (.A(_13473_),
    .Y(_13474_));
 NAND2x1p5_ASAP7_75t_SL _21732_ (.A(_13474_),
    .B(_00671_),
    .Y(_13475_));
 NAND2x1_ASAP7_75t_L _21733_ (.A(_10691_),
    .B(_13473_),
    .Y(_13476_));
 INVx2_ASAP7_75t_R _21734_ (.A(_13463_),
    .Y(_13477_));
 NAND3x1_ASAP7_75t_R _21735_ (.A(_13475_),
    .B(_13476_),
    .C(_13477_),
    .Y(_13478_));
 AOI21x1_ASAP7_75t_SL _21736_ (.A1(_13476_),
    .A2(_13475_),
    .B(_13477_),
    .Y(_13479_));
 INVx2_ASAP7_75t_SL _21737_ (.A(_13479_),
    .Y(_13480_));
 AOI21x1_ASAP7_75t_SL _21738_ (.A1(_13480_),
    .A2(_13478_),
    .B(_10675_),
    .Y(_13481_));
 OAI21x1_ASAP7_75t_R _21739_ (.A1(_13472_),
    .A2(_13481_),
    .B(_00845_),
    .Y(_13482_));
 XOR2x2_ASAP7_75t_SL _21740_ (.A(_13473_),
    .B(_00671_),
    .Y(_13483_));
 NOR2x1_ASAP7_75t_L _21741_ (.A(_13463_),
    .B(_13483_),
    .Y(_13484_));
 OAI21x1_ASAP7_75t_SL _21742_ (.A1(_13484_),
    .A2(_13479_),
    .B(_00574_),
    .Y(_13485_));
 INVx1_ASAP7_75t_R _21743_ (.A(_00845_),
    .Y(_13486_));
 INVx1_ASAP7_75t_R _21744_ (.A(_13472_),
    .Y(_13487_));
 NAND3x1_ASAP7_75t_R _21745_ (.A(_13485_),
    .B(_13486_),
    .C(_13487_),
    .Y(_13488_));
 NAND2x1_ASAP7_75t_SL _21746_ (.A(_13482_),
    .B(_13488_),
    .Y(_13489_));
 NOR2x1_ASAP7_75t_SL _21748_ (.A(_00574_),
    .B(_00458_),
    .Y(_13490_));
 INVx1_ASAP7_75t_SL _21749_ (.A(_13490_),
    .Y(_13491_));
 INVx1_ASAP7_75t_SL _21750_ (.A(_00577_),
    .Y(_13492_));
 NOR2x1_ASAP7_75t_SL _21751_ (.A(_13492_),
    .B(_10714_),
    .Y(_13493_));
 NOR2x1_ASAP7_75t_SL _21752_ (.A(_00577_),
    .B(_10710_),
    .Y(_13494_));
 OAI21x1_ASAP7_75t_SL _21753_ (.A1(_13493_),
    .A2(_13494_),
    .B(_10667_),
    .Y(_13495_));
 INVx1_ASAP7_75t_SL _21754_ (.A(_13495_),
    .Y(_13496_));
 NOR3x1_ASAP7_75t_SL _21755_ (.A(_13494_),
    .B(_13493_),
    .C(_10667_),
    .Y(_13497_));
 OAI21x1_ASAP7_75t_SL _21756_ (.A1(_13496_),
    .A2(_13497_),
    .B(_00574_),
    .Y(_13498_));
 INVx1_ASAP7_75t_SL _21757_ (.A(_00847_),
    .Y(_13499_));
 AOI21x1_ASAP7_75t_SL _21758_ (.A1(_13491_),
    .A2(_13498_),
    .B(_13499_),
    .Y(_13500_));
 NAND2x1_ASAP7_75t_SL _21759_ (.A(_00458_),
    .B(_10675_),
    .Y(_13501_));
 INVx1_ASAP7_75t_SL _21760_ (.A(_10667_),
    .Y(_13502_));
 XOR2x2_ASAP7_75t_SL _21761_ (.A(_10714_),
    .B(_13492_),
    .Y(_13503_));
 NAND2x1_ASAP7_75t_SL _21762_ (.A(_13502_),
    .B(_13503_),
    .Y(_13504_));
 NAND3x1_ASAP7_75t_SL _21763_ (.A(_13504_),
    .B(_00574_),
    .C(_13495_),
    .Y(_13505_));
 AOI21x1_ASAP7_75t_SL _21764_ (.A1(_13501_),
    .A2(_13505_),
    .B(_00847_),
    .Y(_13506_));
 NOR2x2_ASAP7_75t_SL _21765_ (.A(_13500_),
    .B(_13506_),
    .Y(_13507_));
 OAI21x1_ASAP7_75t_SL _21767_ (.A1(_13481_),
    .A2(_13472_),
    .B(_13486_),
    .Y(_13508_));
 NAND3x1_ASAP7_75t_SL _21768_ (.A(_13485_),
    .B(_00845_),
    .C(_13487_),
    .Y(_13509_));
 NAND2x2_ASAP7_75t_SL _21769_ (.A(_13509_),
    .B(_13508_),
    .Y(_13510_));
 AOI21x1_ASAP7_75t_SL _21771_ (.A1(_13491_),
    .A2(_13498_),
    .B(_00847_),
    .Y(_13511_));
 AOI21x1_ASAP7_75t_SL _21772_ (.A1(_13501_),
    .A2(_13505_),
    .B(_13499_),
    .Y(_13512_));
 NOR2x2_ASAP7_75t_SL _21773_ (.A(_13511_),
    .B(_13512_),
    .Y(_13513_));
 NAND2x2_ASAP7_75t_SL _21777_ (.A(_01155_),
    .B(_13513_),
    .Y(_13516_));
 NOR2x1_ASAP7_75t_R _21779_ (.A(_00574_),
    .B(_00559_),
    .Y(_13518_));
 XOR2x2_ASAP7_75t_L _21780_ (.A(_00641_),
    .B(_00646_),
    .Y(_13519_));
 XOR2x2_ASAP7_75t_SL _21781_ (.A(_10763_),
    .B(_13519_),
    .Y(_13520_));
 XNOR2x2_ASAP7_75t_L _21782_ (.A(_00578_),
    .B(_10764_),
    .Y(_13521_));
 XOR2x2_ASAP7_75t_SL _21783_ (.A(_13520_),
    .B(_13521_),
    .Y(_13522_));
 NOR2x1_ASAP7_75t_SL _21784_ (.A(_10675_),
    .B(_13522_),
    .Y(_13523_));
 INVx1_ASAP7_75t_R _21785_ (.A(_00848_),
    .Y(_13524_));
 OAI21x1_ASAP7_75t_R _21786_ (.A1(_13518_),
    .A2(_13523_),
    .B(_13524_),
    .Y(_13525_));
 NOR2x1_ASAP7_75t_L _21787_ (.A(_13521_),
    .B(_13520_),
    .Y(_13526_));
 AND2x2_ASAP7_75t_SL _21788_ (.A(_13520_),
    .B(_13521_),
    .Y(_13527_));
 OAI21x1_ASAP7_75t_SL _21789_ (.A1(_13526_),
    .A2(_13527_),
    .B(_00574_),
    .Y(_13528_));
 INVx1_ASAP7_75t_R _21790_ (.A(_13518_),
    .Y(_13529_));
 NAND3x1_ASAP7_75t_SL _21791_ (.A(_13528_),
    .B(_00848_),
    .C(_13529_),
    .Y(_13530_));
 NAND2x1_ASAP7_75t_SL _21792_ (.A(_13525_),
    .B(_13530_),
    .Y(_13531_));
 NOR2x1_ASAP7_75t_L _21794_ (.A(_13489_),
    .B(_13513_),
    .Y(_13533_));
 NOR2x1_ASAP7_75t_SL _21795_ (.A(_13531_),
    .B(_13533_),
    .Y(_13534_));
 NAND2x1_ASAP7_75t_SL _21796_ (.A(_13516_),
    .B(_13534_),
    .Y(_13535_));
 XNOR2x2_ASAP7_75t_SL _21798_ (.A(_13470_),
    .B(_00846_),
    .Y(_13537_));
 NOR2x2_ASAP7_75t_SL _21800_ (.A(_13537_),
    .B(_13489_),
    .Y(_13538_));
 NAND2x1_ASAP7_75t_R _21801_ (.A(_13507_),
    .B(_13538_),
    .Y(_13539_));
 OAI21x1_ASAP7_75t_SL _21802_ (.A1(_13518_),
    .A2(_13523_),
    .B(_00848_),
    .Y(_13540_));
 NAND3x1_ASAP7_75t_SL _21803_ (.A(_13528_),
    .B(_13524_),
    .C(_13529_),
    .Y(_13541_));
 NAND2x1_ASAP7_75t_SL _21804_ (.A(_13540_),
    .B(_13541_),
    .Y(_13542_));
 NOR2x1_ASAP7_75t_SL _21806_ (.A(_13471_),
    .B(_13507_),
    .Y(_13544_));
 NOR2x1_ASAP7_75t_SL _21807_ (.A(_13542_),
    .B(_13544_),
    .Y(_13545_));
 AND2x2_ASAP7_75t_R _21808_ (.A(_10675_),
    .B(_00558_),
    .Y(_13546_));
 XOR2x2_ASAP7_75t_R _21809_ (.A(_00579_),
    .B(_00643_),
    .Y(_13547_));
 XOR2x2_ASAP7_75t_SL _21810_ (.A(_10746_),
    .B(_13547_),
    .Y(_13548_));
 XOR2x2_ASAP7_75t_L _21811_ (.A(_00642_),
    .B(_00646_),
    .Y(_13549_));
 INVx1_ASAP7_75t_R _21812_ (.A(_00675_),
    .Y(_13550_));
 XOR2x2_ASAP7_75t_SL _21813_ (.A(_13549_),
    .B(_13550_),
    .Y(_13551_));
 XOR2x2_ASAP7_75t_SL _21814_ (.A(_13548_),
    .B(_13551_),
    .Y(_13552_));
 NOR2x1_ASAP7_75t_R _21815_ (.A(_10675_),
    .B(_13552_),
    .Y(_13553_));
 OAI21x1_ASAP7_75t_R _21816_ (.A1(_13546_),
    .A2(_13553_),
    .B(_00850_),
    .Y(_13554_));
 NOR2x1_ASAP7_75t_R _21817_ (.A(_00574_),
    .B(_00558_),
    .Y(_13555_));
 XNOR2x2_ASAP7_75t_SL _21818_ (.A(_13551_),
    .B(_13548_),
    .Y(_13556_));
 NOR2x1_ASAP7_75t_R _21819_ (.A(_10675_),
    .B(_13556_),
    .Y(_13557_));
 INVx1_ASAP7_75t_R _21820_ (.A(_00850_),
    .Y(_13558_));
 OAI21x1_ASAP7_75t_R _21821_ (.A1(_13555_),
    .A2(_13557_),
    .B(_13558_),
    .Y(_13559_));
 NAND2x2_ASAP7_75t_SL _21822_ (.A(_13554_),
    .B(_13559_),
    .Y(_13560_));
 AOI21x1_ASAP7_75t_SL _21824_ (.A1(_13539_),
    .A2(_13545_),
    .B(_13560_),
    .Y(_13562_));
 NAND2x1_ASAP7_75t_SL _21825_ (.A(_13535_),
    .B(_13562_),
    .Y(_13563_));
 INVx1_ASAP7_75t_SL _21826_ (.A(_01148_),
    .Y(_13564_));
 OAI21x1_ASAP7_75t_R _21827_ (.A1(_13500_),
    .A2(_13506_),
    .B(_13564_),
    .Y(_13565_));
 OAI21x1_ASAP7_75t_SL _21828_ (.A1(_13565_),
    .A2(_13542_),
    .B(_13560_),
    .Y(_13566_));
 NAND2x1_ASAP7_75t_SL _21829_ (.A(_13537_),
    .B(_13507_),
    .Y(_13567_));
 NOR2x1_ASAP7_75t_SL _21830_ (.A(_13542_),
    .B(_13567_),
    .Y(_13568_));
 NOR2x1_ASAP7_75t_SL _21831_ (.A(_13566_),
    .B(_13568_),
    .Y(_13569_));
 NOR2x2_ASAP7_75t_SL _21832_ (.A(_13537_),
    .B(_13510_),
    .Y(_13570_));
 NAND2x2_ASAP7_75t_SL _21833_ (.A(_13513_),
    .B(_13570_),
    .Y(_13571_));
 NAND2x1_ASAP7_75t_SL _21834_ (.A(_13571_),
    .B(_13534_),
    .Y(_13572_));
 XOR2x2_ASAP7_75t_R _21835_ (.A(_00643_),
    .B(_00644_),
    .Y(_13573_));
 INVx1_ASAP7_75t_R _21836_ (.A(_00676_),
    .Y(_13574_));
 XOR2x2_ASAP7_75t_SL _21837_ (.A(_13573_),
    .B(_13574_),
    .Y(_13575_));
 XNOR2x2_ASAP7_75t_R _21838_ (.A(_00580_),
    .B(_00611_),
    .Y(_13576_));
 XOR2x2_ASAP7_75t_SL _21839_ (.A(_13575_),
    .B(_13576_),
    .Y(_13577_));
 NOR2x1_ASAP7_75t_R _21841_ (.A(_00574_),
    .B(_00557_),
    .Y(_13579_));
 INVx1_ASAP7_75t_R _21842_ (.A(_13579_),
    .Y(_13580_));
 OA21x2_ASAP7_75t_R _21843_ (.A1(_13577_),
    .A2(_10675_),
    .B(_13580_),
    .Y(_13581_));
 XOR2x2_ASAP7_75t_SL _21844_ (.A(_13581_),
    .B(_00851_),
    .Y(_13582_));
 AOI21x1_ASAP7_75t_SL _21845_ (.A1(_13569_),
    .A2(_13572_),
    .B(_13582_),
    .Y(_13583_));
 NAND2x1_ASAP7_75t_SL _21846_ (.A(_13563_),
    .B(_13583_),
    .Y(_13584_));
 NAND2x2_ASAP7_75t_L _21847_ (.A(_01147_),
    .B(_13513_),
    .Y(_13585_));
 AOI21x1_ASAP7_75t_R _21848_ (.A1(_13495_),
    .A2(_13504_),
    .B(_10675_),
    .Y(_13586_));
 OAI21x1_ASAP7_75t_R _21849_ (.A1(_13490_),
    .A2(_13586_),
    .B(_13499_),
    .Y(_13587_));
 NAND3x1_ASAP7_75t_R _21850_ (.A(_13498_),
    .B(_00847_),
    .C(_13491_),
    .Y(_13588_));
 INVx2_ASAP7_75t_R _21851_ (.A(_01155_),
    .Y(_13589_));
 AOI21x1_ASAP7_75t_SL _21852_ (.A1(_13587_),
    .A2(_13588_),
    .B(_13589_),
    .Y(_13590_));
 NOR2x1_ASAP7_75t_SL _21853_ (.A(_13531_),
    .B(_13590_),
    .Y(_13591_));
 NAND2x1_ASAP7_75t_SL _21854_ (.A(_13585_),
    .B(_13591_),
    .Y(_13592_));
 AO21x1_ASAP7_75t_R _21856_ (.A1(_13507_),
    .A2(_13537_),
    .B(_13489_),
    .Y(_13594_));
 AOI21x1_ASAP7_75t_SL _21857_ (.A1(_13531_),
    .A2(_13594_),
    .B(_13560_),
    .Y(_13595_));
 NAND2x1_ASAP7_75t_SL _21858_ (.A(_13592_),
    .B(_13595_),
    .Y(_13596_));
 INVx2_ASAP7_75t_SL _21859_ (.A(_13560_),
    .Y(_13597_));
 AOI21x1_ASAP7_75t_R _21861_ (.A1(_13510_),
    .A2(_13507_),
    .B(_13542_),
    .Y(_13599_));
 NOR2x1_ASAP7_75t_SL _21862_ (.A(_13597_),
    .B(_13599_),
    .Y(_13600_));
 AOI21x1_ASAP7_75t_SL _21865_ (.A1(_01150_),
    .A2(_13513_),
    .B(_13531_),
    .Y(_13603_));
 NAND2x1_ASAP7_75t_SL _21866_ (.A(_13603_),
    .B(_13539_),
    .Y(_13604_));
 XNOR2x2_ASAP7_75t_SL _21867_ (.A(_00851_),
    .B(_13581_),
    .Y(_13605_));
 AOI21x1_ASAP7_75t_SL _21869_ (.A1(_13600_),
    .A2(_13604_),
    .B(_13605_),
    .Y(_13607_));
 XOR2x2_ASAP7_75t_SL _21870_ (.A(_00645_),
    .B(_00677_),
    .Y(_13608_));
 XOR2x2_ASAP7_75t_R _21871_ (.A(_10826_),
    .B(_00581_),
    .Y(_13609_));
 XNOR2x2_ASAP7_75t_R _21872_ (.A(_13608_),
    .B(_13609_),
    .Y(_13610_));
 NOR2x1_ASAP7_75t_R _21873_ (.A(_00574_),
    .B(_00556_),
    .Y(_13611_));
 AO21x1_ASAP7_75t_SL _21874_ (.A1(_13610_),
    .A2(_00574_),
    .B(_13611_),
    .Y(_13612_));
 XOR2x2_ASAP7_75t_SL _21875_ (.A(_13612_),
    .B(_00852_),
    .Y(_13613_));
 AOI21x1_ASAP7_75t_SL _21877_ (.A1(_13596_),
    .A2(_13607_),
    .B(_13613_),
    .Y(_13615_));
 XNOR2x2_ASAP7_75t_R _21878_ (.A(_00582_),
    .B(_00613_),
    .Y(_13616_));
 XOR2x2_ASAP7_75t_R _21879_ (.A(_00645_),
    .B(_00646_),
    .Y(_13617_));
 XOR2x2_ASAP7_75t_R _21880_ (.A(_13617_),
    .B(_10879_),
    .Y(_13618_));
 XNOR2x2_ASAP7_75t_R _21881_ (.A(_13616_),
    .B(_13618_),
    .Y(_13619_));
 NOR2x1_ASAP7_75t_R _21882_ (.A(_00574_),
    .B(_00555_),
    .Y(_13620_));
 AO21x1_ASAP7_75t_SL _21883_ (.A1(_13619_),
    .A2(_00574_),
    .B(_13620_),
    .Y(_13621_));
 XOR2x2_ASAP7_75t_SL _21884_ (.A(_13621_),
    .B(_00853_),
    .Y(_13622_));
 INVx2_ASAP7_75t_SL _21885_ (.A(_13622_),
    .Y(_13623_));
 AOI21x1_ASAP7_75t_SL _21886_ (.A1(_13584_),
    .A2(_13615_),
    .B(_13623_),
    .Y(_13624_));
 NOR2x1_ASAP7_75t_SL _21887_ (.A(_13510_),
    .B(_13513_),
    .Y(_13625_));
 OAI21x1_ASAP7_75t_SL _21889_ (.A1(_13538_),
    .A2(_13625_),
    .B(_13531_),
    .Y(_13627_));
 NAND2x1_ASAP7_75t_R _21890_ (.A(_13489_),
    .B(_13507_),
    .Y(_13628_));
 AOI21x1_ASAP7_75t_R _21891_ (.A1(_13471_),
    .A2(_13510_),
    .B(_13531_),
    .Y(_13629_));
 AOI21x1_ASAP7_75t_SL _21892_ (.A1(_13628_),
    .A2(_13629_),
    .B(_13560_),
    .Y(_13630_));
 NAND2x1_ASAP7_75t_SL _21893_ (.A(_13627_),
    .B(_13630_),
    .Y(_13631_));
 NAND2x1_ASAP7_75t_R _21894_ (.A(_13507_),
    .B(_13570_),
    .Y(_13632_));
 INVx2_ASAP7_75t_SL _21895_ (.A(_01147_),
    .Y(_13633_));
 NOR2x1_ASAP7_75t_SL _21896_ (.A(_13633_),
    .B(_13507_),
    .Y(_13634_));
 NOR2x1_ASAP7_75t_SL _21897_ (.A(_13542_),
    .B(_13634_),
    .Y(_13635_));
 NAND2x1_ASAP7_75t_SL _21898_ (.A(_13632_),
    .B(_13635_),
    .Y(_13636_));
 INVx1_ASAP7_75t_SL _21900_ (.A(_01152_),
    .Y(_13638_));
 OAI21x1_ASAP7_75t_SL _21901_ (.A1(_13511_),
    .A2(_13512_),
    .B(_01146_),
    .Y(_13639_));
 OAI21x1_ASAP7_75t_R _21902_ (.A1(_13638_),
    .A2(_13507_),
    .B(_13639_),
    .Y(_13640_));
 AOI21x1_ASAP7_75t_SL _21903_ (.A1(_13542_),
    .A2(_13640_),
    .B(_13597_),
    .Y(_13641_));
 AOI21x1_ASAP7_75t_SL _21904_ (.A1(_13636_),
    .A2(_13641_),
    .B(_13605_),
    .Y(_13642_));
 NAND2x1_ASAP7_75t_SL _21905_ (.A(_13631_),
    .B(_13642_),
    .Y(_13643_));
 NOR2x2_ASAP7_75t_L _21906_ (.A(_13537_),
    .B(_13513_),
    .Y(_13644_));
 OAI21x1_ASAP7_75t_SL _21907_ (.A1(_13500_),
    .A2(_13506_),
    .B(_13633_),
    .Y(_13645_));
 NAND2x1p5_ASAP7_75t_SL _21908_ (.A(_13531_),
    .B(_13645_),
    .Y(_13646_));
 NOR2x1_ASAP7_75t_SL _21909_ (.A(_13644_),
    .B(_13646_),
    .Y(_13647_));
 NAND2x1_ASAP7_75t_SL _21912_ (.A(_01147_),
    .B(_13507_),
    .Y(_13650_));
 AOI21x1_ASAP7_75t_SL _21913_ (.A1(_13542_),
    .A2(_13650_),
    .B(_13560_),
    .Y(_13651_));
 INVx1_ASAP7_75t_SL _21914_ (.A(_13651_),
    .Y(_13652_));
 NOR2x1_ASAP7_75t_SL _21915_ (.A(_13647_),
    .B(_13652_),
    .Y(_13653_));
 AO21x1_ASAP7_75t_SL _21917_ (.A1(_13639_),
    .A2(_13645_),
    .B(_13531_),
    .Y(_13655_));
 OAI21x1_ASAP7_75t_SL _21918_ (.A1(_13500_),
    .A2(_13506_),
    .B(_01146_),
    .Y(_13656_));
 INVx1_ASAP7_75t_SL _21919_ (.A(_13656_),
    .Y(_13657_));
 NOR2x1_ASAP7_75t_SL _21920_ (.A(_13638_),
    .B(_13513_),
    .Y(_13658_));
 OAI21x1_ASAP7_75t_SL _21922_ (.A1(_13657_),
    .A2(_13658_),
    .B(_13531_),
    .Y(_13660_));
 AOI21x1_ASAP7_75t_SL _21924_ (.A1(_13655_),
    .A2(_13660_),
    .B(_13597_),
    .Y(_13662_));
 OAI21x1_ASAP7_75t_SL _21925_ (.A1(_13653_),
    .A2(_13662_),
    .B(_13605_),
    .Y(_13663_));
 NAND3x1_ASAP7_75t_SL _21927_ (.A(_13643_),
    .B(_13663_),
    .C(_13613_),
    .Y(_13665_));
 NAND2x1_ASAP7_75t_SL _21928_ (.A(_13624_),
    .B(_13665_),
    .Y(_13666_));
 AND2x2_ASAP7_75t_R _21932_ (.A(_01148_),
    .B(_01150_),
    .Y(_13670_));
 NOR2x1_ASAP7_75t_SL _21933_ (.A(_13670_),
    .B(_13513_),
    .Y(_13671_));
 AOI21x1_ASAP7_75t_R _21934_ (.A1(_13471_),
    .A2(_13510_),
    .B(_13507_),
    .Y(_13672_));
 NOR2x1_ASAP7_75t_SL _21935_ (.A(_13671_),
    .B(_13672_),
    .Y(_13673_));
 OAI21x1_ASAP7_75t_SL _21937_ (.A1(_13657_),
    .A2(_13625_),
    .B(_13542_),
    .Y(_13675_));
 OAI21x1_ASAP7_75t_SL _21938_ (.A1(_13542_),
    .A2(_13673_),
    .B(_13675_),
    .Y(_13676_));
 AO21x1_ASAP7_75t_SL _21939_ (.A1(_13541_),
    .A2(_13540_),
    .B(_01160_),
    .Y(_13677_));
 OAI21x1_ASAP7_75t_SL _21940_ (.A1(_13511_),
    .A2(_13512_),
    .B(_13633_),
    .Y(_13678_));
 OA21x2_ASAP7_75t_SL _21941_ (.A1(_13542_),
    .A2(_13678_),
    .B(_13597_),
    .Y(_13679_));
 AOI21x1_ASAP7_75t_SL _21943_ (.A1(_13677_),
    .A2(_13679_),
    .B(_13582_),
    .Y(_13681_));
 OAI21x1_ASAP7_75t_SL _21944_ (.A1(_13597_),
    .A2(_13676_),
    .B(_13681_),
    .Y(_13682_));
 NAND2x2_ASAP7_75t_SL _21945_ (.A(_13513_),
    .B(_13538_),
    .Y(_13683_));
 AOI21x1_ASAP7_75t_SL _21946_ (.A1(_13638_),
    .A2(_13507_),
    .B(_13542_),
    .Y(_13684_));
 OAI21x1_ASAP7_75t_SL _21947_ (.A1(_13531_),
    .A2(_13565_),
    .B(_13597_),
    .Y(_13685_));
 AO21x1_ASAP7_75t_SL _21948_ (.A1(_13683_),
    .A2(_13684_),
    .B(_13685_),
    .Y(_13686_));
 INVx1_ASAP7_75t_SL _21949_ (.A(_13566_),
    .Y(_13687_));
 INVx1_ASAP7_75t_R _21950_ (.A(_01153_),
    .Y(_13688_));
 AOI21x1_ASAP7_75t_SL _21951_ (.A1(_13587_),
    .A2(_13588_),
    .B(_13688_),
    .Y(_13689_));
 NOR2x1p5_ASAP7_75t_SL _21952_ (.A(_13531_),
    .B(_13689_),
    .Y(_13690_));
 NAND2x1_ASAP7_75t_SL _21953_ (.A(_13690_),
    .B(_13683_),
    .Y(_13691_));
 AOI21x1_ASAP7_75t_SL _21954_ (.A1(_13687_),
    .A2(_13691_),
    .B(_13605_),
    .Y(_13692_));
 NAND2x1_ASAP7_75t_SL _21955_ (.A(_13686_),
    .B(_13692_),
    .Y(_13693_));
 INVx1_ASAP7_75t_SL _21956_ (.A(_13613_),
    .Y(_13694_));
 AOI21x1_ASAP7_75t_SL _21958_ (.A1(_13682_),
    .A2(_13693_),
    .B(_13694_),
    .Y(_13696_));
 INVx1_ASAP7_75t_SL _21959_ (.A(_13603_),
    .Y(_13697_));
 AO21x1_ASAP7_75t_SL _21961_ (.A1(_13565_),
    .A2(_13639_),
    .B(_13542_),
    .Y(_13699_));
 AOI21x1_ASAP7_75t_SL _21963_ (.A1(_13697_),
    .A2(_13699_),
    .B(_13560_),
    .Y(_13701_));
 NOR2x2_ASAP7_75t_SL _21964_ (.A(_13513_),
    .B(_13633_),
    .Y(_13702_));
 OAI21x1_ASAP7_75t_SL _21965_ (.A1(_13544_),
    .A2(_13702_),
    .B(_13531_),
    .Y(_13703_));
 NOR2x1_ASAP7_75t_SL _21966_ (.A(_13510_),
    .B(_13507_),
    .Y(_13704_));
 OAI21x1_ASAP7_75t_SL _21967_ (.A1(_13658_),
    .A2(_13704_),
    .B(_13542_),
    .Y(_13705_));
 AOI21x1_ASAP7_75t_SL _21969_ (.A1(_13703_),
    .A2(_13705_),
    .B(_13597_),
    .Y(_13707_));
 OAI21x1_ASAP7_75t_SL _21971_ (.A1(_13701_),
    .A2(_13707_),
    .B(_13582_),
    .Y(_13709_));
 INVx2_ASAP7_75t_SL _21972_ (.A(_01150_),
    .Y(_13710_));
 OAI21x1_ASAP7_75t_SL _21973_ (.A1(_13511_),
    .A2(_13512_),
    .B(_13710_),
    .Y(_13711_));
 OA21x2_ASAP7_75t_R _21974_ (.A1(_13711_),
    .A2(_13542_),
    .B(_13597_),
    .Y(_13712_));
 NAND2x2_ASAP7_75t_SL _21975_ (.A(_13688_),
    .B(_13513_),
    .Y(_13713_));
 NOR2x1_ASAP7_75t_SL _21976_ (.A(_13542_),
    .B(_13713_),
    .Y(_13714_));
 NOR2x1p5_ASAP7_75t_SL _21977_ (.A(_13531_),
    .B(_13634_),
    .Y(_13715_));
 NOR2x1_ASAP7_75t_SL _21978_ (.A(_13714_),
    .B(_13715_),
    .Y(_13716_));
 NAND2x1_ASAP7_75t_SL _21979_ (.A(_13712_),
    .B(_13716_),
    .Y(_13717_));
 OAI21x1_ASAP7_75t_SL _21980_ (.A1(_13711_),
    .A2(_13542_),
    .B(_13560_),
    .Y(_13718_));
 AOI21x1_ASAP7_75t_SL _21981_ (.A1(_13571_),
    .A2(_13534_),
    .B(_13718_),
    .Y(_13719_));
 NOR2x1_ASAP7_75t_SL _21982_ (.A(_13582_),
    .B(_13719_),
    .Y(_13720_));
 NAND2x1_ASAP7_75t_SL _21983_ (.A(_13717_),
    .B(_13720_),
    .Y(_13721_));
 AOI21x1_ASAP7_75t_SL _21984_ (.A1(_13709_),
    .A2(_13721_),
    .B(_13613_),
    .Y(_13722_));
 OAI21x1_ASAP7_75t_SL _21985_ (.A1(_13696_),
    .A2(_13722_),
    .B(_13623_),
    .Y(_13723_));
 NAND2x1_ASAP7_75t_SL _21986_ (.A(_13666_),
    .B(_13723_),
    .Y(_00064_));
 AND3x1_ASAP7_75t_SL _21987_ (.A(_13530_),
    .B(_01162_),
    .C(_13525_),
    .Y(_13724_));
 AOI21x1_ASAP7_75t_SL _21989_ (.A1(_13605_),
    .A2(_13724_),
    .B(_13597_),
    .Y(_13726_));
 NAND2x1_ASAP7_75t_SL _21990_ (.A(_13684_),
    .B(_13571_),
    .Y(_13727_));
 AO21x1_ASAP7_75t_SL _21991_ (.A1(_13726_),
    .A2(_13727_),
    .B(_13694_),
    .Y(_13728_));
 NAND2x2_ASAP7_75t_SL _21992_ (.A(_13489_),
    .B(_13513_),
    .Y(_13729_));
 NAND2x1_ASAP7_75t_SL _21993_ (.A(_13531_),
    .B(_13729_),
    .Y(_13730_));
 OAI21x1_ASAP7_75t_SL _21994_ (.A1(_13644_),
    .A2(_13730_),
    .B(_13605_),
    .Y(_13731_));
 NOR2x1_ASAP7_75t_SL _21995_ (.A(_01150_),
    .B(_13507_),
    .Y(_13732_));
 OAI21x1_ASAP7_75t_SL _21997_ (.A1(_13644_),
    .A2(_13732_),
    .B(_13542_),
    .Y(_13734_));
 NAND2x1_ASAP7_75t_SL _21998_ (.A(_13597_),
    .B(_13734_),
    .Y(_13735_));
 NOR2x1_ASAP7_75t_SL _21999_ (.A(_13731_),
    .B(_13735_),
    .Y(_13736_));
 AO21x1_ASAP7_75t_SL _22000_ (.A1(_13510_),
    .A2(_13471_),
    .B(_13513_),
    .Y(_13737_));
 AOI21x1_ASAP7_75t_SL _22001_ (.A1(_13471_),
    .A2(_13489_),
    .B(_13507_),
    .Y(_13738_));
 INVx1_ASAP7_75t_SL _22002_ (.A(_13738_),
    .Y(_13739_));
 AOI21x1_ASAP7_75t_SL _22004_ (.A1(_13737_),
    .A2(_13739_),
    .B(_13531_),
    .Y(_13741_));
 NOR2x1_ASAP7_75t_SL _22005_ (.A(_13489_),
    .B(_13507_),
    .Y(_13742_));
 INVx1_ASAP7_75t_R _22006_ (.A(_01146_),
    .Y(_13743_));
 AO21x1_ASAP7_75t_SL _22007_ (.A1(_13743_),
    .A2(_13507_),
    .B(_13542_),
    .Y(_13744_));
 NOR2x1_ASAP7_75t_SL _22008_ (.A(_13560_),
    .B(_13605_),
    .Y(_13745_));
 OAI21x1_ASAP7_75t_SL _22009_ (.A1(_13742_),
    .A2(_13744_),
    .B(_13745_),
    .Y(_13746_));
 NOR2x1_ASAP7_75t_SL _22010_ (.A(_13741_),
    .B(_13746_),
    .Y(_13747_));
 NOR3x1_ASAP7_75t_SL _22011_ (.A(_13728_),
    .B(_13736_),
    .C(_13747_),
    .Y(_13748_));
 OAI21x1_ASAP7_75t_R _22012_ (.A1(_13511_),
    .A2(_13512_),
    .B(_13564_),
    .Y(_13749_));
 OAI21x1_ASAP7_75t_SL _22013_ (.A1(_01155_),
    .A2(_13507_),
    .B(_13749_),
    .Y(_13750_));
 AOI21x1_ASAP7_75t_SL _22014_ (.A1(_13531_),
    .A2(_13750_),
    .B(_13560_),
    .Y(_13751_));
 OAI21x1_ASAP7_75t_SL _22015_ (.A1(_13537_),
    .A2(_13510_),
    .B(_13507_),
    .Y(_13752_));
 AO21x1_ASAP7_75t_SL _22016_ (.A1(_13752_),
    .A2(_13585_),
    .B(_13531_),
    .Y(_13753_));
 NAND2x1_ASAP7_75t_SL _22017_ (.A(_13751_),
    .B(_13753_),
    .Y(_13754_));
 AOI21x1_ASAP7_75t_SL _22018_ (.A1(_13542_),
    .A2(_13585_),
    .B(_13597_),
    .Y(_13755_));
 NAND2x1_ASAP7_75t_SL _22019_ (.A(_13599_),
    .B(_13571_),
    .Y(_13756_));
 AOI21x1_ASAP7_75t_SL _22020_ (.A1(_13755_),
    .A2(_13756_),
    .B(_13582_),
    .Y(_13757_));
 NAND2x1_ASAP7_75t_SL _22021_ (.A(_13754_),
    .B(_13757_),
    .Y(_13758_));
 AO21x1_ASAP7_75t_SL _22022_ (.A1(_13678_),
    .A2(_13656_),
    .B(_13531_),
    .Y(_13759_));
 INVx1_ASAP7_75t_SL _22023_ (.A(_13565_),
    .Y(_13760_));
 OAI21x1_ASAP7_75t_SL _22024_ (.A1(_13760_),
    .A2(_13625_),
    .B(_13531_),
    .Y(_13761_));
 AOI21x1_ASAP7_75t_SL _22025_ (.A1(_13759_),
    .A2(_13761_),
    .B(_13560_),
    .Y(_13762_));
 INVx1_ASAP7_75t_SL _22026_ (.A(_13639_),
    .Y(_13763_));
 OAI21x1_ASAP7_75t_SL _22027_ (.A1(_13763_),
    .A2(_13742_),
    .B(_13531_),
    .Y(_13764_));
 AOI21x1_ASAP7_75t_SL _22028_ (.A1(_13764_),
    .A2(_13734_),
    .B(_13597_),
    .Y(_13765_));
 OAI21x1_ASAP7_75t_SL _22029_ (.A1(_13762_),
    .A2(_13765_),
    .B(_13582_),
    .Y(_13766_));
 AOI21x1_ASAP7_75t_SL _22030_ (.A1(_13758_),
    .A2(_13766_),
    .B(_13613_),
    .Y(_13767_));
 OAI21x1_ASAP7_75t_SL _22032_ (.A1(_13748_),
    .A2(_13767_),
    .B(_13622_),
    .Y(_13769_));
 NAND2x1_ASAP7_75t_SL _22033_ (.A(_13710_),
    .B(_13513_),
    .Y(_13770_));
 OA21x2_ASAP7_75t_SL _22034_ (.A1(_13770_),
    .A2(_13542_),
    .B(_13560_),
    .Y(_13771_));
 NAND2x1_ASAP7_75t_SL _22035_ (.A(_13771_),
    .B(_13753_),
    .Y(_13772_));
 NAND2x1_ASAP7_75t_SL _22036_ (.A(_13531_),
    .B(_13738_),
    .Y(_13773_));
 NAND2x2_ASAP7_75t_SL _22037_ (.A(_13537_),
    .B(_13513_),
    .Y(_13774_));
 AOI21x1_ASAP7_75t_SL _22039_ (.A1(_13774_),
    .A2(_13591_),
    .B(_13560_),
    .Y(_13776_));
 AOI21x1_ASAP7_75t_SL _22040_ (.A1(_13773_),
    .A2(_13776_),
    .B(_13605_),
    .Y(_13777_));
 NAND2x1_ASAP7_75t_SL _22041_ (.A(_13772_),
    .B(_13777_),
    .Y(_13778_));
 INVx1_ASAP7_75t_SL _22042_ (.A(_13711_),
    .Y(_13779_));
 OAI21x1_ASAP7_75t_SL _22043_ (.A1(_13779_),
    .A2(_13634_),
    .B(_13542_),
    .Y(_13780_));
 OAI21x1_ASAP7_75t_SL _22044_ (.A1(_13657_),
    .A2(_13625_),
    .B(_13531_),
    .Y(_13781_));
 AOI21x1_ASAP7_75t_SL _22045_ (.A1(_13780_),
    .A2(_13781_),
    .B(_13560_),
    .Y(_13782_));
 OAI21x1_ASAP7_75t_SL _22046_ (.A1(_13570_),
    .A2(_13742_),
    .B(_13542_),
    .Y(_13783_));
 OAI21x1_ASAP7_75t_SL _22047_ (.A1(_13702_),
    .A2(_13704_),
    .B(_13531_),
    .Y(_13784_));
 AOI21x1_ASAP7_75t_SL _22048_ (.A1(_13783_),
    .A2(_13784_),
    .B(_13597_),
    .Y(_13785_));
 OAI21x1_ASAP7_75t_SL _22050_ (.A1(_13782_),
    .A2(_13785_),
    .B(_13605_),
    .Y(_13787_));
 AOI21x1_ASAP7_75t_SL _22051_ (.A1(_13778_),
    .A2(_13787_),
    .B(_13613_),
    .Y(_13788_));
 OAI21x1_ASAP7_75t_SL _22052_ (.A1(_13779_),
    .A2(_13672_),
    .B(_13531_),
    .Y(_13789_));
 NOR2x1p5_ASAP7_75t_SL _22053_ (.A(_13531_),
    .B(_13702_),
    .Y(_13790_));
 AOI21x1_ASAP7_75t_SL _22054_ (.A1(_13516_),
    .A2(_13790_),
    .B(_13597_),
    .Y(_13791_));
 NAND2x1_ASAP7_75t_SL _22055_ (.A(_13789_),
    .B(_13791_),
    .Y(_13792_));
 OA21x2_ASAP7_75t_SL _22056_ (.A1(_13644_),
    .A2(_13531_),
    .B(_13774_),
    .Y(_13793_));
 AOI21x1_ASAP7_75t_SL _22057_ (.A1(_13712_),
    .A2(_13793_),
    .B(_13582_),
    .Y(_13794_));
 NAND2x1_ASAP7_75t_SL _22058_ (.A(_13792_),
    .B(_13794_),
    .Y(_13795_));
 NOR2x2_ASAP7_75t_SL _22059_ (.A(_13513_),
    .B(_13531_),
    .Y(_13796_));
 INVx1_ASAP7_75t_R _22060_ (.A(_13538_),
    .Y(_13797_));
 NAND2x1_ASAP7_75t_SL _22061_ (.A(_13796_),
    .B(_13797_),
    .Y(_13798_));
 NOR2x1_ASAP7_75t_SL _22062_ (.A(_13471_),
    .B(_13510_),
    .Y(_13799_));
 OAI21x1_ASAP7_75t_SL _22063_ (.A1(_13799_),
    .A2(_13644_),
    .B(_13531_),
    .Y(_13800_));
 AOI21x1_ASAP7_75t_SL _22064_ (.A1(_13798_),
    .A2(_13800_),
    .B(_13597_),
    .Y(_13801_));
 OAI21x1_ASAP7_75t_SL _22065_ (.A1(_13732_),
    .A2(_13533_),
    .B(_13531_),
    .Y(_13802_));
 OAI21x1_ASAP7_75t_SL _22066_ (.A1(_13510_),
    .A2(_13513_),
    .B(_13645_),
    .Y(_13803_));
 NAND2x1_ASAP7_75t_SL _22067_ (.A(_13542_),
    .B(_13803_),
    .Y(_13804_));
 AOI21x1_ASAP7_75t_SL _22068_ (.A1(_13802_),
    .A2(_13804_),
    .B(_13560_),
    .Y(_13805_));
 OAI21x1_ASAP7_75t_SL _22069_ (.A1(_13801_),
    .A2(_13805_),
    .B(_13582_),
    .Y(_13806_));
 AOI21x1_ASAP7_75t_SL _22070_ (.A1(_13795_),
    .A2(_13806_),
    .B(_13694_),
    .Y(_13807_));
 OAI21x1_ASAP7_75t_SL _22071_ (.A1(_13788_),
    .A2(_13807_),
    .B(_13623_),
    .Y(_13808_));
 NAND2x1_ASAP7_75t_SL _22072_ (.A(_13769_),
    .B(_13808_),
    .Y(_00065_));
 NAND2x1_ASAP7_75t_SL _22073_ (.A(_01150_),
    .B(_13507_),
    .Y(_13809_));
 AOI21x1_ASAP7_75t_SL _22074_ (.A1(_13809_),
    .A2(_13683_),
    .B(_13531_),
    .Y(_13810_));
 NOR2x1_ASAP7_75t_SL _22075_ (.A(_13597_),
    .B(_13810_),
    .Y(_13811_));
 NOR2x1_ASAP7_75t_SL _22076_ (.A(_01155_),
    .B(_13513_),
    .Y(_13812_));
 OAI21x1_ASAP7_75t_SL _22077_ (.A1(_13812_),
    .A2(_13732_),
    .B(_13531_),
    .Y(_13813_));
 NAND2x1_ASAP7_75t_SL _22078_ (.A(_13471_),
    .B(_13513_),
    .Y(_13814_));
 NAND2x1_ASAP7_75t_SL _22079_ (.A(_13814_),
    .B(_13629_),
    .Y(_13815_));
 AOI21x1_ASAP7_75t_SL _22080_ (.A1(_13813_),
    .A2(_13815_),
    .B(_13560_),
    .Y(_13816_));
 AOI21x1_ASAP7_75t_SL _22081_ (.A1(_13703_),
    .A2(_13811_),
    .B(_13816_),
    .Y(_13817_));
 NOR2x1_ASAP7_75t_SL _22082_ (.A(_13471_),
    .B(_13513_),
    .Y(_13818_));
 OAI21x1_ASAP7_75t_SL _22083_ (.A1(_13646_),
    .A2(_13818_),
    .B(_13745_),
    .Y(_13819_));
 AND3x1_ASAP7_75t_SL _22084_ (.A(_13729_),
    .B(_13542_),
    .C(_13749_),
    .Y(_13820_));
 OAI21x1_ASAP7_75t_SL _22085_ (.A1(_13820_),
    .A2(_13819_),
    .B(_13613_),
    .Y(_13821_));
 AO21x1_ASAP7_75t_SL _22086_ (.A1(_13538_),
    .A2(_13507_),
    .B(_13542_),
    .Y(_13822_));
 NAND2x1_ASAP7_75t_SL _22087_ (.A(_13589_),
    .B(_13513_),
    .Y(_13823_));
 AO21x1_ASAP7_75t_SL _22088_ (.A1(_13752_),
    .A2(_13823_),
    .B(_13531_),
    .Y(_13824_));
 NOR2x1_ASAP7_75t_SL _22089_ (.A(_13597_),
    .B(_13605_),
    .Y(_13825_));
 INVx1_ASAP7_75t_SL _22090_ (.A(_13825_),
    .Y(_13826_));
 AOI21x1_ASAP7_75t_SL _22091_ (.A1(_13822_),
    .A2(_13824_),
    .B(_13826_),
    .Y(_13827_));
 NOR2x1_ASAP7_75t_SL _22092_ (.A(_13827_),
    .B(_13821_),
    .Y(_13828_));
 OAI21x1_ASAP7_75t_SL _22093_ (.A1(_13582_),
    .A2(_13817_),
    .B(_13828_),
    .Y(_13829_));
 AO21x1_ASAP7_75t_SL _22094_ (.A1(_13814_),
    .A2(_13711_),
    .B(_13531_),
    .Y(_13830_));
 NOR2x1_ASAP7_75t_SL _22095_ (.A(_13718_),
    .B(_13714_),
    .Y(_13831_));
 AOI21x1_ASAP7_75t_SL _22096_ (.A1(_13830_),
    .A2(_13831_),
    .B(_13582_),
    .Y(_13832_));
 NOR2x1_ASAP7_75t_R _22097_ (.A(_01153_),
    .B(_13507_),
    .Y(_13833_));
 NAND2x1_ASAP7_75t_SL _22098_ (.A(_13589_),
    .B(_13507_),
    .Y(_13834_));
 NAND2x1_ASAP7_75t_SL _22099_ (.A(_13531_),
    .B(_13834_),
    .Y(_13835_));
 NOR2x1_ASAP7_75t_SL _22100_ (.A(_13833_),
    .B(_13835_),
    .Y(_13836_));
 AND3x1_ASAP7_75t_SL _22101_ (.A(_13729_),
    .B(_13542_),
    .C(_13711_),
    .Y(_13837_));
 OAI21x1_ASAP7_75t_SL _22102_ (.A1(_13836_),
    .A2(_13837_),
    .B(_13597_),
    .Y(_13838_));
 NAND2x1_ASAP7_75t_SL _22103_ (.A(_13832_),
    .B(_13838_),
    .Y(_13839_));
 NAND2x2_ASAP7_75t_SL _22104_ (.A(_13510_),
    .B(_13513_),
    .Y(_13840_));
 INVx1_ASAP7_75t_SL _22105_ (.A(_13689_),
    .Y(_13841_));
 NAND3x1_ASAP7_75t_SL _22106_ (.A(_13840_),
    .B(_13841_),
    .C(_13531_),
    .Y(_13842_));
 AO21x1_ASAP7_75t_SL _22107_ (.A1(_13645_),
    .A2(_13650_),
    .B(_13531_),
    .Y(_13843_));
 AOI21x1_ASAP7_75t_SL _22108_ (.A1(_13842_),
    .A2(_13843_),
    .B(_13826_),
    .Y(_13844_));
 OAI21x1_ASAP7_75t_SL _22109_ (.A1(_13704_),
    .A2(_13835_),
    .B(_13597_),
    .Y(_13845_));
 NAND2x1_ASAP7_75t_SL _22110_ (.A(_13542_),
    .B(_13713_),
    .Y(_13846_));
 OAI21x1_ASAP7_75t_SL _22111_ (.A1(_13818_),
    .A2(_13846_),
    .B(_13582_),
    .Y(_13847_));
 OAI21x1_ASAP7_75t_SL _22112_ (.A1(_13845_),
    .A2(_13847_),
    .B(_13694_),
    .Y(_13848_));
 NOR2x1_ASAP7_75t_SL _22113_ (.A(_13848_),
    .B(_13844_),
    .Y(_13849_));
 AOI21x1_ASAP7_75t_SL _22114_ (.A1(_13849_),
    .A2(_13839_),
    .B(_13623_),
    .Y(_13850_));
 NAND2x1_ASAP7_75t_SL _22115_ (.A(_13829_),
    .B(_13850_),
    .Y(_13851_));
 NAND2x1_ASAP7_75t_SL _22116_ (.A(_01159_),
    .B(_13542_),
    .Y(_13852_));
 AOI21x1_ASAP7_75t_SL _22117_ (.A1(_13852_),
    .A2(_13822_),
    .B(_13597_),
    .Y(_13853_));
 NOR2x1_ASAP7_75t_SL _22118_ (.A(_01164_),
    .B(_13542_),
    .Y(_13854_));
 AOI21x1_ASAP7_75t_SL _22119_ (.A1(_13814_),
    .A2(_13629_),
    .B(_13854_),
    .Y(_13855_));
 OAI21x1_ASAP7_75t_SL _22120_ (.A1(_13560_),
    .A2(_13855_),
    .B(_13613_),
    .Y(_13856_));
 NOR2x1_ASAP7_75t_SL _22121_ (.A(_13853_),
    .B(_13856_),
    .Y(_13857_));
 NOR2x1_ASAP7_75t_SL _22122_ (.A(_13638_),
    .B(_13507_),
    .Y(_13858_));
 NAND2x1p5_ASAP7_75t_SL _22123_ (.A(_13542_),
    .B(_13678_),
    .Y(_13859_));
 NOR2x1_ASAP7_75t_SL _22124_ (.A(_13858_),
    .B(_13859_),
    .Y(_13860_));
 NOR2x1_ASAP7_75t_SL _22125_ (.A(_13537_),
    .B(_13507_),
    .Y(_13861_));
 NOR3x1_ASAP7_75t_SL _22126_ (.A(_13861_),
    .B(_13763_),
    .C(_13542_),
    .Y(_13862_));
 OAI21x1_ASAP7_75t_SL _22127_ (.A1(_13862_),
    .A2(_13860_),
    .B(_13597_),
    .Y(_13863_));
 NAND2x1_ASAP7_75t_SL _22128_ (.A(_01162_),
    .B(_13531_),
    .Y(_13864_));
 NOR2x2_ASAP7_75t_SL _22129_ (.A(_13471_),
    .B(_13489_),
    .Y(_13865_));
 NOR2x1_ASAP7_75t_SL _22130_ (.A(_13865_),
    .B(_13861_),
    .Y(_13866_));
 AOI21x1_ASAP7_75t_SL _22131_ (.A1(_13542_),
    .A2(_13866_),
    .B(_13597_),
    .Y(_13867_));
 NAND2x1_ASAP7_75t_SL _22132_ (.A(_13864_),
    .B(_13867_),
    .Y(_13868_));
 AOI21x1_ASAP7_75t_SL _22133_ (.A1(_13868_),
    .A2(_13863_),
    .B(_13613_),
    .Y(_13869_));
 OAI21x1_ASAP7_75t_SL _22134_ (.A1(_13869_),
    .A2(_13857_),
    .B(_13605_),
    .Y(_13870_));
 NAND2x1_ASAP7_75t_SL _22135_ (.A(_13542_),
    .B(_13840_),
    .Y(_13871_));
 OAI21x1_ASAP7_75t_SL _22136_ (.A1(_13871_),
    .A2(_13818_),
    .B(_13703_),
    .Y(_13872_));
 OA21x2_ASAP7_75t_SL _22137_ (.A1(_13542_),
    .A2(_01160_),
    .B(_13560_),
    .Y(_13873_));
 NAND2x1_ASAP7_75t_SL _22138_ (.A(_13683_),
    .B(_13790_),
    .Y(_13874_));
 AOI21x1_ASAP7_75t_SL _22139_ (.A1(_13873_),
    .A2(_13874_),
    .B(_13613_),
    .Y(_13875_));
 OAI21x1_ASAP7_75t_SL _22140_ (.A1(_13560_),
    .A2(_13872_),
    .B(_13875_),
    .Y(_13876_));
 AO21x1_ASAP7_75t_SL _22141_ (.A1(_13645_),
    .A2(_13711_),
    .B(_13531_),
    .Y(_13877_));
 NOR2x1_ASAP7_75t_SL _22142_ (.A(_13656_),
    .B(_13542_),
    .Y(_13878_));
 NOR2x1_ASAP7_75t_SL _22143_ (.A(_13597_),
    .B(_13878_),
    .Y(_13879_));
 AOI21x1_ASAP7_75t_SL _22144_ (.A1(_13877_),
    .A2(_13879_),
    .B(_13694_),
    .Y(_13880_));
 NOR2x1_ASAP7_75t_SL _22145_ (.A(_13670_),
    .B(_13507_),
    .Y(_13881_));
 AOI21x1_ASAP7_75t_R _22146_ (.A1(_13471_),
    .A2(_13489_),
    .B(_13513_),
    .Y(_13882_));
 OAI21x1_ASAP7_75t_SL _22147_ (.A1(_13881_),
    .A2(_13882_),
    .B(_13542_),
    .Y(_13883_));
 AOI21x1_ASAP7_75t_SL _22148_ (.A1(_13684_),
    .A2(_13571_),
    .B(_13560_),
    .Y(_13884_));
 NAND2x1_ASAP7_75t_SL _22149_ (.A(_13883_),
    .B(_13884_),
    .Y(_13885_));
 AOI21x1_ASAP7_75t_SL _22150_ (.A1(_13885_),
    .A2(_13880_),
    .B(_13605_),
    .Y(_13886_));
 AOI21x1_ASAP7_75t_SL _22151_ (.A1(_13886_),
    .A2(_13876_),
    .B(_13622_),
    .Y(_13887_));
 NAND2x1_ASAP7_75t_SL _22152_ (.A(_13870_),
    .B(_13887_),
    .Y(_13888_));
 NAND2x1_ASAP7_75t_SL _22153_ (.A(_13888_),
    .B(_13851_),
    .Y(_00066_));
 NAND2x1_ASAP7_75t_SL _22154_ (.A(_01152_),
    .B(_13507_),
    .Y(_13889_));
 NAND2x1_ASAP7_75t_SL _22155_ (.A(_13889_),
    .B(_13635_),
    .Y(_13890_));
 NAND2x1_ASAP7_75t_SL _22156_ (.A(_13890_),
    .B(_13630_),
    .Y(_13891_));
 NOR2x1_ASAP7_75t_SL _22157_ (.A(_13531_),
    .B(_13818_),
    .Y(_13892_));
 NOR2x1_ASAP7_75t_SL _22158_ (.A(_13858_),
    .B(_13625_),
    .Y(_13893_));
 NAND2x1_ASAP7_75t_SL _22159_ (.A(_13892_),
    .B(_13893_),
    .Y(_13894_));
 NAND2x1_ASAP7_75t_SL _22160_ (.A(_13678_),
    .B(_13531_),
    .Y(_13895_));
 OA21x2_ASAP7_75t_SL _22161_ (.A1(_13738_),
    .A2(_13895_),
    .B(_13560_),
    .Y(_13896_));
 NAND2x1_ASAP7_75t_SL _22162_ (.A(_13894_),
    .B(_13896_),
    .Y(_13897_));
 AOI21x1_ASAP7_75t_SL _22163_ (.A1(_13891_),
    .A2(_13897_),
    .B(_13613_),
    .Y(_13898_));
 NAND2x1_ASAP7_75t_SL _22164_ (.A(_13656_),
    .B(_13790_),
    .Y(_13899_));
 NAND2x1_ASAP7_75t_SL _22166_ (.A(_13531_),
    .B(_13893_),
    .Y(_13901_));
 AOI21x1_ASAP7_75t_SL _22167_ (.A1(_13899_),
    .A2(_13901_),
    .B(_13560_),
    .Y(_13902_));
 OAI21x1_ASAP7_75t_SL _22168_ (.A1(_13818_),
    .A2(_13646_),
    .B(_13560_),
    .Y(_13903_));
 AND3x1_ASAP7_75t_SL _22169_ (.A(_13809_),
    .B(_13516_),
    .C(_13542_),
    .Y(_13904_));
 OAI21x1_ASAP7_75t_SL _22170_ (.A1(_13903_),
    .A2(_13904_),
    .B(_13613_),
    .Y(_13905_));
 NOR2x1_ASAP7_75t_SL _22171_ (.A(_13902_),
    .B(_13905_),
    .Y(_13906_));
 NOR3x1_ASAP7_75t_SL _22172_ (.A(_13898_),
    .B(_13622_),
    .C(_13906_),
    .Y(_13907_));
 NOR2x1_ASAP7_75t_SL _22173_ (.A(_13542_),
    .B(_13585_),
    .Y(_13908_));
 OA21x2_ASAP7_75t_SL _22174_ (.A1(_13685_),
    .A2(_13908_),
    .B(_13613_),
    .Y(_13909_));
 OA21x2_ASAP7_75t_SL _22175_ (.A1(_13713_),
    .A2(_13531_),
    .B(_13560_),
    .Y(_13910_));
 NAND2x1_ASAP7_75t_SL _22176_ (.A(_13842_),
    .B(_13910_),
    .Y(_13911_));
 AO21x1_ASAP7_75t_SL _22177_ (.A1(_13909_),
    .A2(_13911_),
    .B(_13623_),
    .Y(_13912_));
 INVx1_ASAP7_75t_SL _22178_ (.A(_13590_),
    .Y(_13913_));
 OA21x2_ASAP7_75t_SL _22179_ (.A1(_13533_),
    .A2(_13833_),
    .B(_13542_),
    .Y(_13914_));
 AOI21x1_ASAP7_75t_SL _22180_ (.A1(_13913_),
    .A2(_13635_),
    .B(_13914_),
    .Y(_13915_));
 NAND2x1_ASAP7_75t_SL _22181_ (.A(_13675_),
    .B(_13800_),
    .Y(_13916_));
 OAI21x1_ASAP7_75t_SL _22182_ (.A1(_13597_),
    .A2(_13916_),
    .B(_13694_),
    .Y(_13917_));
 AOI21x1_ASAP7_75t_SL _22183_ (.A1(_13597_),
    .A2(_13915_),
    .B(_13917_),
    .Y(_13918_));
 OAI21x1_ASAP7_75t_SL _22184_ (.A1(_13912_),
    .A2(_13918_),
    .B(_13582_),
    .Y(_13919_));
 INVx2_ASAP7_75t_SL _22185_ (.A(_13646_),
    .Y(_13920_));
 NAND2x1p5_ASAP7_75t_SL _22186_ (.A(_13920_),
    .B(_13841_),
    .Y(_13921_));
 NAND2x1p5_ASAP7_75t_SL _22187_ (.A(_13776_),
    .B(_13921_),
    .Y(_13922_));
 NAND2x1_ASAP7_75t_SL _22188_ (.A(_13513_),
    .B(_13542_),
    .Y(_13923_));
 OAI21x1_ASAP7_75t_SL _22189_ (.A1(_13510_),
    .A2(_13513_),
    .B(_13560_),
    .Y(_13924_));
 NOR2x1_ASAP7_75t_SL _22190_ (.A(_13865_),
    .B(_13924_),
    .Y(_13925_));
 AOI21x1_ASAP7_75t_SL _22191_ (.A1(_13923_),
    .A2(_13925_),
    .B(_13613_),
    .Y(_13926_));
 AOI21x1_ASAP7_75t_SL _22192_ (.A1(_13926_),
    .A2(_13922_),
    .B(_13622_),
    .Y(_13927_));
 NAND2x1_ASAP7_75t_SL _22193_ (.A(_13471_),
    .B(_13507_),
    .Y(_13928_));
 AO21x1_ASAP7_75t_SL _22194_ (.A1(_13729_),
    .A2(_13928_),
    .B(_13542_),
    .Y(_13929_));
 AOI21x1_ASAP7_75t_SL _22195_ (.A1(_13651_),
    .A2(_13929_),
    .B(_13694_),
    .Y(_13930_));
 INVx1_ASAP7_75t_SL _22196_ (.A(_13730_),
    .Y(_13931_));
 NAND2x1_ASAP7_75t_SL _22197_ (.A(_13797_),
    .B(_13931_),
    .Y(_13932_));
 AOI21x1_ASAP7_75t_SL _22198_ (.A1(_13567_),
    .A2(_13715_),
    .B(_13597_),
    .Y(_13933_));
 NAND2x1_ASAP7_75t_SL _22199_ (.A(_13932_),
    .B(_13933_),
    .Y(_13934_));
 NAND2x1_ASAP7_75t_SL _22200_ (.A(_13930_),
    .B(_13934_),
    .Y(_13935_));
 AOI21x1_ASAP7_75t_SL _22201_ (.A1(_13935_),
    .A2(_13927_),
    .B(_13582_),
    .Y(_13936_));
 NAND2x1_ASAP7_75t_SL _22202_ (.A(_13694_),
    .B(_13845_),
    .Y(_13937_));
 NAND2x1_ASAP7_75t_SL _22203_ (.A(_13670_),
    .B(_13513_),
    .Y(_13938_));
 NAND2x1_ASAP7_75t_SL _22204_ (.A(_13938_),
    .B(_13690_),
    .Y(_13939_));
 AOI21x1_ASAP7_75t_SL _22205_ (.A1(_13939_),
    .A2(_13727_),
    .B(_13597_),
    .Y(_13940_));
 NOR2x1_ASAP7_75t_SL _22206_ (.A(_13937_),
    .B(_13940_),
    .Y(_13941_));
 NAND2x1_ASAP7_75t_SL _22207_ (.A(_13814_),
    .B(_13684_),
    .Y(_13942_));
 NOR2x1_ASAP7_75t_SL _22208_ (.A(_13531_),
    .B(_13650_),
    .Y(_13943_));
 NOR2x1_ASAP7_75t_SL _22209_ (.A(_13943_),
    .B(_13685_),
    .Y(_13944_));
 NAND2x1_ASAP7_75t_SL _22210_ (.A(_13942_),
    .B(_13944_),
    .Y(_13945_));
 OAI21x1_ASAP7_75t_SL _22211_ (.A1(_13812_),
    .A2(_13881_),
    .B(_13542_),
    .Y(_13946_));
 AOI21x1_ASAP7_75t_SL _22212_ (.A1(_13531_),
    .A2(_13803_),
    .B(_13597_),
    .Y(_13947_));
 NAND2x1_ASAP7_75t_SL _22213_ (.A(_13946_),
    .B(_13947_),
    .Y(_13948_));
 AOI21x1_ASAP7_75t_SL _22214_ (.A1(_13945_),
    .A2(_13948_),
    .B(_13694_),
    .Y(_13949_));
 OAI21x1_ASAP7_75t_SL _22215_ (.A1(_13941_),
    .A2(_13949_),
    .B(_13622_),
    .Y(_13950_));
 NAND2x1_ASAP7_75t_SL _22216_ (.A(_13950_),
    .B(_13936_),
    .Y(_13951_));
 OAI21x1_ASAP7_75t_SL _22217_ (.A1(_13907_),
    .A2(_13919_),
    .B(_13951_),
    .Y(_00067_));
 OAI21x1_ASAP7_75t_SL _22218_ (.A1(_13865_),
    .A2(_13704_),
    .B(_13542_),
    .Y(_13952_));
 NAND2x1_ASAP7_75t_R _22219_ (.A(_13565_),
    .B(_13639_),
    .Y(_13953_));
 AOI21x1_ASAP7_75t_R _22220_ (.A1(_13531_),
    .A2(_13953_),
    .B(_13597_),
    .Y(_13954_));
 NAND2x1_ASAP7_75t_R _22221_ (.A(_13952_),
    .B(_13954_),
    .Y(_13955_));
 NAND2x1_ASAP7_75t_R _22222_ (.A(_13471_),
    .B(_13489_),
    .Y(_13956_));
 AOI21x1_ASAP7_75t_SL _22223_ (.A1(_13956_),
    .A2(_13774_),
    .B(_13542_),
    .Y(_13957_));
 INVx1_ASAP7_75t_R _22224_ (.A(_13957_),
    .Y(_13958_));
 AOI21x1_ASAP7_75t_R _22225_ (.A1(_13729_),
    .A2(_13690_),
    .B(_13560_),
    .Y(_13959_));
 NAND2x1_ASAP7_75t_R _22226_ (.A(_13958_),
    .B(_13959_),
    .Y(_13960_));
 AOI21x1_ASAP7_75t_R _22227_ (.A1(_13955_),
    .A2(_13960_),
    .B(_13582_),
    .Y(_13961_));
 NAND2x1_ASAP7_75t_SL _22228_ (.A(_13774_),
    .B(_13690_),
    .Y(_13962_));
 INVx1_ASAP7_75t_SL _22229_ (.A(_13962_),
    .Y(_13963_));
 NAND2x1_ASAP7_75t_SL _22230_ (.A(_13531_),
    .B(_13704_),
    .Y(_13964_));
 NAND2x1_ASAP7_75t_SL _22231_ (.A(_13531_),
    .B(_13544_),
    .Y(_13965_));
 NAND3x1_ASAP7_75t_R _22232_ (.A(_13964_),
    .B(_13965_),
    .C(_13745_),
    .Y(_13966_));
 NAND2x1_ASAP7_75t_R _22233_ (.A(_01154_),
    .B(_13531_),
    .Y(_13967_));
 NAND2x1_ASAP7_75t_L _22234_ (.A(_13967_),
    .B(_13859_),
    .Y(_13968_));
 OA21x2_ASAP7_75t_SL _22235_ (.A1(_13968_),
    .A2(_13826_),
    .B(_13622_),
    .Y(_13969_));
 OAI21x1_ASAP7_75t_SL _22236_ (.A1(_13963_),
    .A2(_13966_),
    .B(_13969_),
    .Y(_13970_));
 OAI21x1_ASAP7_75t_SL _22237_ (.A1(_13970_),
    .A2(_13961_),
    .B(_13613_),
    .Y(_13971_));
 AND3x1_ASAP7_75t_R _22238_ (.A(_13650_),
    .B(_13516_),
    .C(_13531_),
    .Y(_13972_));
 AO21x1_ASAP7_75t_R _22239_ (.A1(_13683_),
    .A2(_13690_),
    .B(_13597_),
    .Y(_13973_));
 OA21x2_ASAP7_75t_SL _22240_ (.A1(_13678_),
    .A2(_13531_),
    .B(_13713_),
    .Y(_13974_));
 AOI21x1_ASAP7_75t_SL _22241_ (.A1(_13712_),
    .A2(_13974_),
    .B(_13605_),
    .Y(_13975_));
 OAI21x1_ASAP7_75t_SL _22242_ (.A1(_13972_),
    .A2(_13973_),
    .B(_13975_),
    .Y(_13976_));
 NAND2x1_ASAP7_75t_SL _22243_ (.A(_13656_),
    .B(_13928_),
    .Y(_13977_));
 AOI21x1_ASAP7_75t_R _22244_ (.A1(_13542_),
    .A2(_13977_),
    .B(_13597_),
    .Y(_13978_));
 AOI21x1_ASAP7_75t_R _22245_ (.A1(_13789_),
    .A2(_13978_),
    .B(_13582_),
    .Y(_13979_));
 NAND2x1_ASAP7_75t_SL _22246_ (.A(_13683_),
    .B(_13892_),
    .Y(_13980_));
 NAND3x1_ASAP7_75t_SL _22247_ (.A(_13980_),
    .B(_13597_),
    .C(_13813_),
    .Y(_13981_));
 NAND2x1_ASAP7_75t_SL _22248_ (.A(_13979_),
    .B(_13981_),
    .Y(_13982_));
 AOI21x1_ASAP7_75t_SL _22249_ (.A1(_13982_),
    .A2(_13976_),
    .B(_13622_),
    .Y(_13983_));
 NOR2x1_ASAP7_75t_SL _22250_ (.A(_13971_),
    .B(_13983_),
    .Y(_13984_));
 AO21x1_ASAP7_75t_R _22251_ (.A1(_13534_),
    .A2(_13571_),
    .B(_13597_),
    .Y(_13985_));
 INVx2_ASAP7_75t_R _22252_ (.A(_13678_),
    .Y(_13986_));
 AO21x1_ASAP7_75t_SL _22253_ (.A1(_01150_),
    .A2(_13513_),
    .B(_13542_),
    .Y(_13987_));
 OAI21x1_ASAP7_75t_R _22254_ (.A1(_13986_),
    .A2(_13987_),
    .B(_13582_),
    .Y(_13988_));
 AO21x1_ASAP7_75t_R _22255_ (.A1(_13570_),
    .A2(_13507_),
    .B(_13531_),
    .Y(_13989_));
 NAND2x1_ASAP7_75t_SL _22256_ (.A(_13597_),
    .B(_13582_),
    .Y(_13990_));
 OA21x2_ASAP7_75t_SL _22257_ (.A1(_13564_),
    .A2(_13513_),
    .B(_13531_),
    .Y(_13991_));
 NOR2x1_ASAP7_75t_SL _22258_ (.A(_13990_),
    .B(_13991_),
    .Y(_13992_));
 AOI21x1_ASAP7_75t_R _22259_ (.A1(_13989_),
    .A2(_13992_),
    .B(_13623_),
    .Y(_13993_));
 OAI21x1_ASAP7_75t_R _22260_ (.A1(_13985_),
    .A2(_13988_),
    .B(_13993_),
    .Y(_13994_));
 AO21x1_ASAP7_75t_R _22261_ (.A1(_13542_),
    .A2(_13507_),
    .B(_13597_),
    .Y(_13995_));
 AO21x1_ASAP7_75t_R _22262_ (.A1(_13931_),
    .A2(_13913_),
    .B(_13995_),
    .Y(_13996_));
 AO21x1_ASAP7_75t_R _22263_ (.A1(_13567_),
    .A2(_13656_),
    .B(_13542_),
    .Y(_13997_));
 NAND3x1_ASAP7_75t_R _22264_ (.A(_13997_),
    .B(_13597_),
    .C(_13734_),
    .Y(_13998_));
 AOI21x1_ASAP7_75t_R _22265_ (.A1(_13996_),
    .A2(_13998_),
    .B(_13582_),
    .Y(_13999_));
 NOR2x1_ASAP7_75t_SL _22266_ (.A(_13994_),
    .B(_13999_),
    .Y(_14000_));
 NAND2x1_ASAP7_75t_SL _22267_ (.A(_13542_),
    .B(_13928_),
    .Y(_14001_));
 NOR2x1_ASAP7_75t_SL _22268_ (.A(_13742_),
    .B(_14001_),
    .Y(_14002_));
 OAI21x1_ASAP7_75t_R _22269_ (.A1(_13742_),
    .A2(_13744_),
    .B(_13825_),
    .Y(_14003_));
 INVx1_ASAP7_75t_R _22270_ (.A(_13690_),
    .Y(_14004_));
 NOR2x1_ASAP7_75t_SL _22271_ (.A(_13760_),
    .B(_13990_),
    .Y(_14005_));
 AOI21x1_ASAP7_75t_R _22272_ (.A1(_14004_),
    .A2(_14005_),
    .B(_13622_),
    .Y(_14006_));
 OAI21x1_ASAP7_75t_SL _22273_ (.A1(_14002_),
    .A2(_14003_),
    .B(_14006_),
    .Y(_14007_));
 NAND2x1_ASAP7_75t_SL _22274_ (.A(_13542_),
    .B(_13814_),
    .Y(_14008_));
 NOR2x1_ASAP7_75t_R _22275_ (.A(_13763_),
    .B(_14008_),
    .Y(_14009_));
 OAI21x1_ASAP7_75t_R _22276_ (.A1(_13957_),
    .A2(_14009_),
    .B(_13597_),
    .Y(_14010_));
 AO21x1_ASAP7_75t_R _22277_ (.A1(_13840_),
    .A2(_13567_),
    .B(_13542_),
    .Y(_14011_));
 NAND2x1_ASAP7_75t_SL _22278_ (.A(_14011_),
    .B(_13867_),
    .Y(_14012_));
 AOI21x1_ASAP7_75t_R _22279_ (.A1(_14010_),
    .A2(_14012_),
    .B(_13582_),
    .Y(_14013_));
 OAI21x1_ASAP7_75t_R _22280_ (.A1(_14007_),
    .A2(_14013_),
    .B(_13694_),
    .Y(_14014_));
 NOR2x1_ASAP7_75t_SL _22281_ (.A(_14000_),
    .B(_14014_),
    .Y(_14015_));
 NOR2x1_ASAP7_75t_SL _22282_ (.A(_13984_),
    .B(_14015_),
    .Y(_00068_));
 NOR2x1_ASAP7_75t_SL _22283_ (.A(_13542_),
    .B(_13689_),
    .Y(_14016_));
 AO21x1_ASAP7_75t_SL _22284_ (.A1(_13710_),
    .A2(_13542_),
    .B(_13685_),
    .Y(_14017_));
 AO21x1_ASAP7_75t_SL _22285_ (.A1(_13683_),
    .A2(_14016_),
    .B(_14017_),
    .Y(_14018_));
 AO21x1_ASAP7_75t_SL _22286_ (.A1(_13834_),
    .A2(_13770_),
    .B(_13531_),
    .Y(_14019_));
 AOI21x1_ASAP7_75t_SL _22287_ (.A1(_14019_),
    .A2(_13569_),
    .B(_13605_),
    .Y(_14020_));
 AO21x1_ASAP7_75t_SL _22288_ (.A1(_13585_),
    .A2(_13531_),
    .B(_13597_),
    .Y(_14021_));
 OAI21x1_ASAP7_75t_SL _22289_ (.A1(_14021_),
    .A2(_13914_),
    .B(_13605_),
    .Y(_14022_));
 AND3x1_ASAP7_75t_SL _22290_ (.A(_13798_),
    .B(_13597_),
    .C(_13987_),
    .Y(_14023_));
 OAI21x1_ASAP7_75t_SL _22291_ (.A1(_14022_),
    .A2(_14023_),
    .B(_13694_),
    .Y(_14024_));
 AOI21x1_ASAP7_75t_SL _22292_ (.A1(_14018_),
    .A2(_14020_),
    .B(_14024_),
    .Y(_14025_));
 NOR2x1_ASAP7_75t_SL _22293_ (.A(_13658_),
    .B(_13738_),
    .Y(_14026_));
 OAI21x1_ASAP7_75t_R _22294_ (.A1(_13570_),
    .A2(_13533_),
    .B(_13531_),
    .Y(_14027_));
 OAI21x1_ASAP7_75t_SL _22295_ (.A1(_13531_),
    .A2(_14026_),
    .B(_14027_),
    .Y(_14028_));
 NOR2x1_ASAP7_75t_R _22296_ (.A(_13471_),
    .B(_13531_),
    .Y(_14029_));
 OAI21x1_ASAP7_75t_SL _22297_ (.A1(_14029_),
    .A2(_13957_),
    .B(_13825_),
    .Y(_14030_));
 OAI21x1_ASAP7_75t_SL _22298_ (.A1(_13990_),
    .A2(_14028_),
    .B(_14030_),
    .Y(_14031_));
 NAND2x1_ASAP7_75t_R _22299_ (.A(_13542_),
    .B(_13986_),
    .Y(_14032_));
 AO21x1_ASAP7_75t_L _22300_ (.A1(_13774_),
    .A2(_13749_),
    .B(_13542_),
    .Y(_14033_));
 AOI21x1_ASAP7_75t_SL _22301_ (.A1(_14032_),
    .A2(_14033_),
    .B(_13560_),
    .Y(_14034_));
 AO21x1_ASAP7_75t_R _22302_ (.A1(_13834_),
    .A2(_13531_),
    .B(_13597_),
    .Y(_14035_));
 AND3x1_ASAP7_75t_SL _22303_ (.A(_13585_),
    .B(_13542_),
    .C(_13639_),
    .Y(_14036_));
 OAI21x1_ASAP7_75t_SL _22304_ (.A1(_14035_),
    .A2(_14036_),
    .B(_13605_),
    .Y(_14037_));
 NOR2x1_ASAP7_75t_SL _22305_ (.A(_14034_),
    .B(_14037_),
    .Y(_14038_));
 OAI21x1_ASAP7_75t_SL _22306_ (.A1(_14031_),
    .A2(_14038_),
    .B(_13613_),
    .Y(_14039_));
 NAND2x1_ASAP7_75t_SL _22307_ (.A(_13623_),
    .B(_14039_),
    .Y(_14040_));
 INVx1_ASAP7_75t_R _22308_ (.A(_13591_),
    .Y(_14041_));
 AOI21x1_ASAP7_75t_SL _22309_ (.A1(_14041_),
    .A2(_13712_),
    .B(_13605_),
    .Y(_14042_));
 INVx1_ASAP7_75t_SL _22310_ (.A(_13571_),
    .Y(_14043_));
 AOI21x1_ASAP7_75t_SL _22311_ (.A1(_13542_),
    .A2(_13938_),
    .B(_13597_),
    .Y(_14044_));
 OAI21x1_ASAP7_75t_SL _22312_ (.A1(_14043_),
    .A2(_13822_),
    .B(_14044_),
    .Y(_14045_));
 AOI21x1_ASAP7_75t_SL _22313_ (.A1(_14042_),
    .A2(_14045_),
    .B(_13694_),
    .Y(_14046_));
 NAND2x1p5_ASAP7_75t_SL _22314_ (.A(_13913_),
    .B(_13920_),
    .Y(_14047_));
 AO21x1_ASAP7_75t_SL _22315_ (.A1(_13889_),
    .A2(_13645_),
    .B(_13531_),
    .Y(_14048_));
 AOI21x1_ASAP7_75t_SL _22316_ (.A1(_14048_),
    .A2(_14047_),
    .B(_13560_),
    .Y(_14049_));
 AO21x1_ASAP7_75t_SL _22317_ (.A1(_13541_),
    .A2(_13540_),
    .B(_13638_),
    .Y(_14050_));
 AO21x1_ASAP7_75t_SL _22318_ (.A1(_13570_),
    .A2(_13513_),
    .B(_13542_),
    .Y(_14051_));
 AOI21x1_ASAP7_75t_SL _22319_ (.A1(_14050_),
    .A2(_14051_),
    .B(_13597_),
    .Y(_14052_));
 OAI21x1_ASAP7_75t_SL _22320_ (.A1(_14052_),
    .A2(_14049_),
    .B(_13605_),
    .Y(_14053_));
 NAND2x1_ASAP7_75t_SL _22321_ (.A(_14046_),
    .B(_14053_),
    .Y(_14054_));
 OA21x2_ASAP7_75t_SL _22322_ (.A1(_13531_),
    .A2(_13510_),
    .B(_13560_),
    .Y(_14055_));
 AOI21x1_ASAP7_75t_SL _22323_ (.A1(_14055_),
    .A2(_13627_),
    .B(_13605_),
    .Y(_14056_));
 AOI21x1_ASAP7_75t_SL _22324_ (.A1(_13774_),
    .A2(_14016_),
    .B(_13560_),
    .Y(_14057_));
 NAND2x1_ASAP7_75t_SL _22325_ (.A(_13539_),
    .B(_13715_),
    .Y(_14058_));
 NAND2x1_ASAP7_75t_SL _22326_ (.A(_14057_),
    .B(_14058_),
    .Y(_14059_));
 AOI21x1_ASAP7_75t_SL _22327_ (.A1(_14056_),
    .A2(_14059_),
    .B(_13613_),
    .Y(_14060_));
 OAI21x1_ASAP7_75t_SL _22328_ (.A1(_13812_),
    .A2(_13738_),
    .B(_13531_),
    .Y(_14061_));
 OA21x2_ASAP7_75t_SL _22329_ (.A1(_13889_),
    .A2(_13531_),
    .B(_13597_),
    .Y(_14062_));
 AOI21x1_ASAP7_75t_SL _22330_ (.A1(_14061_),
    .A2(_14062_),
    .B(_13582_),
    .Y(_14063_));
 NAND2x1_ASAP7_75t_SL _22331_ (.A(_13964_),
    .B(_13719_),
    .Y(_14064_));
 NAND2x1_ASAP7_75t_SL _22332_ (.A(_14063_),
    .B(_14064_),
    .Y(_14065_));
 AOI21x1_ASAP7_75t_SL _22333_ (.A1(_14060_),
    .A2(_14065_),
    .B(_13623_),
    .Y(_14066_));
 NAND2x1_ASAP7_75t_SL _22334_ (.A(_14054_),
    .B(_14066_),
    .Y(_14067_));
 OAI21x1_ASAP7_75t_SL _22335_ (.A1(_14025_),
    .A2(_14040_),
    .B(_14067_),
    .Y(_00069_));
 AOI21x1_ASAP7_75t_SL _22336_ (.A1(_13510_),
    .A2(_13796_),
    .B(_13597_),
    .Y(_14068_));
 NAND2x1p5_ASAP7_75t_SL _22337_ (.A(_13846_),
    .B(_13646_),
    .Y(_14069_));
 NAND2x1_ASAP7_75t_SL _22338_ (.A(_14069_),
    .B(_14068_),
    .Y(_14070_));
 NAND2x1_ASAP7_75t_SL _22339_ (.A(_14001_),
    .B(_13595_),
    .Y(_14071_));
 AOI21x1_ASAP7_75t_SL _22340_ (.A1(_14071_),
    .A2(_14070_),
    .B(_13613_),
    .Y(_14072_));
 INVx1_ASAP7_75t_SL _22341_ (.A(_13684_),
    .Y(_14073_));
 AOI21x1_ASAP7_75t_SL _22342_ (.A1(_14073_),
    .A2(_13962_),
    .B(_13560_),
    .Y(_14074_));
 OAI21x1_ASAP7_75t_SL _22343_ (.A1(_13597_),
    .A2(_13810_),
    .B(_13613_),
    .Y(_14075_));
 NOR2x1_ASAP7_75t_SL _22344_ (.A(_14074_),
    .B(_14075_),
    .Y(_14076_));
 OAI21x1_ASAP7_75t_SL _22345_ (.A1(_14076_),
    .A2(_14072_),
    .B(_13605_),
    .Y(_14077_));
 AO21x1_ASAP7_75t_SL _22346_ (.A1(_13542_),
    .A2(_01158_),
    .B(_13597_),
    .Y(_14078_));
 AO21x1_ASAP7_75t_SL _22347_ (.A1(_13774_),
    .A2(_14016_),
    .B(_14078_),
    .Y(_14079_));
 NAND2x1_ASAP7_75t_SL _22348_ (.A(_13591_),
    .B(_13645_),
    .Y(_14080_));
 OA21x2_ASAP7_75t_SL _22349_ (.A1(_13628_),
    .A2(_13542_),
    .B(_13597_),
    .Y(_14081_));
 AOI21x1_ASAP7_75t_SL _22350_ (.A1(_14080_),
    .A2(_14081_),
    .B(_13694_),
    .Y(_14082_));
 NAND2x1_ASAP7_75t_SL _22351_ (.A(_14079_),
    .B(_14082_),
    .Y(_14083_));
 NAND2x1_ASAP7_75t_SL _22352_ (.A(_13537_),
    .B(_13531_),
    .Y(_14084_));
 AOI21x1_ASAP7_75t_SL _22353_ (.A1(_14084_),
    .A2(_13925_),
    .B(_13613_),
    .Y(_14085_));
 NOR2x1_ASAP7_75t_SL _22354_ (.A(_13531_),
    .B(_13865_),
    .Y(_14086_));
 NOR2x1_ASAP7_75t_SL _22355_ (.A(_13589_),
    .B(_13507_),
    .Y(_14087_));
 NOR2x1_ASAP7_75t_SL _22356_ (.A(_13542_),
    .B(_14087_),
    .Y(_14088_));
 NOR2x1_ASAP7_75t_SL _22357_ (.A(_14086_),
    .B(_14088_),
    .Y(_14089_));
 OAI21x1_ASAP7_75t_SL _22358_ (.A1(_13625_),
    .A2(_14089_),
    .B(_13597_),
    .Y(_14090_));
 AOI21x1_ASAP7_75t_SL _22359_ (.A1(_14085_),
    .A2(_14090_),
    .B(_13605_),
    .Y(_14091_));
 AOI21x1_ASAP7_75t_SL _22360_ (.A1(_14083_),
    .A2(_14091_),
    .B(_13623_),
    .Y(_14092_));
 NAND2x1_ASAP7_75t_SL _22361_ (.A(_14077_),
    .B(_14092_),
    .Y(_14093_));
 AO21x1_ASAP7_75t_SL _22362_ (.A1(_13538_),
    .A2(_13507_),
    .B(_13531_),
    .Y(_14094_));
 AO21x1_ASAP7_75t_SL _22363_ (.A1(_13585_),
    .A2(_13749_),
    .B(_13542_),
    .Y(_14095_));
 OAI21x1_ASAP7_75t_SL _22364_ (.A1(_13544_),
    .A2(_14094_),
    .B(_14095_),
    .Y(_14096_));
 OAI21x1_ASAP7_75t_SL _22365_ (.A1(_13542_),
    .A2(_13585_),
    .B(_13597_),
    .Y(_14097_));
 AOI21x1_ASAP7_75t_SL _22366_ (.A1(_13852_),
    .A2(_13822_),
    .B(_14097_),
    .Y(_14098_));
 AOI21x1_ASAP7_75t_SL _22367_ (.A1(_13560_),
    .A2(_14096_),
    .B(_14098_),
    .Y(_14099_));
 NAND2x1_ASAP7_75t_SL _22368_ (.A(_01157_),
    .B(_01163_),
    .Y(_14100_));
 AO21x1_ASAP7_75t_SL _22369_ (.A1(_13531_),
    .A2(_14100_),
    .B(_13597_),
    .Y(_14101_));
 AO21x1_ASAP7_75t_SL _22370_ (.A1(_13797_),
    .A2(_13892_),
    .B(_14101_),
    .Y(_14102_));
 AOI21x1_ASAP7_75t_SL _22371_ (.A1(_13564_),
    .A2(_13796_),
    .B(_13878_),
    .Y(_14103_));
 OA21x2_ASAP7_75t_SL _22372_ (.A1(_13713_),
    .A2(_13531_),
    .B(_13597_),
    .Y(_14104_));
 AOI21x1_ASAP7_75t_SL _22373_ (.A1(_14103_),
    .A2(_14104_),
    .B(_13613_),
    .Y(_14105_));
 AOI21x1_ASAP7_75t_SL _22374_ (.A1(_14102_),
    .A2(_14105_),
    .B(_13605_),
    .Y(_14106_));
 OAI21x1_ASAP7_75t_SL _22375_ (.A1(_13694_),
    .A2(_14099_),
    .B(_14106_),
    .Y(_14107_));
 NAND2x1_ASAP7_75t_SL _22376_ (.A(_13516_),
    .B(_14016_),
    .Y(_14108_));
 OAI21x1_ASAP7_75t_SL _22377_ (.A1(_13760_),
    .A2(_13882_),
    .B(_13542_),
    .Y(_14109_));
 AOI21x1_ASAP7_75t_SL _22378_ (.A1(_14108_),
    .A2(_14109_),
    .B(_13597_),
    .Y(_14110_));
 NOR2x1_ASAP7_75t_SL _22379_ (.A(_13671_),
    .B(_13846_),
    .Y(_14111_));
 NAND2x1_ASAP7_75t_SL _22380_ (.A(_13964_),
    .B(_13679_),
    .Y(_14112_));
 NOR2x1_ASAP7_75t_SL _22381_ (.A(_14111_),
    .B(_14112_),
    .Y(_14113_));
 OAI21x1_ASAP7_75t_SL _22382_ (.A1(_14113_),
    .A2(_14110_),
    .B(_13694_),
    .Y(_14114_));
 AO21x1_ASAP7_75t_SL _22383_ (.A1(_13729_),
    .A2(_13471_),
    .B(_13531_),
    .Y(_14115_));
 OA21x2_ASAP7_75t_SL _22384_ (.A1(_13889_),
    .A2(_13542_),
    .B(_13597_),
    .Y(_14116_));
 AOI21x1_ASAP7_75t_SL _22385_ (.A1(_14115_),
    .A2(_14116_),
    .B(_13694_),
    .Y(_14117_));
 OAI21x1_ASAP7_75t_SL _22386_ (.A1(_13702_),
    .A2(_13881_),
    .B(_13531_),
    .Y(_14118_));
 NAND3x1_ASAP7_75t_SL _22387_ (.A(_14068_),
    .B(_13952_),
    .C(_14118_),
    .Y(_14119_));
 AOI21x1_ASAP7_75t_SL _22388_ (.A1(_14117_),
    .A2(_14119_),
    .B(_13582_),
    .Y(_14120_));
 AOI21x1_ASAP7_75t_SL _22389_ (.A1(_14120_),
    .A2(_14114_),
    .B(_13622_),
    .Y(_14121_));
 NAND2x1_ASAP7_75t_SL _22390_ (.A(_14121_),
    .B(_14107_),
    .Y(_14122_));
 NAND2x1_ASAP7_75t_SL _22391_ (.A(_14122_),
    .B(_14093_),
    .Y(_00070_));
 OAI21x1_ASAP7_75t_SL _22392_ (.A1(_14088_),
    .A2(_13963_),
    .B(_13825_),
    .Y(_14123_));
 NAND3x1_ASAP7_75t_SL _22393_ (.A(_13752_),
    .B(_13542_),
    .C(_13656_),
    .Y(_14124_));
 NOR2x1_ASAP7_75t_SL _22394_ (.A(_13489_),
    .B(_13542_),
    .Y(_14125_));
 AOI21x1_ASAP7_75t_SL _22395_ (.A1(_13774_),
    .A2(_14125_),
    .B(_13990_),
    .Y(_14126_));
 AOI21x1_ASAP7_75t_SL _22396_ (.A1(_14124_),
    .A2(_14126_),
    .B(_13613_),
    .Y(_14127_));
 NAND2x1_ASAP7_75t_SL _22397_ (.A(_14123_),
    .B(_14127_),
    .Y(_14128_));
 AND2x2_ASAP7_75t_SL _22398_ (.A(_13803_),
    .B(_13531_),
    .Y(_14129_));
 NAND2x1_ASAP7_75t_SL _22399_ (.A(_13542_),
    .B(_13650_),
    .Y(_14130_));
 OAI21x1_ASAP7_75t_SL _22400_ (.A1(_14087_),
    .A2(_14130_),
    .B(_13597_),
    .Y(_14131_));
 OAI21x1_ASAP7_75t_SL _22401_ (.A1(_14129_),
    .A2(_14131_),
    .B(_13605_),
    .Y(_14132_));
 OAI21x1_ASAP7_75t_SL _22402_ (.A1(_13871_),
    .A2(_13818_),
    .B(_14108_),
    .Y(_14133_));
 NOR2x1_ASAP7_75t_SL _22403_ (.A(_13597_),
    .B(_14133_),
    .Y(_14134_));
 NOR2x1_ASAP7_75t_SL _22404_ (.A(_14132_),
    .B(_14134_),
    .Y(_14135_));
 OAI21x1_ASAP7_75t_SL _22405_ (.A1(_14128_),
    .A2(_14135_),
    .B(_13622_),
    .Y(_14136_));
 NOR2x1_ASAP7_75t_SL _22406_ (.A(_13570_),
    .B(_13923_),
    .Y(_14137_));
 AO21x1_ASAP7_75t_SL _22407_ (.A1(_13634_),
    .A2(_13531_),
    .B(_13597_),
    .Y(_14138_));
 OAI21x1_ASAP7_75t_SL _22408_ (.A1(_14137_),
    .A2(_14138_),
    .B(_13605_),
    .Y(_14139_));
 AO21x1_ASAP7_75t_SL _22409_ (.A1(_13542_),
    .A2(_13507_),
    .B(_13560_),
    .Y(_14140_));
 AOI211x1_ASAP7_75t_SL _22410_ (.A1(_13920_),
    .A2(_13632_),
    .B(_13629_),
    .C(_14140_),
    .Y(_14141_));
 OAI21x1_ASAP7_75t_SL _22411_ (.A1(_14141_),
    .A2(_14139_),
    .B(_13613_),
    .Y(_14142_));
 OAI21x1_ASAP7_75t_SL _22412_ (.A1(_13865_),
    .A2(_14008_),
    .B(_13560_),
    .Y(_14143_));
 AND2x2_ASAP7_75t_SL _22413_ (.A(_13545_),
    .B(_13632_),
    .Y(_14144_));
 OAI21x1_ASAP7_75t_SL _22414_ (.A1(_14143_),
    .A2(_14144_),
    .B(_13582_),
    .Y(_14145_));
 OA21x2_ASAP7_75t_SL _22415_ (.A1(_14002_),
    .A2(_14125_),
    .B(_13597_),
    .Y(_14146_));
 NOR2x1_ASAP7_75t_SL _22416_ (.A(_14145_),
    .B(_14146_),
    .Y(_14147_));
 NOR2x1_ASAP7_75t_SL _22417_ (.A(_14147_),
    .B(_14142_),
    .Y(_14148_));
 AO21x1_ASAP7_75t_SL _22418_ (.A1(_13531_),
    .A2(_13710_),
    .B(_13560_),
    .Y(_14149_));
 AO21x1_ASAP7_75t_SL _22419_ (.A1(_13797_),
    .A2(_13892_),
    .B(_14149_),
    .Y(_14150_));
 NAND2x1_ASAP7_75t_SL _22420_ (.A(_13542_),
    .B(_13818_),
    .Y(_14151_));
 NAND2x1_ASAP7_75t_SL _22421_ (.A(_13560_),
    .B(_13656_),
    .Y(_14152_));
 NOR2x1_ASAP7_75t_SL _22422_ (.A(_13749_),
    .B(_13542_),
    .Y(_14153_));
 NOR2x1_ASAP7_75t_SL _22423_ (.A(_14152_),
    .B(_14153_),
    .Y(_14154_));
 AOI21x1_ASAP7_75t_SL _22424_ (.A1(_14151_),
    .A2(_14154_),
    .B(_13613_),
    .Y(_14155_));
 AO21x1_ASAP7_75t_SL _22425_ (.A1(_14150_),
    .A2(_14155_),
    .B(_13582_),
    .Y(_14156_));
 AOI22x1_ASAP7_75t_SL _22426_ (.A1(_13599_),
    .A2(_13774_),
    .B1(_13790_),
    .B2(_13645_),
    .Y(_14157_));
 AO21x1_ASAP7_75t_SL _22427_ (.A1(_13833_),
    .A2(_13531_),
    .B(_13597_),
    .Y(_14158_));
 NOR2x1_ASAP7_75t_SL _22428_ (.A(_01163_),
    .B(_13531_),
    .Y(_14159_));
 AO21x1_ASAP7_75t_SL _22429_ (.A1(_13531_),
    .A2(_13702_),
    .B(_14159_),
    .Y(_14160_));
 OAI21x1_ASAP7_75t_SL _22430_ (.A1(_14158_),
    .A2(_14160_),
    .B(_13613_),
    .Y(_14161_));
 AOI21x1_ASAP7_75t_SL _22431_ (.A1(_13597_),
    .A2(_14157_),
    .B(_14161_),
    .Y(_14162_));
 NOR2x1_ASAP7_75t_SL _22432_ (.A(_14156_),
    .B(_14162_),
    .Y(_14163_));
 AO21x1_ASAP7_75t_SL _22433_ (.A1(_13542_),
    .A2(_01154_),
    .B(_13597_),
    .Y(_14164_));
 OAI21x1_ASAP7_75t_SL _22434_ (.A1(_14153_),
    .A2(_14164_),
    .B(_13613_),
    .Y(_14165_));
 INVx1_ASAP7_75t_SL _22435_ (.A(_13734_),
    .Y(_14166_));
 AOI21x1_ASAP7_75t_SL _22436_ (.A1(_13537_),
    .A2(_13531_),
    .B(_13560_),
    .Y(_14167_));
 NAND2x1_ASAP7_75t_SL _22437_ (.A(_14167_),
    .B(_13964_),
    .Y(_14168_));
 NOR2x1_ASAP7_75t_SL _22438_ (.A(_14166_),
    .B(_14168_),
    .Y(_14169_));
 OAI21x1_ASAP7_75t_SL _22439_ (.A1(_14165_),
    .A2(_14169_),
    .B(_13582_),
    .Y(_14170_));
 INVx1_ASAP7_75t_SL _22440_ (.A(_13939_),
    .Y(_14171_));
 NAND2x1_ASAP7_75t_SL _22441_ (.A(_13531_),
    .B(_13533_),
    .Y(_14172_));
 NAND2x1_ASAP7_75t_SL _22442_ (.A(_14167_),
    .B(_14172_),
    .Y(_14173_));
 OAI21x1_ASAP7_75t_SL _22443_ (.A1(_14171_),
    .A2(_14173_),
    .B(_13694_),
    .Y(_14174_));
 NAND2x1_ASAP7_75t_SL _22444_ (.A(_13889_),
    .B(_13715_),
    .Y(_14175_));
 NAND3x1_ASAP7_75t_SL _22445_ (.A(_13752_),
    .B(_13531_),
    .C(_13656_),
    .Y(_14176_));
 AOI21x1_ASAP7_75t_SL _22446_ (.A1(_14175_),
    .A2(_14176_),
    .B(_13597_),
    .Y(_14177_));
 NOR2x1_ASAP7_75t_SL _22447_ (.A(_14174_),
    .B(_14177_),
    .Y(_14178_));
 OAI21x1_ASAP7_75t_SL _22448_ (.A1(_14170_),
    .A2(_14178_),
    .B(_13623_),
    .Y(_14179_));
 OAI22x1_ASAP7_75t_SL _22449_ (.A1(_14148_),
    .A2(_14136_),
    .B1(_14163_),
    .B2(_14179_),
    .Y(_00071_));
 XOR2x2_ASAP7_75t_SL _22450_ (.A(_00654_),
    .B(_00647_),
    .Y(_14180_));
 XOR2x1_ASAP7_75t_SL _22451_ (.A(_00648_),
    .Y(_14181_),
    .B(_00680_));
 XOR2x2_ASAP7_75t_SL _22452_ (.A(_14181_),
    .B(_14180_),
    .Y(_14182_));
 XOR2x2_ASAP7_75t_SL _22453_ (.A(_00584_),
    .B(_11386_),
    .Y(_14183_));
 AND2x2_ASAP7_75t_SL _22454_ (.A(_14182_),
    .B(_14183_),
    .Y(_14184_));
 OAI21x1_ASAP7_75t_SL _22455_ (.A1(_14183_),
    .A2(_14182_),
    .B(_00574_),
    .Y(_14185_));
 NAND2x1_ASAP7_75t_R _22456_ (.A(_00459_),
    .B(_10675_),
    .Y(_14186_));
 OAI21x1_ASAP7_75t_SL _22457_ (.A1(_14185_),
    .A2(_14184_),
    .B(_14186_),
    .Y(_14187_));
 XOR2x2_ASAP7_75t_SL _22458_ (.A(_14187_),
    .B(_00878_),
    .Y(_14188_));
 NOR2x1_ASAP7_75t_R _22460_ (.A(_00574_),
    .B(_00460_),
    .Y(_14189_));
 INVx1_ASAP7_75t_R _22461_ (.A(_14189_),
    .Y(_14190_));
 XOR2x2_ASAP7_75t_R _22462_ (.A(_00583_),
    .B(_00622_),
    .Y(_14191_));
 NAND2x1_ASAP7_75t_R _22463_ (.A(_11408_),
    .B(_14191_),
    .Y(_14192_));
 XNOR2x2_ASAP7_75t_R _22464_ (.A(_00583_),
    .B(_00622_),
    .Y(_14193_));
 NAND2x1_ASAP7_75t_R _22465_ (.A(_00679_),
    .B(_14193_),
    .Y(_14194_));
 INVx1_ASAP7_75t_R _22466_ (.A(_14180_),
    .Y(_14195_));
 AOI21x1_ASAP7_75t_R _22467_ (.A1(_14192_),
    .A2(_14194_),
    .B(_14195_),
    .Y(_14196_));
 XOR2x2_ASAP7_75t_R _22468_ (.A(_00622_),
    .B(_00679_),
    .Y(_14197_));
 NAND2x1_ASAP7_75t_R _22469_ (.A(_00583_),
    .B(_14197_),
    .Y(_14198_));
 INVx1_ASAP7_75t_R _22470_ (.A(_00583_),
    .Y(_14199_));
 XNOR2x2_ASAP7_75t_R _22471_ (.A(_00622_),
    .B(_00679_),
    .Y(_14200_));
 NAND2x1_ASAP7_75t_R _22472_ (.A(_14199_),
    .B(_14200_),
    .Y(_14201_));
 AOI21x1_ASAP7_75t_R _22473_ (.A1(_14198_),
    .A2(_14201_),
    .B(_14180_),
    .Y(_14202_));
 OAI21x1_ASAP7_75t_SL _22474_ (.A1(_14196_),
    .A2(_14202_),
    .B(_00574_),
    .Y(_14203_));
 NAND2x1_ASAP7_75t_SL _22475_ (.A(_14190_),
    .B(_14203_),
    .Y(_14204_));
 XNOR2x2_ASAP7_75t_SL _22476_ (.A(_00877_),
    .B(_14204_),
    .Y(_14205_));
 OR2x2_ASAP7_75t_R _22478_ (.A(_00574_),
    .B(_00461_),
    .Y(_14206_));
 INVx1_ASAP7_75t_R _22479_ (.A(_00585_),
    .Y(_14207_));
 NOR2x1_ASAP7_75t_SL _22480_ (.A(_14207_),
    .B(_11441_),
    .Y(_14208_));
 NOR2x1_ASAP7_75t_SL _22481_ (.A(_00585_),
    .B(_11430_),
    .Y(_14209_));
 OAI21x1_ASAP7_75t_SL _22482_ (.A1(_14208_),
    .A2(_14209_),
    .B(_11389_),
    .Y(_14210_));
 INVx1_ASAP7_75t_SL _22483_ (.A(_14210_),
    .Y(_14211_));
 NOR3x1_ASAP7_75t_L _22484_ (.A(_14209_),
    .B(_14208_),
    .C(_11389_),
    .Y(_14212_));
 OAI21x1_ASAP7_75t_SL _22485_ (.A1(_14211_),
    .A2(_14212_),
    .B(_00574_),
    .Y(_14213_));
 INVx1_ASAP7_75t_R _22486_ (.A(_00879_),
    .Y(_14214_));
 AOI21x1_ASAP7_75t_SL _22487_ (.A1(_14206_),
    .A2(_14213_),
    .B(_14214_),
    .Y(_14215_));
 NAND2x1_ASAP7_75t_R _22488_ (.A(_00461_),
    .B(_10675_),
    .Y(_14216_));
 INVx1_ASAP7_75t_R _22489_ (.A(_11389_),
    .Y(_14217_));
 XOR2x2_ASAP7_75t_SL _22490_ (.A(_11441_),
    .B(_14207_),
    .Y(_14218_));
 NAND2x1_ASAP7_75t_SL _22491_ (.A(_14217_),
    .B(_14218_),
    .Y(_14219_));
 NAND3x1_ASAP7_75t_SL _22492_ (.A(_14219_),
    .B(_00574_),
    .C(_14210_),
    .Y(_14220_));
 AOI21x1_ASAP7_75t_SL _22493_ (.A1(_14216_),
    .A2(_14220_),
    .B(_00879_),
    .Y(_14221_));
 NOR2x2_ASAP7_75t_SL _22494_ (.A(_14215_),
    .B(_14221_),
    .Y(_14222_));
 NAND3x1_ASAP7_75t_L _22498_ (.A(_14203_),
    .B(_00877_),
    .C(_14190_),
    .Y(_14225_));
 AO21x1_ASAP7_75t_SL _22499_ (.A1(_14190_),
    .A2(_14203_),
    .B(_00877_),
    .Y(_14226_));
 NAND2x1p5_ASAP7_75t_SL _22500_ (.A(_14226_),
    .B(_14225_),
    .Y(_14227_));
 AOI21x1_ASAP7_75t_SL _22502_ (.A1(_14206_),
    .A2(_14213_),
    .B(_00879_),
    .Y(_14228_));
 AOI21x1_ASAP7_75t_SL _22503_ (.A1(_14216_),
    .A2(_14220_),
    .B(_14214_),
    .Y(_14229_));
 NOR2x2_ASAP7_75t_SL _22504_ (.A(_14228_),
    .B(_14229_),
    .Y(_14230_));
 NAND3x1_ASAP7_75t_R _22507_ (.A(_14213_),
    .B(_00879_),
    .C(_14206_),
    .Y(_14232_));
 INVx1_ASAP7_75t_R _22508_ (.A(_14228_),
    .Y(_14233_));
 INVx4_ASAP7_75t_SL _22510_ (.A(_01168_),
    .Y(_14235_));
 AOI21x1_ASAP7_75t_SL _22511_ (.A1(_14232_),
    .A2(_14233_),
    .B(_14235_),
    .Y(_14236_));
 NOR2x1_ASAP7_75t_SL _22512_ (.A(_14188_),
    .B(_14222_),
    .Y(_14237_));
 NOR2x1_ASAP7_75t_R _22513_ (.A(_00574_),
    .B(_00499_),
    .Y(_14238_));
 XOR2x2_ASAP7_75t_L _22514_ (.A(_00649_),
    .B(_00654_),
    .Y(_14239_));
 XNOR2x2_ASAP7_75t_SL _22515_ (.A(_11455_),
    .B(_14239_),
    .Y(_14240_));
 XNOR2x2_ASAP7_75t_SL _22516_ (.A(_00586_),
    .B(_11454_),
    .Y(_14241_));
 XOR2x2_ASAP7_75t_SL _22517_ (.A(_14240_),
    .B(_14241_),
    .Y(_14242_));
 NOR2x1_ASAP7_75t_SL _22518_ (.A(_10675_),
    .B(_14242_),
    .Y(_14243_));
 INVx1_ASAP7_75t_R _22519_ (.A(_00880_),
    .Y(_14244_));
 OAI21x1_ASAP7_75t_R _22520_ (.A1(_14238_),
    .A2(_14243_),
    .B(_14244_),
    .Y(_14245_));
 NOR2x1_ASAP7_75t_R _22521_ (.A(_14241_),
    .B(_14240_),
    .Y(_14246_));
 AND2x2_ASAP7_75t_SL _22522_ (.A(_14240_),
    .B(_14241_),
    .Y(_14247_));
 OAI21x1_ASAP7_75t_R _22523_ (.A1(_14246_),
    .A2(_14247_),
    .B(_00574_),
    .Y(_14248_));
 INVx1_ASAP7_75t_R _22524_ (.A(_14238_),
    .Y(_14249_));
 NAND3x1_ASAP7_75t_SL _22525_ (.A(_14248_),
    .B(_00880_),
    .C(_14249_),
    .Y(_14250_));
 NAND2x2_ASAP7_75t_SL _22526_ (.A(_14245_),
    .B(_14250_),
    .Y(_14251_));
 OAI21x1_ASAP7_75t_SL _22528_ (.A1(_14237_),
    .A2(_14236_),
    .B(_14251_),
    .Y(_14253_));
 NOR2x1_ASAP7_75t_SL _22529_ (.A(_14227_),
    .B(_14222_),
    .Y(_14254_));
 INVx1_ASAP7_75t_SL _22530_ (.A(_01173_),
    .Y(_14255_));
 NOR2x1_ASAP7_75t_SL _22532_ (.A(_14255_),
    .B(_14230_),
    .Y(_14257_));
 OAI21x1_ASAP7_75t_SL _22533_ (.A1(_14238_),
    .A2(_14243_),
    .B(_00880_),
    .Y(_14258_));
 NAND3x1_ASAP7_75t_SL _22534_ (.A(_14248_),
    .B(_14244_),
    .C(_14249_),
    .Y(_14259_));
 NAND2x1_ASAP7_75t_SL _22535_ (.A(_14258_),
    .B(_14259_),
    .Y(_14260_));
 OAI21x1_ASAP7_75t_SL _22538_ (.A1(_14254_),
    .A2(_14257_),
    .B(_14260_),
    .Y(_14263_));
 AND2x2_ASAP7_75t_R _22539_ (.A(_10675_),
    .B(_00498_),
    .Y(_14264_));
 XOR2x2_ASAP7_75t_R _22540_ (.A(_00587_),
    .B(_00651_),
    .Y(_14265_));
 XOR2x2_ASAP7_75t_SL _22541_ (.A(_11481_),
    .B(_14265_),
    .Y(_14266_));
 XOR2x2_ASAP7_75t_L _22542_ (.A(_00650_),
    .B(_00654_),
    .Y(_14267_));
 INVx1_ASAP7_75t_R _22543_ (.A(_00683_),
    .Y(_14268_));
 XOR2x2_ASAP7_75t_SL _22544_ (.A(_14267_),
    .B(_14268_),
    .Y(_14269_));
 XOR2x2_ASAP7_75t_SL _22545_ (.A(_14266_),
    .B(_14269_),
    .Y(_14270_));
 NOR2x1_ASAP7_75t_R _22546_ (.A(_10675_),
    .B(_14270_),
    .Y(_14271_));
 INVx1_ASAP7_75t_R _22547_ (.A(_00882_),
    .Y(_14272_));
 OAI21x1_ASAP7_75t_R _22548_ (.A1(_14264_),
    .A2(_14271_),
    .B(_14272_),
    .Y(_14273_));
 NOR2x1_ASAP7_75t_R _22549_ (.A(_00574_),
    .B(_00498_),
    .Y(_14274_));
 XNOR2x2_ASAP7_75t_SL _22550_ (.A(_14269_),
    .B(_14266_),
    .Y(_14275_));
 NOR2x1_ASAP7_75t_R _22551_ (.A(_10675_),
    .B(_14275_),
    .Y(_14276_));
 OAI21x1_ASAP7_75t_R _22552_ (.A1(_14274_),
    .A2(_14276_),
    .B(_00882_),
    .Y(_14277_));
 NAND2x2_ASAP7_75t_SL _22553_ (.A(_14273_),
    .B(_14277_),
    .Y(_14278_));
 AOI21x1_ASAP7_75t_SL _22555_ (.A1(_14253_),
    .A2(_14263_),
    .B(_14278_),
    .Y(_14280_));
 AOI21x1_ASAP7_75t_SL _22556_ (.A1(_01171_),
    .A2(_14230_),
    .B(_14251_),
    .Y(_14281_));
 INVx1_ASAP7_75t_SL _22557_ (.A(_14281_),
    .Y(_14282_));
 INVx1_ASAP7_75t_R _22558_ (.A(_01167_),
    .Y(_14283_));
 NOR2x1_ASAP7_75t_SL _22559_ (.A(_14283_),
    .B(_14230_),
    .Y(_14284_));
 NOR2x1_ASAP7_75t_SL _22560_ (.A(_01169_),
    .B(_14222_),
    .Y(_14285_));
 OAI21x1_ASAP7_75t_SL _22563_ (.A1(_14284_),
    .A2(_14285_),
    .B(_14251_),
    .Y(_14288_));
 INVx3_ASAP7_75t_SL _22564_ (.A(_14278_),
    .Y(_14289_));
 AOI21x1_ASAP7_75t_SL _22567_ (.A1(_14282_),
    .A2(_14288_),
    .B(_14289_),
    .Y(_14292_));
 XNOR2x2_ASAP7_75t_R _22568_ (.A(_00588_),
    .B(_00619_),
    .Y(_14293_));
 XOR2x2_ASAP7_75t_SL _22569_ (.A(_00651_),
    .B(_00652_),
    .Y(_14294_));
 INVx1_ASAP7_75t_R _22570_ (.A(_00684_),
    .Y(_14295_));
 XOR2x2_ASAP7_75t_R _22571_ (.A(_14294_),
    .B(_14295_),
    .Y(_14296_));
 XNOR2x2_ASAP7_75t_L _22572_ (.A(_14293_),
    .B(_14296_),
    .Y(_14297_));
 NOR2x1_ASAP7_75t_R _22573_ (.A(_00574_),
    .B(_00497_),
    .Y(_14298_));
 AOI21x1_ASAP7_75t_R _22574_ (.A1(_00574_),
    .A2(_14297_),
    .B(_14298_),
    .Y(_14299_));
 XNOR2x2_ASAP7_75t_SL _22575_ (.A(_00883_),
    .B(_14299_),
    .Y(_14300_));
 INVx1_ASAP7_75t_SL _22576_ (.A(_14300_),
    .Y(_14301_));
 OAI21x1_ASAP7_75t_SL _22578_ (.A1(_14280_),
    .A2(_14292_),
    .B(_14301_),
    .Y(_14303_));
 INVx1_ASAP7_75t_SL _22579_ (.A(_01171_),
    .Y(_14304_));
 OAI21x1_ASAP7_75t_SL _22580_ (.A1(_14228_),
    .A2(_14229_),
    .B(_14304_),
    .Y(_14305_));
 OAI21x1_ASAP7_75t_SL _22581_ (.A1(_14260_),
    .A2(_14305_),
    .B(_14289_),
    .Y(_14306_));
 INVx1_ASAP7_75t_SL _22582_ (.A(_14306_),
    .Y(_14307_));
 XNOR2x2_ASAP7_75t_SL _22583_ (.A(_14187_),
    .B(_00878_),
    .Y(_14308_));
 OAI21x1_ASAP7_75t_SL _22584_ (.A1(_14308_),
    .A2(_14227_),
    .B(_14230_),
    .Y(_14309_));
 NAND2x2_ASAP7_75t_SL _22585_ (.A(_14205_),
    .B(_14222_),
    .Y(_14310_));
 AO21x1_ASAP7_75t_SL _22586_ (.A1(_14309_),
    .A2(_14310_),
    .B(_14251_),
    .Y(_14311_));
 NAND2x1_ASAP7_75t_SL _22587_ (.A(_14307_),
    .B(_14311_),
    .Y(_14312_));
 OA21x2_ASAP7_75t_SL _22589_ (.A1(_14260_),
    .A2(_14305_),
    .B(_14278_),
    .Y(_14314_));
 INVx1_ASAP7_75t_SL _22590_ (.A(_01174_),
    .Y(_14315_));
 OAI21x1_ASAP7_75t_R _22591_ (.A1(_14215_),
    .A2(_14221_),
    .B(_14315_),
    .Y(_14316_));
 NOR2x1_ASAP7_75t_R _22592_ (.A(_14316_),
    .B(_14260_),
    .Y(_14317_));
 OAI21x1_ASAP7_75t_SL _22593_ (.A1(_14215_),
    .A2(_14221_),
    .B(_01168_),
    .Y(_14318_));
 NAND2x1p5_ASAP7_75t_SL _22594_ (.A(_14260_),
    .B(_14318_),
    .Y(_14319_));
 INVx3_ASAP7_75t_SL _22595_ (.A(_14319_),
    .Y(_14320_));
 NOR2x1_ASAP7_75t_SL _22596_ (.A(_14317_),
    .B(_14320_),
    .Y(_14321_));
 AOI21x1_ASAP7_75t_SL _22598_ (.A1(_14321_),
    .A2(_14314_),
    .B(_14301_),
    .Y(_14323_));
 NAND2x1_ASAP7_75t_SL _22599_ (.A(_14312_),
    .B(_14323_),
    .Y(_14324_));
 XOR2x2_ASAP7_75t_R _22600_ (.A(_00653_),
    .B(_00685_),
    .Y(_14325_));
 XOR2x2_ASAP7_75t_R _22601_ (.A(_11543_),
    .B(_00589_),
    .Y(_14326_));
 XNOR2x2_ASAP7_75t_R _22602_ (.A(_14325_),
    .B(_14326_),
    .Y(_14327_));
 NOR2x1_ASAP7_75t_R _22604_ (.A(_00574_),
    .B(_00496_),
    .Y(_14329_));
 AO21x1_ASAP7_75t_SL _22605_ (.A1(_14327_),
    .A2(_00574_),
    .B(_14329_),
    .Y(_14330_));
 XOR2x2_ASAP7_75t_SL _22606_ (.A(_14330_),
    .B(_00884_),
    .Y(_14331_));
 INVx2_ASAP7_75t_SL _22607_ (.A(_14331_),
    .Y(_14332_));
 NAND3x1_ASAP7_75t_SL _22609_ (.A(_14324_),
    .B(_14303_),
    .C(_14332_),
    .Y(_14334_));
 NAND2x1_ASAP7_75t_SL _22610_ (.A(_14188_),
    .B(_14227_),
    .Y(_14335_));
 NAND2x1_ASAP7_75t_SL _22611_ (.A(_14230_),
    .B(_14335_),
    .Y(_14336_));
 AOI21x1_ASAP7_75t_SL _22612_ (.A1(_14305_),
    .A2(_14336_),
    .B(_14260_),
    .Y(_14337_));
 NOR2x1_ASAP7_75t_SL _22613_ (.A(_01169_),
    .B(_14230_),
    .Y(_14338_));
 AOI21x1_ASAP7_75t_SL _22614_ (.A1(_14251_),
    .A2(_14338_),
    .B(_14278_),
    .Y(_14339_));
 NAND2x2_ASAP7_75t_SL _22616_ (.A(_01167_),
    .B(_14230_),
    .Y(_14341_));
 AO21x1_ASAP7_75t_SL _22618_ (.A1(_14310_),
    .A2(_14341_),
    .B(_14251_),
    .Y(_14343_));
 NAND2x1_ASAP7_75t_SL _22619_ (.A(_14339_),
    .B(_14343_),
    .Y(_14344_));
 AO21x1_ASAP7_75t_SL _22620_ (.A1(_14259_),
    .A2(_14258_),
    .B(_01181_),
    .Y(_14345_));
 NAND2x1p5_ASAP7_75t_SL _22621_ (.A(_14235_),
    .B(_14222_),
    .Y(_14346_));
 OA21x2_ASAP7_75t_SL _22624_ (.A1(_14346_),
    .A2(_14260_),
    .B(_14278_),
    .Y(_14349_));
 AOI21x1_ASAP7_75t_SL _22626_ (.A1(_14345_),
    .A2(_14349_),
    .B(_14301_),
    .Y(_14351_));
 OAI21x1_ASAP7_75t_SL _22627_ (.A1(_14337_),
    .A2(_14344_),
    .B(_14351_),
    .Y(_14352_));
 INVx1_ASAP7_75t_SL _22628_ (.A(_01169_),
    .Y(_14353_));
 NAND2x1_ASAP7_75t_SL _22629_ (.A(_14353_),
    .B(_14230_),
    .Y(_14354_));
 OA21x2_ASAP7_75t_SL _22631_ (.A1(_14354_),
    .A2(_14260_),
    .B(_14289_),
    .Y(_14356_));
 NOR2x2_ASAP7_75t_SL _22632_ (.A(_14308_),
    .B(_14205_),
    .Y(_14357_));
 NAND2x1_ASAP7_75t_SL _22633_ (.A(_14230_),
    .B(_14357_),
    .Y(_14358_));
 NOR2x1_ASAP7_75t_L _22634_ (.A(_14315_),
    .B(_14230_),
    .Y(_14359_));
 NOR2x1_ASAP7_75t_SL _22635_ (.A(_14251_),
    .B(_14359_),
    .Y(_14360_));
 NAND2x1_ASAP7_75t_SL _22636_ (.A(_14358_),
    .B(_14360_),
    .Y(_14361_));
 NAND2x1_ASAP7_75t_SL _22637_ (.A(_14356_),
    .B(_14361_),
    .Y(_14362_));
 AOI21x1_ASAP7_75t_R _22638_ (.A1(_14232_),
    .A2(_14233_),
    .B(_01173_),
    .Y(_14363_));
 NOR2x1_ASAP7_75t_SL _22639_ (.A(_14260_),
    .B(_14363_),
    .Y(_14364_));
 NAND2x1_ASAP7_75t_SL _22640_ (.A(_14364_),
    .B(_14358_),
    .Y(_14365_));
 OA21x2_ASAP7_75t_SL _22641_ (.A1(_14354_),
    .A2(_14251_),
    .B(_14278_),
    .Y(_14366_));
 AOI21x1_ASAP7_75t_SL _22643_ (.A1(_14365_),
    .A2(_14366_),
    .B(_14300_),
    .Y(_14368_));
 AOI21x1_ASAP7_75t_SL _22644_ (.A1(_14362_),
    .A2(_14368_),
    .B(_14332_),
    .Y(_14369_));
 XNOR2x2_ASAP7_75t_R _22645_ (.A(_00590_),
    .B(_00621_),
    .Y(_14370_));
 XOR2x2_ASAP7_75t_L _22646_ (.A(_00653_),
    .B(_00654_),
    .Y(_14371_));
 XOR2x2_ASAP7_75t_R _22647_ (.A(_14371_),
    .B(_11589_),
    .Y(_14372_));
 XNOR2x2_ASAP7_75t_R _22648_ (.A(_14370_),
    .B(_14372_),
    .Y(_14373_));
 NOR2x1_ASAP7_75t_R _22649_ (.A(_00574_),
    .B(_00495_),
    .Y(_14374_));
 AO21x1_ASAP7_75t_SL _22650_ (.A1(_14373_),
    .A2(_00574_),
    .B(_14374_),
    .Y(_14375_));
 XOR2x2_ASAP7_75t_SL _22651_ (.A(_14375_),
    .B(_00885_),
    .Y(_14376_));
 AOI21x1_ASAP7_75t_SL _22652_ (.A1(_14352_),
    .A2(_14369_),
    .B(_14376_),
    .Y(_14377_));
 NAND2x1_ASAP7_75t_SL _22653_ (.A(_14334_),
    .B(_14377_),
    .Y(_14378_));
 NAND2x1_ASAP7_75t_SL _22654_ (.A(_01167_),
    .B(_14222_),
    .Y(_14379_));
 OAI21x1_ASAP7_75t_SL _22655_ (.A1(_14215_),
    .A2(_14221_),
    .B(_14235_),
    .Y(_14380_));
 AO21x1_ASAP7_75t_SL _22657_ (.A1(_14380_),
    .A2(_14379_),
    .B(_14251_),
    .Y(_14382_));
 NAND2x1_ASAP7_75t_SL _22658_ (.A(_01173_),
    .B(_14222_),
    .Y(_14383_));
 AO21x1_ASAP7_75t_SL _22659_ (.A1(_14341_),
    .A2(_14383_),
    .B(_14260_),
    .Y(_14384_));
 AOI21x1_ASAP7_75t_SL _22660_ (.A1(_14384_),
    .A2(_14382_),
    .B(_14278_),
    .Y(_14385_));
 NOR2x1p5_ASAP7_75t_SL _22661_ (.A(_14236_),
    .B(_14251_),
    .Y(_14386_));
 NOR2x1p5_ASAP7_75t_SL _22662_ (.A(_14386_),
    .B(_14289_),
    .Y(_14387_));
 INVx2_ASAP7_75t_SL _22663_ (.A(_14387_),
    .Y(_14388_));
 NAND2x2_ASAP7_75t_SL _22664_ (.A(_14308_),
    .B(_14222_),
    .Y(_14389_));
 INVx1_ASAP7_75t_SL _22665_ (.A(_14389_),
    .Y(_14390_));
 NOR2x1p5_ASAP7_75t_SL _22666_ (.A(_14260_),
    .B(_14318_),
    .Y(_14391_));
 AO21x1_ASAP7_75t_SL _22667_ (.A1(_14390_),
    .A2(_14251_),
    .B(_14391_),
    .Y(_14392_));
 OAI21x1_ASAP7_75t_SL _22668_ (.A1(_14388_),
    .A2(_14392_),
    .B(_14300_),
    .Y(_14393_));
 NOR2x1_ASAP7_75t_SL _22669_ (.A(_14393_),
    .B(_14385_),
    .Y(_14394_));
 AO21x1_ASAP7_75t_SL _22670_ (.A1(_14310_),
    .A2(_14335_),
    .B(_14260_),
    .Y(_14395_));
 NOR2x1_ASAP7_75t_SL _22671_ (.A(_14251_),
    .B(_14357_),
    .Y(_14396_));
 AOI21x1_ASAP7_75t_SL _22673_ (.A1(_14310_),
    .A2(_14396_),
    .B(_14289_),
    .Y(_14398_));
 NAND2x1_ASAP7_75t_SL _22674_ (.A(_14395_),
    .B(_14398_),
    .Y(_14399_));
 NOR2x2_ASAP7_75t_SL _22675_ (.A(_14308_),
    .B(_14227_),
    .Y(_14400_));
 NAND2x1p5_ASAP7_75t_SL _22676_ (.A(_14251_),
    .B(_14318_),
    .Y(_14401_));
 AO21x1_ASAP7_75t_SL _22677_ (.A1(_14222_),
    .A2(_14400_),
    .B(_14401_),
    .Y(_14402_));
 NAND2x1_ASAP7_75t_SL _22678_ (.A(_01173_),
    .B(_14230_),
    .Y(_14403_));
 NAND2x1_ASAP7_75t_SL _22679_ (.A(_14379_),
    .B(_14403_),
    .Y(_14404_));
 AOI21x1_ASAP7_75t_SL _22681_ (.A1(_14260_),
    .A2(_14404_),
    .B(_14278_),
    .Y(_14406_));
 NAND2x1_ASAP7_75t_SL _22682_ (.A(_14402_),
    .B(_14406_),
    .Y(_14407_));
 AOI21x1_ASAP7_75t_SL _22684_ (.A1(_14399_),
    .A2(_14407_),
    .B(_14300_),
    .Y(_14409_));
 OAI21x1_ASAP7_75t_SL _22686_ (.A1(_14409_),
    .A2(_14394_),
    .B(_14331_),
    .Y(_14411_));
 OAI21x1_ASAP7_75t_SL _22687_ (.A1(_14188_),
    .A2(_14230_),
    .B(_14227_),
    .Y(_14412_));
 NAND2x1_ASAP7_75t_SL _22688_ (.A(_14251_),
    .B(_14412_),
    .Y(_14413_));
 NAND2x1_ASAP7_75t_SL _22689_ (.A(_01176_),
    .B(_14222_),
    .Y(_14414_));
 AOI21x1_ASAP7_75t_SL _22691_ (.A1(_14414_),
    .A2(_14320_),
    .B(_14289_),
    .Y(_14416_));
 NAND2x1_ASAP7_75t_SL _22692_ (.A(_14416_),
    .B(_14413_),
    .Y(_14417_));
 NAND2x1_ASAP7_75t_SL _22694_ (.A(_14227_),
    .B(_14222_),
    .Y(_14419_));
 AOI21x1_ASAP7_75t_SL _22695_ (.A1(_14251_),
    .A2(_14419_),
    .B(_14278_),
    .Y(_14420_));
 NAND2x1_ASAP7_75t_SL _22696_ (.A(_14222_),
    .B(_14357_),
    .Y(_14421_));
 NAND2x1_ASAP7_75t_SL _22697_ (.A(_14421_),
    .B(_14281_),
    .Y(_14422_));
 AOI21x1_ASAP7_75t_SL _22698_ (.A1(_14420_),
    .A2(_14422_),
    .B(_14300_),
    .Y(_14423_));
 AOI21x1_ASAP7_75t_SL _22699_ (.A1(_14423_),
    .A2(_14417_),
    .B(_14331_),
    .Y(_14424_));
 INVx1_ASAP7_75t_SL _22700_ (.A(_01176_),
    .Y(_14425_));
 NAND2x1_ASAP7_75t_SL _22701_ (.A(_14425_),
    .B(_14230_),
    .Y(_14426_));
 AO21x1_ASAP7_75t_SL _22702_ (.A1(_14310_),
    .A2(_14426_),
    .B(_14251_),
    .Y(_14427_));
 NOR2x1_ASAP7_75t_SL _22703_ (.A(_14260_),
    .B(_14237_),
    .Y(_14428_));
 AOI21x1_ASAP7_75t_SL _22704_ (.A1(_14421_),
    .A2(_14428_),
    .B(_14289_),
    .Y(_14429_));
 AOI21x1_ASAP7_75t_SL _22705_ (.A1(_14427_),
    .A2(_14429_),
    .B(_14301_),
    .Y(_14430_));
 AO21x1_ASAP7_75t_SL _22706_ (.A1(_14389_),
    .A2(_14354_),
    .B(_14260_),
    .Y(_14431_));
 NAND3x1_ASAP7_75t_SL _22707_ (.A(_14311_),
    .B(_14289_),
    .C(_14431_),
    .Y(_14432_));
 NAND2x1_ASAP7_75t_SL _22708_ (.A(_14430_),
    .B(_14432_),
    .Y(_14433_));
 INVx1_ASAP7_75t_SL _22709_ (.A(_14376_),
    .Y(_14434_));
 AOI21x1_ASAP7_75t_SL _22710_ (.A1(_14433_),
    .A2(_14424_),
    .B(_14434_),
    .Y(_14435_));
 NAND2x1_ASAP7_75t_SL _22711_ (.A(_14411_),
    .B(_14435_),
    .Y(_14436_));
 NAND2x1_ASAP7_75t_SL _22712_ (.A(_14378_),
    .B(_14436_),
    .Y(_00072_));
 AOI21x1_ASAP7_75t_SL _22714_ (.A1(_14341_),
    .A2(_14346_),
    .B(_14251_),
    .Y(_14438_));
 AOI21x1_ASAP7_75t_SL _22716_ (.A1(_14310_),
    .A2(_14354_),
    .B(_14260_),
    .Y(_14440_));
 OAI21x1_ASAP7_75t_SL _22718_ (.A1(_14438_),
    .A2(_14440_),
    .B(_14278_),
    .Y(_14442_));
 NAND2x1_ASAP7_75t_SL _22719_ (.A(_14188_),
    .B(_14222_),
    .Y(_14443_));
 NAND2x1_ASAP7_75t_SL _22720_ (.A(_14304_),
    .B(_14230_),
    .Y(_14444_));
 AOI21x1_ASAP7_75t_SL _22721_ (.A1(_14443_),
    .A2(_14444_),
    .B(_14251_),
    .Y(_14445_));
 NOR2x1_ASAP7_75t_SL _22722_ (.A(_01167_),
    .B(_14230_),
    .Y(_14446_));
 NAND2x2_ASAP7_75t_SL _22724_ (.A(_14205_),
    .B(_14230_),
    .Y(_14448_));
 NAND2x1_ASAP7_75t_SL _22725_ (.A(_14251_),
    .B(_14448_),
    .Y(_14449_));
 NOR2x1_ASAP7_75t_SL _22726_ (.A(_14446_),
    .B(_14449_),
    .Y(_14450_));
 OAI21x1_ASAP7_75t_SL _22728_ (.A1(_14445_),
    .A2(_14450_),
    .B(_14289_),
    .Y(_14452_));
 AOI21x1_ASAP7_75t_SL _22730_ (.A1(_14442_),
    .A2(_14452_),
    .B(_14300_),
    .Y(_14454_));
 NAND2x1_ASAP7_75t_R _22731_ (.A(_14188_),
    .B(_14205_),
    .Y(_14455_));
 NAND2x1_ASAP7_75t_SL _22732_ (.A(_14222_),
    .B(_14455_),
    .Y(_14456_));
 AOI21x1_ASAP7_75t_SL _22733_ (.A1(_14318_),
    .A2(_14456_),
    .B(_14251_),
    .Y(_14457_));
 NOR2x1_ASAP7_75t_SL _22734_ (.A(_14353_),
    .B(_14230_),
    .Y(_14458_));
 NAND2x2_ASAP7_75t_SL _22735_ (.A(_01176_),
    .B(_14230_),
    .Y(_14459_));
 NAND2x1_ASAP7_75t_SL _22736_ (.A(_14251_),
    .B(_14459_),
    .Y(_14460_));
 OAI21x1_ASAP7_75t_SL _22737_ (.A1(_14458_),
    .A2(_14460_),
    .B(_14278_),
    .Y(_14461_));
 NOR2x1_ASAP7_75t_SL _22738_ (.A(_14457_),
    .B(_14461_),
    .Y(_14462_));
 AO21x1_ASAP7_75t_SL _22739_ (.A1(_14260_),
    .A2(_14318_),
    .B(_14278_),
    .Y(_14463_));
 NOR2x1_ASAP7_75t_SL _22740_ (.A(_14222_),
    .B(_14455_),
    .Y(_14464_));
 NAND2x1_ASAP7_75t_SL _22741_ (.A(_14251_),
    .B(_14419_),
    .Y(_14465_));
 NOR2x1_ASAP7_75t_SL _22742_ (.A(_14464_),
    .B(_14465_),
    .Y(_14466_));
 OAI21x1_ASAP7_75t_SL _22743_ (.A1(_14463_),
    .A2(_14466_),
    .B(_14300_),
    .Y(_14467_));
 OAI21x1_ASAP7_75t_SL _22744_ (.A1(_14462_),
    .A2(_14467_),
    .B(_14332_),
    .Y(_14468_));
 OAI21x1_ASAP7_75t_SL _22745_ (.A1(_14454_),
    .A2(_14468_),
    .B(_14376_),
    .Y(_14469_));
 NAND2x1_ASAP7_75t_SL _22746_ (.A(_01183_),
    .B(_14300_),
    .Y(_14470_));
 NAND2x1_ASAP7_75t_R _22747_ (.A(_14230_),
    .B(_14400_),
    .Y(_14471_));
 AOI21x1_ASAP7_75t_SL _22748_ (.A1(_14364_),
    .A2(_14471_),
    .B(_14278_),
    .Y(_14472_));
 OAI21x1_ASAP7_75t_SL _22749_ (.A1(_14251_),
    .A2(_14470_),
    .B(_14472_),
    .Y(_14473_));
 NOR2x1_ASAP7_75t_R _22750_ (.A(_14205_),
    .B(_14222_),
    .Y(_14474_));
 OAI21x1_ASAP7_75t_SL _22751_ (.A1(_01167_),
    .A2(_14230_),
    .B(_14251_),
    .Y(_14475_));
 OAI21x1_ASAP7_75t_SL _22752_ (.A1(_14474_),
    .A2(_14475_),
    .B(_14301_),
    .Y(_14476_));
 NAND2x1_ASAP7_75t_SL _22753_ (.A(_14222_),
    .B(_14335_),
    .Y(_14477_));
 AOI21x1_ASAP7_75t_SL _22754_ (.A1(_14309_),
    .A2(_14477_),
    .B(_14251_),
    .Y(_14478_));
 NOR2x1_ASAP7_75t_SL _22755_ (.A(_14476_),
    .B(_14478_),
    .Y(_14479_));
 NOR2x1_ASAP7_75t_SL _22757_ (.A(_14308_),
    .B(_14230_),
    .Y(_14480_));
 OAI21x1_ASAP7_75t_SL _22758_ (.A1(_14480_),
    .A2(_14449_),
    .B(_14300_),
    .Y(_14481_));
 NOR2x1_ASAP7_75t_SL _22759_ (.A(_14445_),
    .B(_14481_),
    .Y(_14482_));
 OAI21x1_ASAP7_75t_SL _22760_ (.A1(_14479_),
    .A2(_14482_),
    .B(_14278_),
    .Y(_14483_));
 AOI21x1_ASAP7_75t_SL _22761_ (.A1(_14473_),
    .A2(_14483_),
    .B(_14332_),
    .Y(_14484_));
 INVx1_ASAP7_75t_SL _22762_ (.A(_14309_),
    .Y(_14485_));
 NAND2x1_ASAP7_75t_SL _22763_ (.A(_14251_),
    .B(_14485_),
    .Y(_14486_));
 OAI21x1_ASAP7_75t_R _22764_ (.A1(_14228_),
    .A2(_14229_),
    .B(_14425_),
    .Y(_14487_));
 NAND2x1_ASAP7_75t_SL _22765_ (.A(_14188_),
    .B(_14230_),
    .Y(_14488_));
 NAND2x1_ASAP7_75t_R _22766_ (.A(_14487_),
    .B(_14488_),
    .Y(_14489_));
 AOI21x1_ASAP7_75t_SL _22767_ (.A1(_14260_),
    .A2(_14489_),
    .B(_14289_),
    .Y(_14490_));
 OAI21x1_ASAP7_75t_SL _22769_ (.A1(_14260_),
    .A2(_14444_),
    .B(_14289_),
    .Y(_14492_));
 OAI21x1_ASAP7_75t_SL _22770_ (.A1(_14492_),
    .A2(_14457_),
    .B(_14301_),
    .Y(_14493_));
 AOI21x1_ASAP7_75t_SL _22771_ (.A1(_14486_),
    .A2(_14490_),
    .B(_14493_),
    .Y(_14494_));
 NAND2x1p5_ASAP7_75t_SL _22772_ (.A(_14305_),
    .B(_14320_),
    .Y(_14495_));
 NAND3x1_ASAP7_75t_SL _22773_ (.A(_14310_),
    .B(_14341_),
    .C(_14251_),
    .Y(_14496_));
 AOI21x1_ASAP7_75t_SL _22774_ (.A1(_14496_),
    .A2(_14495_),
    .B(_14289_),
    .Y(_14497_));
 NAND2x1_ASAP7_75t_SL _22776_ (.A(_14308_),
    .B(_14205_),
    .Y(_14499_));
 AND3x1_ASAP7_75t_SL _22777_ (.A(_14419_),
    .B(_14260_),
    .C(_14499_),
    .Y(_14500_));
 NAND2x1_ASAP7_75t_SL _22778_ (.A(_14251_),
    .B(_14346_),
    .Y(_14501_));
 OAI21x1_ASAP7_75t_SL _22779_ (.A1(_14474_),
    .A2(_14501_),
    .B(_14289_),
    .Y(_14502_));
 OAI21x1_ASAP7_75t_SL _22780_ (.A1(_14500_),
    .A2(_14502_),
    .B(_14300_),
    .Y(_14503_));
 OAI21x1_ASAP7_75t_SL _22781_ (.A1(_14503_),
    .A2(_14497_),
    .B(_14332_),
    .Y(_14504_));
 NOR2x1_ASAP7_75t_SL _22782_ (.A(_14494_),
    .B(_14504_),
    .Y(_14505_));
 AOI21x1_ASAP7_75t_R _22783_ (.A1(_14499_),
    .A2(_14443_),
    .B(_14260_),
    .Y(_14506_));
 NAND2x1_ASAP7_75t_SL _22784_ (.A(_14222_),
    .B(_14260_),
    .Y(_14507_));
 NOR2x1_ASAP7_75t_SL _22785_ (.A(_14357_),
    .B(_14507_),
    .Y(_14508_));
 OAI21x1_ASAP7_75t_SL _22786_ (.A1(_14506_),
    .A2(_14508_),
    .B(_14289_),
    .Y(_14509_));
 AOI21x1_ASAP7_75t_SL _22787_ (.A1(_14310_),
    .A2(_14380_),
    .B(_14251_),
    .Y(_14510_));
 AOI21x1_ASAP7_75t_SL _22788_ (.A1(_14419_),
    .A2(_14444_),
    .B(_14260_),
    .Y(_14511_));
 OAI21x1_ASAP7_75t_SL _22789_ (.A1(_14510_),
    .A2(_14511_),
    .B(_14278_),
    .Y(_14512_));
 AOI21x1_ASAP7_75t_SL _22790_ (.A1(_14512_),
    .A2(_14509_),
    .B(_14300_),
    .Y(_14513_));
 NAND2x1_ASAP7_75t_SL _22791_ (.A(_14308_),
    .B(_14230_),
    .Y(_14514_));
 OAI21x1_ASAP7_75t_SL _22792_ (.A1(_14260_),
    .A2(_14305_),
    .B(_14514_),
    .Y(_14515_));
 AOI21x1_ASAP7_75t_SL _22793_ (.A1(_14260_),
    .A2(_14443_),
    .B(_14289_),
    .Y(_14516_));
 INVx1_ASAP7_75t_SL _22794_ (.A(_14516_),
    .Y(_14517_));
 OAI21x1_ASAP7_75t_SL _22795_ (.A1(_14515_),
    .A2(_14517_),
    .B(_14300_),
    .Y(_14518_));
 NOR2x1_ASAP7_75t_R _22796_ (.A(_14425_),
    .B(_14222_),
    .Y(_14519_));
 OAI21x1_ASAP7_75t_SL _22797_ (.A1(_14228_),
    .A2(_14229_),
    .B(_01168_),
    .Y(_14520_));
 NAND2x1_ASAP7_75t_L _22798_ (.A(_14520_),
    .B(_14260_),
    .Y(_14521_));
 OAI21x1_ASAP7_75t_SL _22799_ (.A1(_14519_),
    .A2(_14521_),
    .B(_14289_),
    .Y(_14522_));
 NOR2x1_ASAP7_75t_SL _22800_ (.A(_14522_),
    .B(_14337_),
    .Y(_14523_));
 OAI21x1_ASAP7_75t_SL _22801_ (.A1(_14518_),
    .A2(_14523_),
    .B(_14331_),
    .Y(_14524_));
 OAI21x1_ASAP7_75t_SL _22802_ (.A1(_14513_),
    .A2(_14524_),
    .B(_14434_),
    .Y(_14525_));
 OAI22x1_ASAP7_75t_SL _22803_ (.A1(_14469_),
    .A2(_14484_),
    .B1(_14505_),
    .B2(_14525_),
    .Y(_00073_));
 AO21x1_ASAP7_75t_SL _22804_ (.A1(_14488_),
    .A2(_14305_),
    .B(_14251_),
    .Y(_14526_));
 NOR2x1_ASAP7_75t_SL _22805_ (.A(_14317_),
    .B(_14306_),
    .Y(_14527_));
 NAND2x1_ASAP7_75t_SL _22806_ (.A(_14526_),
    .B(_14527_),
    .Y(_14528_));
 NOR2x1_ASAP7_75t_SL _22807_ (.A(_14289_),
    .B(_14317_),
    .Y(_14529_));
 NAND2x1_ASAP7_75t_SL _22808_ (.A(_14305_),
    .B(_14260_),
    .Y(_14530_));
 NAND2x1_ASAP7_75t_SL _22809_ (.A(_14487_),
    .B(_14251_),
    .Y(_14531_));
 OAI21x1_ASAP7_75t_SL _22810_ (.A1(_14254_),
    .A2(_14530_),
    .B(_14531_),
    .Y(_14532_));
 AOI21x1_ASAP7_75t_SL _22811_ (.A1(_14529_),
    .A2(_14532_),
    .B(_14301_),
    .Y(_14533_));
 NAND2x1_ASAP7_75t_SL _22812_ (.A(_14528_),
    .B(_14533_),
    .Y(_14534_));
 NAND2x1_ASAP7_75t_SL _22813_ (.A(_14316_),
    .B(_14260_),
    .Y(_14535_));
 NOR2x1_ASAP7_75t_SL _22814_ (.A(_14390_),
    .B(_14535_),
    .Y(_14536_));
 OAI21x1_ASAP7_75t_SL _22815_ (.A1(_14254_),
    .A2(_14531_),
    .B(_14278_),
    .Y(_14537_));
 NOR2x1_ASAP7_75t_SL _22816_ (.A(_14536_),
    .B(_14537_),
    .Y(_14538_));
 AO21x1_ASAP7_75t_SL _22817_ (.A1(_14520_),
    .A2(_14380_),
    .B(_14251_),
    .Y(_14539_));
 NOR2x1_ASAP7_75t_R _22818_ (.A(_01174_),
    .B(_14230_),
    .Y(_14540_));
 OAI21x1_ASAP7_75t_SL _22819_ (.A1(_14254_),
    .A2(_14540_),
    .B(_14251_),
    .Y(_14541_));
 AOI21x1_ASAP7_75t_SL _22821_ (.A1(_14539_),
    .A2(_14541_),
    .B(_14278_),
    .Y(_14543_));
 OAI21x1_ASAP7_75t_SL _22822_ (.A1(_14543_),
    .A2(_14538_),
    .B(_14301_),
    .Y(_14544_));
 AOI21x1_ASAP7_75t_SL _22823_ (.A1(_14544_),
    .A2(_14534_),
    .B(_14331_),
    .Y(_14545_));
 OAI21x1_ASAP7_75t_SL _22824_ (.A1(_01169_),
    .A2(_14230_),
    .B(_14260_),
    .Y(_14546_));
 NOR2x1_ASAP7_75t_SL _22825_ (.A(_14254_),
    .B(_14546_),
    .Y(_14547_));
 NAND2x1p5_ASAP7_75t_SL _22826_ (.A(_14251_),
    .B(_14380_),
    .Y(_14548_));
 OAI21x1_ASAP7_75t_SL _22827_ (.A1(_14548_),
    .A2(_14390_),
    .B(_14278_),
    .Y(_14549_));
 OAI21x1_ASAP7_75t_SL _22828_ (.A1(_14549_),
    .A2(_14547_),
    .B(_14301_),
    .Y(_14550_));
 OAI21x1_ASAP7_75t_SL _22829_ (.A1(_14230_),
    .A2(_14335_),
    .B(_14251_),
    .Y(_14551_));
 INVx1_ASAP7_75t_SL _22830_ (.A(_14426_),
    .Y(_14552_));
 AOI21x1_ASAP7_75t_SL _22831_ (.A1(_14188_),
    .A2(_14205_),
    .B(_14230_),
    .Y(_14553_));
 OAI21x1_ASAP7_75t_SL _22832_ (.A1(_14552_),
    .A2(_14553_),
    .B(_14260_),
    .Y(_14554_));
 AOI21x1_ASAP7_75t_SL _22833_ (.A1(_14551_),
    .A2(_14554_),
    .B(_14278_),
    .Y(_14555_));
 OAI21x1_ASAP7_75t_SL _22834_ (.A1(_14550_),
    .A2(_14555_),
    .B(_14331_),
    .Y(_14556_));
 NOR3x1_ASAP7_75t_SL _22835_ (.A(_14530_),
    .B(_14254_),
    .C(_14237_),
    .Y(_14557_));
 NAND2x1_ASAP7_75t_SL _22836_ (.A(_14289_),
    .B(_14253_),
    .Y(_14558_));
 NOR2x1_ASAP7_75t_SL _22837_ (.A(_14557_),
    .B(_14558_),
    .Y(_14559_));
 AOI21x1_ASAP7_75t_SL _22838_ (.A1(_14487_),
    .A2(_14444_),
    .B(_14260_),
    .Y(_14560_));
 AOI21x1_ASAP7_75t_R _22839_ (.A1(_14205_),
    .A2(_14222_),
    .B(_14308_),
    .Y(_14561_));
 NOR2x1_ASAP7_75t_SL _22840_ (.A(_14251_),
    .B(_14561_),
    .Y(_14562_));
 NOR2x1_ASAP7_75t_SL _22841_ (.A(_14560_),
    .B(_14562_),
    .Y(_14563_));
 OAI21x1_ASAP7_75t_SL _22842_ (.A1(_14289_),
    .A2(_14563_),
    .B(_14300_),
    .Y(_14564_));
 NOR2x1_ASAP7_75t_SL _22843_ (.A(_14559_),
    .B(_14564_),
    .Y(_14565_));
 NOR2x1_ASAP7_75t_SL _22844_ (.A(_14556_),
    .B(_14565_),
    .Y(_14566_));
 OAI21x1_ASAP7_75t_SL _22845_ (.A1(_14566_),
    .A2(_14545_),
    .B(_14376_),
    .Y(_14567_));
 NAND2x1_ASAP7_75t_SL _22846_ (.A(_01183_),
    .B(_14251_),
    .Y(_14568_));
 NOR2x1_ASAP7_75t_SL _22847_ (.A(_14188_),
    .B(_14227_),
    .Y(_14569_));
 OAI21x1_ASAP7_75t_SL _22849_ (.A1(_14569_),
    .A2(_14480_),
    .B(_14260_),
    .Y(_14571_));
 AOI21x1_ASAP7_75t_SL _22850_ (.A1(_14568_),
    .A2(_14571_),
    .B(_14278_),
    .Y(_14572_));
 NOR3x1_ASAP7_75t_SL _22851_ (.A(_14229_),
    .B(_14228_),
    .C(_14255_),
    .Y(_14573_));
 NOR2x1_ASAP7_75t_SL _22852_ (.A(_01168_),
    .B(_14230_),
    .Y(_14574_));
 OAI21x1_ASAP7_75t_SL _22853_ (.A1(_14573_),
    .A2(_14574_),
    .B(_14260_),
    .Y(_14575_));
 NOR2x1_ASAP7_75t_SL _22854_ (.A(_14308_),
    .B(_14222_),
    .Y(_14576_));
 OAI21x1_ASAP7_75t_SL _22855_ (.A1(_14284_),
    .A2(_14576_),
    .B(_14251_),
    .Y(_14577_));
 AOI21x1_ASAP7_75t_SL _22856_ (.A1(_14575_),
    .A2(_14577_),
    .B(_14289_),
    .Y(_14578_));
 OAI21x1_ASAP7_75t_SL _22857_ (.A1(_14572_),
    .A2(_14578_),
    .B(_14300_),
    .Y(_14579_));
 OA21x2_ASAP7_75t_SL _22858_ (.A1(_14260_),
    .A2(_01181_),
    .B(_14289_),
    .Y(_14580_));
 NAND2x1_ASAP7_75t_SL _22859_ (.A(_14386_),
    .B(_14358_),
    .Y(_14581_));
 AOI21x1_ASAP7_75t_SL _22860_ (.A1(_14580_),
    .A2(_14581_),
    .B(_14300_),
    .Y(_14582_));
 AO21x1_ASAP7_75t_SL _22861_ (.A1(_14448_),
    .A2(_14443_),
    .B(_14251_),
    .Y(_14583_));
 NAND2x1_ASAP7_75t_SL _22862_ (.A(_14520_),
    .B(_14514_),
    .Y(_14584_));
 AOI21x1_ASAP7_75t_SL _22863_ (.A1(_14251_),
    .A2(_14584_),
    .B(_14289_),
    .Y(_14585_));
 NAND2x1_ASAP7_75t_SL _22864_ (.A(_14583_),
    .B(_14585_),
    .Y(_14586_));
 NAND2x1_ASAP7_75t_SL _22865_ (.A(_14582_),
    .B(_14586_),
    .Y(_14587_));
 AOI21x1_ASAP7_75t_SL _22866_ (.A1(_14579_),
    .A2(_14587_),
    .B(_14331_),
    .Y(_14588_));
 NAND2x1_ASAP7_75t_SL _22867_ (.A(_01180_),
    .B(_14260_),
    .Y(_14589_));
 AOI21x1_ASAP7_75t_SL _22868_ (.A1(_14589_),
    .A2(_14551_),
    .B(_14278_),
    .Y(_14590_));
 AO21x1_ASAP7_75t_SL _22869_ (.A1(_14250_),
    .A2(_14245_),
    .B(_01185_),
    .Y(_14591_));
 OAI21x1_ASAP7_75t_SL _22870_ (.A1(_14227_),
    .A2(_14230_),
    .B(_14188_),
    .Y(_14592_));
 NAND2x1_ASAP7_75t_SL _22871_ (.A(_14260_),
    .B(_14592_),
    .Y(_14593_));
 AOI21x1_ASAP7_75t_SL _22872_ (.A1(_14591_),
    .A2(_14593_),
    .B(_14289_),
    .Y(_14594_));
 OAI21x1_ASAP7_75t_SL _22873_ (.A1(_14590_),
    .A2(_14594_),
    .B(_14300_),
    .Y(_14595_));
 NOR2x1_ASAP7_75t_SL _22874_ (.A(_14260_),
    .B(_14341_),
    .Y(_14596_));
 INVx1_ASAP7_75t_SL _22875_ (.A(_14596_),
    .Y(_14597_));
 AO21x1_ASAP7_75t_SL _22876_ (.A1(_14305_),
    .A2(_14380_),
    .B(_14251_),
    .Y(_14598_));
 NAND3x1_ASAP7_75t_SL _22877_ (.A(_14598_),
    .B(_14597_),
    .C(_14289_),
    .Y(_14599_));
 AND2x2_ASAP7_75t_R _22878_ (.A(_01171_),
    .B(_01169_),
    .Y(_14600_));
 INVx1_ASAP7_75t_SL _22879_ (.A(_14600_),
    .Y(_14601_));
 NAND2x1_ASAP7_75t_SL _22880_ (.A(_14601_),
    .B(_14230_),
    .Y(_14602_));
 INVx1_ASAP7_75t_SL _22881_ (.A(_14602_),
    .Y(_14603_));
 OAI21x1_ASAP7_75t_SL _22882_ (.A1(_14603_),
    .A2(_14553_),
    .B(_14260_),
    .Y(_14604_));
 AOI21x1_ASAP7_75t_SL _22883_ (.A1(_14364_),
    .A2(_14471_),
    .B(_14289_),
    .Y(_14605_));
 AOI21x1_ASAP7_75t_SL _22884_ (.A1(_14604_),
    .A2(_14605_),
    .B(_14300_),
    .Y(_14606_));
 NAND2x1_ASAP7_75t_SL _22885_ (.A(_14599_),
    .B(_14606_),
    .Y(_14607_));
 AOI21x1_ASAP7_75t_SL _22886_ (.A1(_14607_),
    .A2(_14595_),
    .B(_14332_),
    .Y(_14608_));
 OAI21x1_ASAP7_75t_SL _22887_ (.A1(_14588_),
    .A2(_14608_),
    .B(_14434_),
    .Y(_14609_));
 NAND2x1_ASAP7_75t_SL _22888_ (.A(_14609_),
    .B(_14567_),
    .Y(_00074_));
 NOR2x1_ASAP7_75t_SL _22889_ (.A(_14254_),
    .B(_14531_),
    .Y(_14610_));
 AOI21x1_ASAP7_75t_SL _22890_ (.A1(_14278_),
    .A2(_14610_),
    .B(_14301_),
    .Y(_14611_));
 NAND2x1_ASAP7_75t_R _22891_ (.A(_14315_),
    .B(_14222_),
    .Y(_14612_));
 AO21x1_ASAP7_75t_SL _22892_ (.A1(_14612_),
    .A2(_14602_),
    .B(_14251_),
    .Y(_14613_));
 NAND2x1_ASAP7_75t_SL _22893_ (.A(_14613_),
    .B(_14472_),
    .Y(_14614_));
 AOI21x1_ASAP7_75t_SL _22894_ (.A1(_14611_),
    .A2(_14614_),
    .B(_14331_),
    .Y(_14615_));
 AO21x1_ASAP7_75t_SL _22895_ (.A1(_14487_),
    .A2(_14380_),
    .B(_14260_),
    .Y(_14616_));
 AO21x1_ASAP7_75t_SL _22896_ (.A1(_14419_),
    .A2(_14316_),
    .B(_14251_),
    .Y(_14617_));
 AOI21x1_ASAP7_75t_SL _22897_ (.A1(_14616_),
    .A2(_14617_),
    .B(_14289_),
    .Y(_14618_));
 INVx1_ASAP7_75t_SL _22898_ (.A(_14506_),
    .Y(_14619_));
 AOI21x1_ASAP7_75t_SL _22899_ (.A1(_14619_),
    .A2(_14343_),
    .B(_14278_),
    .Y(_14620_));
 OAI21x1_ASAP7_75t_SL _22900_ (.A1(_14618_),
    .A2(_14620_),
    .B(_14301_),
    .Y(_14621_));
 AOI21x1_ASAP7_75t_SL _22901_ (.A1(_14615_),
    .A2(_14621_),
    .B(_14434_),
    .Y(_14622_));
 OAI21x1_ASAP7_75t_SL _22902_ (.A1(_14318_),
    .A2(_14260_),
    .B(_14301_),
    .Y(_14623_));
 AO21x1_ASAP7_75t_SL _22903_ (.A1(_14236_),
    .A2(_14260_),
    .B(_14301_),
    .Y(_14624_));
 AO21x1_ASAP7_75t_SL _22904_ (.A1(_14488_),
    .A2(_14364_),
    .B(_14624_),
    .Y(_14625_));
 INVx1_ASAP7_75t_SL _22905_ (.A(_14366_),
    .Y(_14626_));
 AOI21x1_ASAP7_75t_SL _22906_ (.A1(_14623_),
    .A2(_14625_),
    .B(_14626_),
    .Y(_14627_));
 INVx1_ASAP7_75t_R _22907_ (.A(_14316_),
    .Y(_14628_));
 NAND2x1_ASAP7_75t_SL _22908_ (.A(_14260_),
    .B(_14628_),
    .Y(_14629_));
 NAND3x1_ASAP7_75t_SL _22909_ (.A(_14541_),
    .B(_14301_),
    .C(_14629_),
    .Y(_14630_));
 AO21x1_ASAP7_75t_SL _22910_ (.A1(_14602_),
    .A2(_14487_),
    .B(_14251_),
    .Y(_14631_));
 NAND2x1_ASAP7_75t_SL _22911_ (.A(_14310_),
    .B(_14380_),
    .Y(_14632_));
 AOI21x1_ASAP7_75t_SL _22912_ (.A1(_14251_),
    .A2(_14632_),
    .B(_14301_),
    .Y(_14633_));
 NAND2x1_ASAP7_75t_SL _22913_ (.A(_14631_),
    .B(_14633_),
    .Y(_14634_));
 AOI21x1_ASAP7_75t_SL _22914_ (.A1(_14630_),
    .A2(_14634_),
    .B(_14278_),
    .Y(_14635_));
 OAI21x1_ASAP7_75t_SL _22915_ (.A1(_14635_),
    .A2(_14627_),
    .B(_14331_),
    .Y(_14636_));
 NAND2x1_ASAP7_75t_SL _22916_ (.A(_14622_),
    .B(_14636_),
    .Y(_14637_));
 AOI211x1_ASAP7_75t_SL _22917_ (.A1(_14335_),
    .A2(_14222_),
    .B(_14251_),
    .C(_14573_),
    .Y(_14638_));
 OAI21x1_ASAP7_75t_SL _22918_ (.A1(_14485_),
    .A2(_14501_),
    .B(_14289_),
    .Y(_14639_));
 NOR2x1_ASAP7_75t_SL _22919_ (.A(_14638_),
    .B(_14639_),
    .Y(_14640_));
 OAI21x1_ASAP7_75t_SL _22920_ (.A1(_14257_),
    .A2(_14401_),
    .B(_14278_),
    .Y(_14641_));
 NAND2x1_ASAP7_75t_SL _22921_ (.A(_14310_),
    .B(_14396_),
    .Y(_14642_));
 INVx1_ASAP7_75t_SL _22922_ (.A(_14642_),
    .Y(_14643_));
 OAI21x1_ASAP7_75t_SL _22923_ (.A1(_14641_),
    .A2(_14643_),
    .B(_14301_),
    .Y(_14644_));
 NOR2x1_ASAP7_75t_SL _22924_ (.A(_14640_),
    .B(_14644_),
    .Y(_14645_));
 INVx1_ASAP7_75t_R _22925_ (.A(_14310_),
    .Y(_14646_));
 NAND2x1_ASAP7_75t_SL _22926_ (.A(_14308_),
    .B(_14227_),
    .Y(_14647_));
 NAND2x1_ASAP7_75t_SL _22927_ (.A(_14289_),
    .B(_14647_),
    .Y(_14648_));
 NOR2x1_ASAP7_75t_SL _22928_ (.A(_14646_),
    .B(_14648_),
    .Y(_14649_));
 OAI21x1_ASAP7_75t_SL _22929_ (.A1(_14222_),
    .A2(_14251_),
    .B(_14649_),
    .Y(_14650_));
 NAND2x1_ASAP7_75t_R _22930_ (.A(_01174_),
    .B(_14222_),
    .Y(_14651_));
 INVx3_ASAP7_75t_SL _22931_ (.A(_14548_),
    .Y(_14652_));
 NAND2x1p5_ASAP7_75t_SL _22932_ (.A(_14651_),
    .B(_14652_),
    .Y(_14653_));
 NAND2x1_ASAP7_75t_SL _22933_ (.A(_14653_),
    .B(_14490_),
    .Y(_14654_));
 AOI21x1_ASAP7_75t_SL _22934_ (.A1(_14654_),
    .A2(_14650_),
    .B(_14301_),
    .Y(_14655_));
 OAI21x1_ASAP7_75t_SL _22935_ (.A1(_14655_),
    .A2(_14645_),
    .B(_14332_),
    .Y(_14656_));
 NAND2x1p5_ASAP7_75t_SL _22936_ (.A(_14389_),
    .B(_14652_),
    .Y(_14657_));
 AO21x1_ASAP7_75t_SL _22937_ (.A1(_14426_),
    .A2(_14305_),
    .B(_14251_),
    .Y(_14658_));
 AOI21x1_ASAP7_75t_SL _22938_ (.A1(_14658_),
    .A2(_14657_),
    .B(_14278_),
    .Y(_14659_));
 AO21x1_ASAP7_75t_SL _22939_ (.A1(_14341_),
    .A2(_14520_),
    .B(_14251_),
    .Y(_14660_));
 AO21x1_ASAP7_75t_SL _22940_ (.A1(_14310_),
    .A2(_14403_),
    .B(_14260_),
    .Y(_14661_));
 AOI21x1_ASAP7_75t_SL _22941_ (.A1(_14660_),
    .A2(_14661_),
    .B(_14289_),
    .Y(_14662_));
 OAI21x1_ASAP7_75t_SL _22942_ (.A1(_14662_),
    .A2(_14659_),
    .B(_14301_),
    .Y(_14663_));
 AO21x1_ASAP7_75t_SL _22943_ (.A1(_14448_),
    .A2(_14443_),
    .B(_14260_),
    .Y(_14664_));
 AOI21x1_ASAP7_75t_SL _22944_ (.A1(_14387_),
    .A2(_14664_),
    .B(_14301_),
    .Y(_14665_));
 AOI21x1_ASAP7_75t_SL _22945_ (.A1(_14389_),
    .A2(_14320_),
    .B(_14278_),
    .Y(_14666_));
 OAI21x1_ASAP7_75t_SL _22946_ (.A1(_14449_),
    .A2(_14357_),
    .B(_14666_),
    .Y(_14667_));
 AOI21x1_ASAP7_75t_SL _22947_ (.A1(_14665_),
    .A2(_14667_),
    .B(_14332_),
    .Y(_14668_));
 AOI21x1_ASAP7_75t_SL _22948_ (.A1(_14668_),
    .A2(_14663_),
    .B(_14376_),
    .Y(_14669_));
 NAND2x1_ASAP7_75t_SL _22949_ (.A(_14669_),
    .B(_14656_),
    .Y(_14670_));
 NAND2x1_ASAP7_75t_SL _22950_ (.A(_14637_),
    .B(_14670_),
    .Y(_00075_));
 AOI21x1_ASAP7_75t_SL _22951_ (.A1(_14288_),
    .A2(_14642_),
    .B(_14278_),
    .Y(_14671_));
 AO21x1_ASAP7_75t_SL _22952_ (.A1(_14514_),
    .A2(_14455_),
    .B(_14260_),
    .Y(_14672_));
 NAND2x1_ASAP7_75t_SL _22953_ (.A(_14448_),
    .B(_14360_),
    .Y(_14673_));
 AOI21x1_ASAP7_75t_SL _22954_ (.A1(_14672_),
    .A2(_14673_),
    .B(_14289_),
    .Y(_14674_));
 OAI21x1_ASAP7_75t_SL _22955_ (.A1(_14671_),
    .A2(_14674_),
    .B(_14300_),
    .Y(_14675_));
 AOI21x1_ASAP7_75t_SL _22956_ (.A1(_14514_),
    .A2(_14360_),
    .B(_14289_),
    .Y(_14676_));
 OAI21x1_ASAP7_75t_SL _22957_ (.A1(_14260_),
    .A2(_14336_),
    .B(_14676_),
    .Y(_14677_));
 OAI22x1_ASAP7_75t_SL _22958_ (.A1(_14507_),
    .A2(_01168_),
    .B1(_01175_),
    .B2(_14260_),
    .Y(_14678_));
 AOI21x1_ASAP7_75t_SL _22959_ (.A1(_14289_),
    .A2(_14678_),
    .B(_14300_),
    .Y(_14679_));
 AOI21x1_ASAP7_75t_SL _22960_ (.A1(_14677_),
    .A2(_14679_),
    .B(_14332_),
    .Y(_14680_));
 NAND2x1_ASAP7_75t_SL _22961_ (.A(_14675_),
    .B(_14680_),
    .Y(_14681_));
 NAND2x1_ASAP7_75t_SL _22962_ (.A(_14289_),
    .B(_14311_),
    .Y(_14682_));
 AO21x1_ASAP7_75t_SL _22963_ (.A1(_01171_),
    .A2(_14230_),
    .B(_14260_),
    .Y(_14683_));
 NOR2x1_ASAP7_75t_SL _22964_ (.A(_14574_),
    .B(_14683_),
    .Y(_14684_));
 AO21x1_ASAP7_75t_SL _22965_ (.A1(_14400_),
    .A2(_14222_),
    .B(_14251_),
    .Y(_14685_));
 OA21x2_ASAP7_75t_SL _22966_ (.A1(_14458_),
    .A2(_14260_),
    .B(_14278_),
    .Y(_14686_));
 AOI21x1_ASAP7_75t_SL _22967_ (.A1(_14685_),
    .A2(_14686_),
    .B(_14300_),
    .Y(_14687_));
 OAI21x1_ASAP7_75t_SL _22968_ (.A1(_14682_),
    .A2(_14684_),
    .B(_14687_),
    .Y(_14688_));
 NOR2x1_ASAP7_75t_SL _22969_ (.A(_14230_),
    .B(_14251_),
    .Y(_14689_));
 NOR2x1_ASAP7_75t_SL _22970_ (.A(_14278_),
    .B(_14689_),
    .Y(_14690_));
 NOR2x1_ASAP7_75t_SL _22971_ (.A(_14260_),
    .B(_14254_),
    .Y(_14691_));
 NAND2x1_ASAP7_75t_SL _22972_ (.A(_14414_),
    .B(_14691_),
    .Y(_14692_));
 AOI21x1_ASAP7_75t_SL _22973_ (.A1(_14690_),
    .A2(_14692_),
    .B(_14301_),
    .Y(_14693_));
 OA21x2_ASAP7_75t_SL _22974_ (.A1(_14389_),
    .A2(_14260_),
    .B(_14278_),
    .Y(_14694_));
 NOR2x1_ASAP7_75t_SL _22975_ (.A(_14596_),
    .B(_14445_),
    .Y(_14695_));
 NAND2x1_ASAP7_75t_SL _22976_ (.A(_14694_),
    .B(_14695_),
    .Y(_14696_));
 AOI21x1_ASAP7_75t_SL _22977_ (.A1(_14693_),
    .A2(_14696_),
    .B(_14331_),
    .Y(_14697_));
 AOI21x1_ASAP7_75t_SL _22978_ (.A1(_14688_),
    .A2(_14697_),
    .B(_14434_),
    .Y(_14698_));
 NAND2x1_ASAP7_75t_SL _22979_ (.A(_14681_),
    .B(_14698_),
    .Y(_14699_));
 AO21x1_ASAP7_75t_SL _22980_ (.A1(_14389_),
    .A2(_14335_),
    .B(_14260_),
    .Y(_14700_));
 AO21x1_ASAP7_75t_SL _22981_ (.A1(_14379_),
    .A2(_14488_),
    .B(_14251_),
    .Y(_14701_));
 AOI21x1_ASAP7_75t_SL _22982_ (.A1(_14700_),
    .A2(_14701_),
    .B(_14289_),
    .Y(_14702_));
 NAND2x1_ASAP7_75t_SL _22983_ (.A(_14443_),
    .B(_14691_),
    .Y(_14703_));
 AOI21x1_ASAP7_75t_SL _22984_ (.A1(_14571_),
    .A2(_14703_),
    .B(_14278_),
    .Y(_14704_));
 OAI21x1_ASAP7_75t_SL _22985_ (.A1(_14702_),
    .A2(_14704_),
    .B(_14300_),
    .Y(_14705_));
 NAND2x1_ASAP7_75t_SL _22986_ (.A(_14278_),
    .B(_14354_),
    .Y(_14706_));
 OA21x2_ASAP7_75t_SL _22987_ (.A1(_14360_),
    .A2(_14706_),
    .B(_14301_),
    .Y(_14707_));
 NAND2x1_ASAP7_75t_SL _22988_ (.A(_14260_),
    .B(_14443_),
    .Y(_14708_));
 AO21x1_ASAP7_75t_SL _22989_ (.A1(_14708_),
    .A2(_14475_),
    .B(_14474_),
    .Y(_14709_));
 NAND2x1_ASAP7_75t_SL _22990_ (.A(_14289_),
    .B(_14709_),
    .Y(_14710_));
 AOI21x1_ASAP7_75t_SL _22991_ (.A1(_14707_),
    .A2(_14710_),
    .B(_14331_),
    .Y(_14711_));
 NAND2x1_ASAP7_75t_SL _22992_ (.A(_14705_),
    .B(_14711_),
    .Y(_14712_));
 INVx1_ASAP7_75t_SL _22993_ (.A(_14337_),
    .Y(_14713_));
 OAI21x1_ASAP7_75t_SL _22994_ (.A1(_14251_),
    .A2(_14341_),
    .B(_14289_),
    .Y(_14714_));
 AND3x1_ASAP7_75t_SL _22995_ (.A(_14260_),
    .B(_14188_),
    .C(_14222_),
    .Y(_14715_));
 NOR2x1_ASAP7_75t_SL _22996_ (.A(_14714_),
    .B(_14715_),
    .Y(_14716_));
 NAND2x1_ASAP7_75t_SL _22997_ (.A(_14713_),
    .B(_14716_),
    .Y(_14717_));
 NOR2x1_ASAP7_75t_SL _22998_ (.A(_14222_),
    .B(_14357_),
    .Y(_14718_));
 OAI21x1_ASAP7_75t_SL _22999_ (.A1(_14480_),
    .A2(_14718_),
    .B(_14260_),
    .Y(_14719_));
 NOR2x1_ASAP7_75t_SL _23000_ (.A(_14289_),
    .B(_14560_),
    .Y(_14720_));
 AOI21x1_ASAP7_75t_SL _23001_ (.A1(_14719_),
    .A2(_14720_),
    .B(_14301_),
    .Y(_14721_));
 NAND2x1_ASAP7_75t_SL _23002_ (.A(_14717_),
    .B(_14721_),
    .Y(_14722_));
 OA21x2_ASAP7_75t_SL _23003_ (.A1(_14346_),
    .A2(_14251_),
    .B(_14316_),
    .Y(_14723_));
 AOI21x1_ASAP7_75t_SL _23004_ (.A1(_14314_),
    .A2(_14723_),
    .B(_14300_),
    .Y(_14724_));
 NOR2x1_ASAP7_75t_SL _23005_ (.A(_14260_),
    .B(_14519_),
    .Y(_14725_));
 AOI21x1_ASAP7_75t_SL _23006_ (.A1(_14520_),
    .A2(_14725_),
    .B(_14278_),
    .Y(_14726_));
 NAND2x1_ASAP7_75t_SL _23007_ (.A(_14361_),
    .B(_14726_),
    .Y(_14727_));
 AOI21x1_ASAP7_75t_SL _23008_ (.A1(_14724_),
    .A2(_14727_),
    .B(_14332_),
    .Y(_14728_));
 AOI21x1_ASAP7_75t_SL _23009_ (.A1(_14722_),
    .A2(_14728_),
    .B(_14376_),
    .Y(_14729_));
 NAND2x1_ASAP7_75t_SL _23010_ (.A(_14712_),
    .B(_14729_),
    .Y(_14730_));
 NAND2x1_ASAP7_75t_SL _23011_ (.A(_14699_),
    .B(_14730_),
    .Y(_00076_));
 NOR2x1_ASAP7_75t_SL _23012_ (.A(_14260_),
    .B(_14448_),
    .Y(_14731_));
 OA21x2_ASAP7_75t_SL _23013_ (.A1(_14383_),
    .A2(_14251_),
    .B(_14278_),
    .Y(_14732_));
 AO21x1_ASAP7_75t_SL _23014_ (.A1(_14309_),
    .A2(_14487_),
    .B(_14260_),
    .Y(_14733_));
 AOI21x1_ASAP7_75t_SL _23015_ (.A1(_14732_),
    .A2(_14733_),
    .B(_14301_),
    .Y(_14734_));
 OA21x2_ASAP7_75t_SL _23016_ (.A1(_14312_),
    .A2(_14731_),
    .B(_14734_),
    .Y(_14735_));
 OA21x2_ASAP7_75t_SL _23017_ (.A1(_14227_),
    .A2(_14251_),
    .B(_14289_),
    .Y(_14736_));
 AO21x1_ASAP7_75t_SL _23018_ (.A1(_14395_),
    .A2(_14736_),
    .B(_14300_),
    .Y(_14737_));
 AO21x1_ASAP7_75t_SL _23019_ (.A1(_14488_),
    .A2(_14612_),
    .B(_14260_),
    .Y(_14738_));
 NAND2x1_ASAP7_75t_SL _23020_ (.A(_14320_),
    .B(_14421_),
    .Y(_14739_));
 AND3x1_ASAP7_75t_SL _23021_ (.A(_14738_),
    .B(_14278_),
    .C(_14739_),
    .Y(_14740_));
 OAI21x1_ASAP7_75t_SL _23022_ (.A1(_14737_),
    .A2(_14740_),
    .B(_14332_),
    .Y(_14741_));
 NAND2x1_ASAP7_75t_SL _23023_ (.A(_14600_),
    .B(_14230_),
    .Y(_14742_));
 AOI21x1_ASAP7_75t_SL _23024_ (.A1(_14260_),
    .A2(_14742_),
    .B(_14278_),
    .Y(_14743_));
 OAI21x1_ASAP7_75t_SL _23025_ (.A1(_14464_),
    .A2(_14551_),
    .B(_14743_),
    .Y(_14744_));
 NAND2x1_ASAP7_75t_SL _23026_ (.A(_14260_),
    .B(_14414_),
    .Y(_14745_));
 AOI21x1_ASAP7_75t_SL _23027_ (.A1(_14745_),
    .A2(_14314_),
    .B(_14300_),
    .Y(_14746_));
 AOI21x1_ASAP7_75t_SL _23028_ (.A1(_14744_),
    .A2(_14746_),
    .B(_14332_),
    .Y(_14747_));
 NOR2x1_ASAP7_75t_SL _23029_ (.A(_14363_),
    .B(_14319_),
    .Y(_14748_));
 AO21x1_ASAP7_75t_SL _23030_ (.A1(_14414_),
    .A2(_14652_),
    .B(_14289_),
    .Y(_14749_));
 OA21x2_ASAP7_75t_SL _23031_ (.A1(_14251_),
    .A2(_14255_),
    .B(_14289_),
    .Y(_14750_));
 AO21x1_ASAP7_75t_SL _23032_ (.A1(_14400_),
    .A2(_14230_),
    .B(_14260_),
    .Y(_14751_));
 AOI21x1_ASAP7_75t_SL _23033_ (.A1(_14750_),
    .A2(_14751_),
    .B(_14301_),
    .Y(_14752_));
 OAI21x1_ASAP7_75t_SL _23034_ (.A1(_14749_),
    .A2(_14748_),
    .B(_14752_),
    .Y(_14753_));
 AOI21x1_ASAP7_75t_SL _23035_ (.A1(_14747_),
    .A2(_14753_),
    .B(_14434_),
    .Y(_14754_));
 OAI21x1_ASAP7_75t_SL _23036_ (.A1(_14735_),
    .A2(_14741_),
    .B(_14754_),
    .Y(_14755_));
 AO21x1_ASAP7_75t_SL _23037_ (.A1(_14354_),
    .A2(_01171_),
    .B(_14251_),
    .Y(_14756_));
 AO21x1_ASAP7_75t_SL _23038_ (.A1(_14336_),
    .A2(_14612_),
    .B(_14260_),
    .Y(_14757_));
 NAND2x1_ASAP7_75t_SL _23039_ (.A(_14756_),
    .B(_14757_),
    .Y(_14758_));
 NAND2x1_ASAP7_75t_SL _23040_ (.A(_14414_),
    .B(_14281_),
    .Y(_14759_));
 NAND2x1_ASAP7_75t_SL _23041_ (.A(_14389_),
    .B(_14354_),
    .Y(_14760_));
 AOI21x1_ASAP7_75t_SL _23042_ (.A1(_14251_),
    .A2(_14760_),
    .B(_14278_),
    .Y(_14761_));
 AOI21x1_ASAP7_75t_SL _23043_ (.A1(_14759_),
    .A2(_14761_),
    .B(_14331_),
    .Y(_14762_));
 OAI21x1_ASAP7_75t_SL _23044_ (.A1(_14289_),
    .A2(_14758_),
    .B(_14762_),
    .Y(_14763_));
 OA21x2_ASAP7_75t_SL _23045_ (.A1(_14251_),
    .A2(_14308_),
    .B(_14289_),
    .Y(_14764_));
 AOI21x1_ASAP7_75t_SL _23046_ (.A1(_14764_),
    .A2(_14700_),
    .B(_14332_),
    .Y(_14765_));
 NOR2x1_ASAP7_75t_SL _23047_ (.A(_14400_),
    .B(_14465_),
    .Y(_14766_));
 AND3x1_ASAP7_75t_SL _23048_ (.A(_14309_),
    .B(_14260_),
    .C(_14383_),
    .Y(_14767_));
 OAI21x1_ASAP7_75t_SL _23049_ (.A1(_14766_),
    .A2(_14767_),
    .B(_14278_),
    .Y(_14768_));
 AOI21x1_ASAP7_75t_SL _23050_ (.A1(_14765_),
    .A2(_14768_),
    .B(_14300_),
    .Y(_14769_));
 NAND2x1_ASAP7_75t_SL _23051_ (.A(_14763_),
    .B(_14769_),
    .Y(_14770_));
 AND2x2_ASAP7_75t_SL _23052_ (.A(_14401_),
    .B(_14289_),
    .Y(_14771_));
 AOI21x1_ASAP7_75t_SL _23053_ (.A1(_14771_),
    .A2(_14617_),
    .B(_14331_),
    .Y(_14772_));
 NOR2x1_ASAP7_75t_SL _23054_ (.A(_14289_),
    .B(_14508_),
    .Y(_14773_));
 NAND2x1_ASAP7_75t_SL _23055_ (.A(_14683_),
    .B(_14773_),
    .Y(_14774_));
 AOI21x1_ASAP7_75t_SL _23056_ (.A1(_14772_),
    .A2(_14774_),
    .B(_14301_),
    .Y(_14775_));
 NAND2x1_ASAP7_75t_SL _23057_ (.A(_14379_),
    .B(_14320_),
    .Y(_14776_));
 AO21x1_ASAP7_75t_SL _23058_ (.A1(_14776_),
    .A2(_14531_),
    .B(_14278_),
    .Y(_14777_));
 OA21x2_ASAP7_75t_SL _23059_ (.A1(_14346_),
    .A2(_14251_),
    .B(_14278_),
    .Y(_14778_));
 OR3x1_ASAP7_75t_SL _23060_ (.A(_14576_),
    .B(_14458_),
    .C(_14260_),
    .Y(_14779_));
 AOI21x1_ASAP7_75t_SL _23061_ (.A1(_14778_),
    .A2(_14779_),
    .B(_14332_),
    .Y(_14780_));
 NAND2x1_ASAP7_75t_SL _23062_ (.A(_14777_),
    .B(_14780_),
    .Y(_14781_));
 AOI21x1_ASAP7_75t_SL _23063_ (.A1(_14775_),
    .A2(_14781_),
    .B(_14376_),
    .Y(_14782_));
 NAND2x1_ASAP7_75t_SL _23064_ (.A(_14770_),
    .B(_14782_),
    .Y(_14783_));
 NAND2x1_ASAP7_75t_SL _23065_ (.A(_14755_),
    .B(_14783_),
    .Y(_00077_));
 INVx1_ASAP7_75t_SL _23066_ (.A(_14458_),
    .Y(_14784_));
 NOR2x1_ASAP7_75t_SL _23067_ (.A(_14251_),
    .B(_14237_),
    .Y(_14785_));
 AOI22x1_ASAP7_75t_SL _23068_ (.A1(_14652_),
    .A2(_14784_),
    .B1(_14785_),
    .B2(_14421_),
    .Y(_14786_));
 NOR2x1_ASAP7_75t_SL _23069_ (.A(_14289_),
    .B(_14391_),
    .Y(_14787_));
 NAND2x1_ASAP7_75t_SL _23070_ (.A(_14589_),
    .B(_14551_),
    .Y(_14788_));
 AOI21x1_ASAP7_75t_SL _23071_ (.A1(_14787_),
    .A2(_14788_),
    .B(_14300_),
    .Y(_14789_));
 OAI21x1_ASAP7_75t_SL _23072_ (.A1(_14278_),
    .A2(_14786_),
    .B(_14789_),
    .Y(_14790_));
 AOI21x1_ASAP7_75t_SL _23073_ (.A1(_14419_),
    .A2(_14336_),
    .B(_14251_),
    .Y(_14791_));
 AND3x1_ASAP7_75t_SL _23074_ (.A(_14346_),
    .B(_14742_),
    .C(_14251_),
    .Y(_14792_));
 OAI21x1_ASAP7_75t_SL _23075_ (.A1(_14791_),
    .A2(_14792_),
    .B(_14289_),
    .Y(_14793_));
 NOR2x1_ASAP7_75t_SL _23076_ (.A(_14260_),
    .B(_14383_),
    .Y(_14794_));
 NOR2x1_ASAP7_75t_SL _23077_ (.A(_14357_),
    .B(_14708_),
    .Y(_14795_));
 OAI21x1_ASAP7_75t_SL _23078_ (.A1(_14794_),
    .A2(_14795_),
    .B(_14278_),
    .Y(_14796_));
 NAND3x1_ASAP7_75t_SL _23079_ (.A(_14793_),
    .B(_14300_),
    .C(_14796_),
    .Y(_14797_));
 AOI21x1_ASAP7_75t_SL _23080_ (.A1(_14797_),
    .A2(_14790_),
    .B(_14332_),
    .Y(_14798_));
 AO21x1_ASAP7_75t_SL _23081_ (.A1(_14514_),
    .A2(_14455_),
    .B(_14251_),
    .Y(_14799_));
 AND2x2_ASAP7_75t_SL _23082_ (.A(_01178_),
    .B(_01184_),
    .Y(_14800_));
 OA21x2_ASAP7_75t_SL _23083_ (.A1(_14260_),
    .A2(_14800_),
    .B(_14289_),
    .Y(_14801_));
 AO21x1_ASAP7_75t_SL _23084_ (.A1(_14799_),
    .A2(_14801_),
    .B(_14300_),
    .Y(_14802_));
 OA21x2_ASAP7_75t_SL _23085_ (.A1(_14338_),
    .A2(_14628_),
    .B(_14260_),
    .Y(_14803_));
 NOR3x1_ASAP7_75t_SL _23086_ (.A(_14803_),
    .B(_14289_),
    .C(_14596_),
    .Y(_14804_));
 OAI21x1_ASAP7_75t_SL _23087_ (.A1(_14802_),
    .A2(_14804_),
    .B(_14332_),
    .Y(_14805_));
 NAND2x1_ASAP7_75t_SL _23088_ (.A(_14601_),
    .B(_14222_),
    .Y(_14806_));
 AO21x1_ASAP7_75t_SL _23089_ (.A1(_14806_),
    .A2(_14316_),
    .B(_14251_),
    .Y(_14807_));
 OAI21x1_ASAP7_75t_SL _23090_ (.A1(_14236_),
    .A2(_14474_),
    .B(_14251_),
    .Y(_14808_));
 AO21x1_ASAP7_75t_SL _23091_ (.A1(_14807_),
    .A2(_14808_),
    .B(_14289_),
    .Y(_14809_));
 AND3x1_ASAP7_75t_SL _23092_ (.A(_14459_),
    .B(_14651_),
    .C(_14251_),
    .Y(_14810_));
 OA21x2_ASAP7_75t_SL _23093_ (.A1(_14553_),
    .A2(_14285_),
    .B(_14260_),
    .Y(_14811_));
 OAI21x1_ASAP7_75t_SL _23094_ (.A1(_14810_),
    .A2(_14811_),
    .B(_14289_),
    .Y(_14812_));
 AOI21x1_ASAP7_75t_SL _23095_ (.A1(_14809_),
    .A2(_14812_),
    .B(_14301_),
    .Y(_14813_));
 OAI21x1_ASAP7_75t_SL _23096_ (.A1(_14805_),
    .A2(_14813_),
    .B(_14434_),
    .Y(_14814_));
 NAND2x1_ASAP7_75t_SL _23097_ (.A(_14289_),
    .B(_14557_),
    .Y(_14815_));
 INVx1_ASAP7_75t_SL _23098_ (.A(_14364_),
    .Y(_14816_));
 AOI21x1_ASAP7_75t_SL _23099_ (.A1(_14816_),
    .A2(_14676_),
    .B(_14301_),
    .Y(_14817_));
 NAND2x1_ASAP7_75t_SL _23100_ (.A(_14815_),
    .B(_14817_),
    .Y(_14818_));
 INVx2_ASAP7_75t_SL _23101_ (.A(_14380_),
    .Y(_14819_));
 OA21x2_ASAP7_75t_SL _23102_ (.A1(_14310_),
    .A2(_14260_),
    .B(_14278_),
    .Y(_14820_));
 OAI21x1_ASAP7_75t_SL _23103_ (.A1(_14819_),
    .A2(_14745_),
    .B(_14820_),
    .Y(_14821_));
 AOI21x1_ASAP7_75t_SL _23104_ (.A1(_01179_),
    .A2(_14260_),
    .B(_14278_),
    .Y(_14822_));
 AOI21x1_ASAP7_75t_SL _23105_ (.A1(_14822_),
    .A2(_14738_),
    .B(_14300_),
    .Y(_14823_));
 AOI21x1_ASAP7_75t_SL _23106_ (.A1(_14821_),
    .A2(_14823_),
    .B(_14332_),
    .Y(_14824_));
 NAND2x1_ASAP7_75t_SL _23107_ (.A(_14818_),
    .B(_14824_),
    .Y(_14825_));
 NAND2x1_ASAP7_75t_SL _23108_ (.A(_14535_),
    .B(_14548_),
    .Y(_14826_));
 AOI21x1_ASAP7_75t_SL _23109_ (.A1(_14227_),
    .A2(_14689_),
    .B(_14278_),
    .Y(_14827_));
 NAND2x1_ASAP7_75t_SL _23110_ (.A(_14827_),
    .B(_14826_),
    .Y(_14828_));
 AOI21x1_ASAP7_75t_SL _23111_ (.A1(_14413_),
    .A2(_14516_),
    .B(_14301_),
    .Y(_14829_));
 AOI21x1_ASAP7_75t_SL _23112_ (.A1(_14829_),
    .A2(_14828_),
    .B(_14331_),
    .Y(_14830_));
 AND2x2_ASAP7_75t_SL _23113_ (.A(_14647_),
    .B(_14260_),
    .Y(_14831_));
 OA21x2_ASAP7_75t_SL _23114_ (.A1(_14831_),
    .A2(_14725_),
    .B(_14310_),
    .Y(_14832_));
 NAND2x1_ASAP7_75t_SL _23115_ (.A(_14308_),
    .B(_14251_),
    .Y(_14833_));
 AOI21x1_ASAP7_75t_SL _23116_ (.A1(_14833_),
    .A2(_14649_),
    .B(_14300_),
    .Y(_14834_));
 OAI21x1_ASAP7_75t_SL _23117_ (.A1(_14289_),
    .A2(_14832_),
    .B(_14834_),
    .Y(_14835_));
 AOI21x1_ASAP7_75t_SL _23118_ (.A1(_14835_),
    .A2(_14830_),
    .B(_14434_),
    .Y(_14836_));
 NAND2x1_ASAP7_75t_SL _23119_ (.A(_14825_),
    .B(_14836_),
    .Y(_14837_));
 OAI21x1_ASAP7_75t_SL _23120_ (.A1(_14798_),
    .A2(_14814_),
    .B(_14837_),
    .Y(_00078_));
 AOI21x1_ASAP7_75t_SL _23121_ (.A1(_14742_),
    .A2(_14360_),
    .B(_14289_),
    .Y(_14838_));
 AO21x1_ASAP7_75t_SL _23122_ (.A1(_14419_),
    .A2(_14188_),
    .B(_14260_),
    .Y(_14839_));
 AO21x1_ASAP7_75t_SL _23123_ (.A1(_14838_),
    .A2(_14839_),
    .B(_14300_),
    .Y(_14840_));
 INVx1_ASAP7_75t_R _23124_ (.A(_14341_),
    .Y(_14841_));
 NOR2x1_ASAP7_75t_SL _23125_ (.A(_14841_),
    .B(_14553_),
    .Y(_14842_));
 AOI22x1_ASAP7_75t_SL _23126_ (.A1(_14320_),
    .A2(_14383_),
    .B1(_14842_),
    .B2(_14251_),
    .Y(_14843_));
 NOR2x1_ASAP7_75t_SL _23127_ (.A(_14278_),
    .B(_14843_),
    .Y(_14844_));
 OA21x2_ASAP7_75t_SL _23128_ (.A1(_14260_),
    .A2(_01171_),
    .B(_14278_),
    .Y(_14845_));
 NAND2x1_ASAP7_75t_SL _23129_ (.A(_14845_),
    .B(_14799_),
    .Y(_14846_));
 OA21x2_ASAP7_75t_SL _23130_ (.A1(_14389_),
    .A2(_14251_),
    .B(_14341_),
    .Y(_14847_));
 AOI21x1_ASAP7_75t_SL _23131_ (.A1(_14339_),
    .A2(_14847_),
    .B(_14301_),
    .Y(_14848_));
 AOI21x1_ASAP7_75t_SL _23132_ (.A1(_14846_),
    .A2(_14848_),
    .B(_14376_),
    .Y(_14849_));
 OAI21x1_ASAP7_75t_SL _23133_ (.A1(_14840_),
    .A2(_14844_),
    .B(_14849_),
    .Y(_14850_));
 NAND2x1_ASAP7_75t_SL _23134_ (.A(_14289_),
    .B(_14583_),
    .Y(_14851_));
 AO21x1_ASAP7_75t_SL _23135_ (.A1(_14380_),
    .A2(_14310_),
    .B(_14260_),
    .Y(_14852_));
 AOI21x1_ASAP7_75t_SL _23136_ (.A1(_14459_),
    .A2(_14386_),
    .B(_14289_),
    .Y(_14853_));
 AOI21x1_ASAP7_75t_SL _23137_ (.A1(_14852_),
    .A2(_14853_),
    .B(_14301_),
    .Y(_14854_));
 OAI21x1_ASAP7_75t_SL _23138_ (.A1(_14810_),
    .A2(_14851_),
    .B(_14854_),
    .Y(_14855_));
 OAI21x1_ASAP7_75t_SL _23139_ (.A1(_14841_),
    .A2(_14553_),
    .B(_14260_),
    .Y(_14856_));
 AO21x1_ASAP7_75t_R _23140_ (.A1(_14230_),
    .A2(_14308_),
    .B(_14205_),
    .Y(_14857_));
 AOI21x1_ASAP7_75t_SL _23141_ (.A1(_14251_),
    .A2(_14857_),
    .B(_14289_),
    .Y(_14858_));
 NAND2x1_ASAP7_75t_SL _23142_ (.A(_14856_),
    .B(_14858_),
    .Y(_14859_));
 AO21x1_ASAP7_75t_SL _23143_ (.A1(_14488_),
    .A2(_14612_),
    .B(_14251_),
    .Y(_14860_));
 OA21x2_ASAP7_75t_SL _23144_ (.A1(_14519_),
    .A2(_14260_),
    .B(_14289_),
    .Y(_14861_));
 AOI21x1_ASAP7_75t_SL _23145_ (.A1(_14860_),
    .A2(_14861_),
    .B(_14300_),
    .Y(_14862_));
 AOI21x1_ASAP7_75t_SL _23146_ (.A1(_14859_),
    .A2(_14862_),
    .B(_14434_),
    .Y(_14863_));
 AOI21x1_ASAP7_75t_SL _23147_ (.A1(_14855_),
    .A2(_14863_),
    .B(_14331_),
    .Y(_14864_));
 NAND2x1_ASAP7_75t_SL _23148_ (.A(_14850_),
    .B(_14864_),
    .Y(_14865_));
 NAND2x1_ASAP7_75t_SL _23149_ (.A(_14251_),
    .B(_14236_),
    .Y(_14866_));
 OAI21x1_ASAP7_75t_R _23150_ (.A1(_01184_),
    .A2(_14251_),
    .B(_14289_),
    .Y(_14867_));
 NOR2x1_ASAP7_75t_SL _23151_ (.A(_14317_),
    .B(_14867_),
    .Y(_14868_));
 AOI21x1_ASAP7_75t_SL _23152_ (.A1(_14866_),
    .A2(_14868_),
    .B(_14301_),
    .Y(_14869_));
 OA21x2_ASAP7_75t_SL _23153_ (.A1(_14819_),
    .A2(_14521_),
    .B(_14278_),
    .Y(_14870_));
 OAI21x1_ASAP7_75t_SL _23154_ (.A1(_14237_),
    .A2(_14465_),
    .B(_14870_),
    .Y(_14871_));
 AOI21x1_ASAP7_75t_SL _23155_ (.A1(_14869_),
    .A2(_14871_),
    .B(_14376_),
    .Y(_14872_));
 AO21x1_ASAP7_75t_SL _23156_ (.A1(_14230_),
    .A2(_14205_),
    .B(_14308_),
    .Y(_14873_));
 AOI21x1_ASAP7_75t_SL _23157_ (.A1(_14251_),
    .A2(_14873_),
    .B(_14445_),
    .Y(_14874_));
 NAND2x1_ASAP7_75t_SL _23158_ (.A(_01175_),
    .B(_14260_),
    .Y(_14875_));
 AO21x1_ASAP7_75t_SL _23159_ (.A1(_14339_),
    .A2(_14875_),
    .B(_14300_),
    .Y(_14876_));
 AO21x1_ASAP7_75t_SL _23160_ (.A1(_14278_),
    .A2(_14874_),
    .B(_14876_),
    .Y(_14877_));
 NAND2x1_ASAP7_75t_SL _23161_ (.A(_14872_),
    .B(_14877_),
    .Y(_14878_));
 NOR2x1_ASAP7_75t_SL _23162_ (.A(_14278_),
    .B(_14391_),
    .Y(_14879_));
 NAND2x1_ASAP7_75t_SL _23163_ (.A(_14260_),
    .B(_14485_),
    .Y(_14880_));
 AOI21x1_ASAP7_75t_SL _23164_ (.A1(_14879_),
    .A2(_14880_),
    .B(_14301_),
    .Y(_14881_));
 NAND2x1_ASAP7_75t_SL _23165_ (.A(_14222_),
    .B(_14400_),
    .Y(_14882_));
 NAND2x1p5_ASAP7_75t_SL _23166_ (.A(_14882_),
    .B(_14652_),
    .Y(_14883_));
 AOI21x1_ASAP7_75t_SL _23167_ (.A1(_14260_),
    .A2(_14358_),
    .B(_14289_),
    .Y(_14884_));
 NAND2x1_ASAP7_75t_SL _23168_ (.A(_14883_),
    .B(_14884_),
    .Y(_14885_));
 AOI21x1_ASAP7_75t_SL _23169_ (.A1(_14881_),
    .A2(_14885_),
    .B(_14434_),
    .Y(_14886_));
 NAND2x1_ASAP7_75t_SL _23170_ (.A(_14227_),
    .B(_14251_),
    .Y(_14887_));
 OAI21x1_ASAP7_75t_SL _23171_ (.A1(_14474_),
    .A2(_14708_),
    .B(_14887_),
    .Y(_14888_));
 NOR2x1_ASAP7_75t_SL _23172_ (.A(_14289_),
    .B(_14888_),
    .Y(_14889_));
 NAND2x1_ASAP7_75t_SL _23173_ (.A(_14882_),
    .B(_14428_),
    .Y(_14890_));
 AOI21x1_ASAP7_75t_SL _23174_ (.A1(_14571_),
    .A2(_14890_),
    .B(_14278_),
    .Y(_14891_));
 OAI21x1_ASAP7_75t_SL _23175_ (.A1(_14889_),
    .A2(_14891_),
    .B(_14301_),
    .Y(_14892_));
 AOI21x1_ASAP7_75t_SL _23176_ (.A1(_14892_),
    .A2(_14886_),
    .B(_14332_),
    .Y(_14893_));
 NAND2x1_ASAP7_75t_SL _23177_ (.A(_14878_),
    .B(_14893_),
    .Y(_14894_));
 NAND2x1_ASAP7_75t_SL _23178_ (.A(_14865_),
    .B(_14894_),
    .Y(_00079_));
 XOR2x2_ASAP7_75t_SL _23179_ (.A(_00655_),
    .B(_00662_),
    .Y(_14895_));
 XOR2x1_ASAP7_75t_SL _23180_ (.A(_00656_),
    .Y(_14896_),
    .B(_00688_));
 XOR2x2_ASAP7_75t_SL _23181_ (.A(_14895_),
    .B(_14896_),
    .Y(_14897_));
 XOR2x2_ASAP7_75t_SL _23182_ (.A(_12076_),
    .B(_00592_),
    .Y(_14898_));
 AND2x2_ASAP7_75t_SL _23183_ (.A(_14897_),
    .B(_14898_),
    .Y(_14899_));
 OAI21x1_ASAP7_75t_SL _23184_ (.A1(_14898_),
    .A2(_14897_),
    .B(_00574_),
    .Y(_14900_));
 NAND2x1_ASAP7_75t_SL _23185_ (.A(_00462_),
    .B(_10675_),
    .Y(_14901_));
 OAI21x1_ASAP7_75t_SL _23186_ (.A1(_14900_),
    .A2(_14899_),
    .B(_14901_),
    .Y(_14902_));
 XOR2x2_ASAP7_75t_SL _23187_ (.A(_14902_),
    .B(_00910_),
    .Y(_14903_));
 NOR2x1_ASAP7_75t_SL _23189_ (.A(_00574_),
    .B(_00463_),
    .Y(_14904_));
 INVx1_ASAP7_75t_SL _23190_ (.A(_14904_),
    .Y(_14905_));
 XOR2x2_ASAP7_75t_L _23191_ (.A(_00591_),
    .B(_00630_),
    .Y(_14906_));
 NAND2x1_ASAP7_75t_SL _23192_ (.A(_12097_),
    .B(_14906_),
    .Y(_14907_));
 XNOR2x2_ASAP7_75t_SL _23193_ (.A(_00591_),
    .B(_00630_),
    .Y(_14908_));
 NAND2x1_ASAP7_75t_SL _23194_ (.A(_00687_),
    .B(_14908_),
    .Y(_14909_));
 INVx1_ASAP7_75t_SL _23195_ (.A(_14895_),
    .Y(_14910_));
 AOI21x1_ASAP7_75t_SL _23196_ (.A1(_14909_),
    .A2(_14907_),
    .B(_14910_),
    .Y(_14911_));
 XOR2x2_ASAP7_75t_L _23197_ (.A(_00630_),
    .B(_00687_),
    .Y(_14912_));
 NAND2x1_ASAP7_75t_SL _23198_ (.A(_00591_),
    .B(_14912_),
    .Y(_14913_));
 INVx1_ASAP7_75t_R _23199_ (.A(_00591_),
    .Y(_14914_));
 XNOR2x2_ASAP7_75t_L _23200_ (.A(_00630_),
    .B(_00687_),
    .Y(_14915_));
 NAND2x1_ASAP7_75t_SL _23201_ (.A(_14914_),
    .B(_14915_),
    .Y(_14916_));
 AOI21x1_ASAP7_75t_SL _23202_ (.A1(_14913_),
    .A2(_14916_),
    .B(_14895_),
    .Y(_14917_));
 OAI21x1_ASAP7_75t_SL _23203_ (.A1(_14917_),
    .A2(_14911_),
    .B(_00574_),
    .Y(_14918_));
 NAND2x1_ASAP7_75t_SL _23204_ (.A(_14905_),
    .B(_14918_),
    .Y(_14919_));
 XNOR2x2_ASAP7_75t_SL _23205_ (.A(_00909_),
    .B(_14919_),
    .Y(_01193_));
 NOR2x1_ASAP7_75t_R _23206_ (.A(_00574_),
    .B(_00464_),
    .Y(_14920_));
 INVx1_ASAP7_75t_SL _23207_ (.A(_14920_),
    .Y(_14921_));
 INVx1_ASAP7_75t_R _23208_ (.A(_00593_),
    .Y(_14922_));
 NOR2x2_ASAP7_75t_SL _23209_ (.A(_14922_),
    .B(_12124_),
    .Y(_14923_));
 NOR2x1_ASAP7_75t_SL _23210_ (.A(_00593_),
    .B(_12120_),
    .Y(_14924_));
 OAI21x1_ASAP7_75t_SL _23211_ (.A1(_14923_),
    .A2(_14924_),
    .B(_12079_),
    .Y(_14925_));
 INVx1_ASAP7_75t_SL _23212_ (.A(_14925_),
    .Y(_14926_));
 NOR3x1_ASAP7_75t_L _23213_ (.A(_14924_),
    .B(_14923_),
    .C(_12079_),
    .Y(_14927_));
 OAI21x1_ASAP7_75t_SL _23214_ (.A1(_14926_),
    .A2(_14927_),
    .B(_00574_),
    .Y(_14928_));
 INVx1_ASAP7_75t_SL _23215_ (.A(_00911_),
    .Y(_14929_));
 AOI21x1_ASAP7_75t_SL _23216_ (.A1(_14921_),
    .A2(_14928_),
    .B(_14929_),
    .Y(_14930_));
 NAND2x1_ASAP7_75t_SL _23217_ (.A(_00464_),
    .B(_10675_),
    .Y(_14931_));
 INVx1_ASAP7_75t_R _23218_ (.A(_12079_),
    .Y(_14932_));
 XOR2x2_ASAP7_75t_SL _23219_ (.A(_12124_),
    .B(_14922_),
    .Y(_14933_));
 NAND2x1_ASAP7_75t_SL _23220_ (.A(_14932_),
    .B(_14933_),
    .Y(_14934_));
 NAND3x1_ASAP7_75t_SL _23221_ (.A(_14934_),
    .B(_00574_),
    .C(_14925_),
    .Y(_14935_));
 AOI21x1_ASAP7_75t_SL _23222_ (.A1(_14931_),
    .A2(_14935_),
    .B(_00911_),
    .Y(_14936_));
 NOR2x2_ASAP7_75t_SL _23223_ (.A(_14930_),
    .B(_14936_),
    .Y(_14937_));
 NAND3x1_ASAP7_75t_L _23225_ (.A(_14905_),
    .B(_00909_),
    .C(_14918_),
    .Y(_14938_));
 AO21x1_ASAP7_75t_SL _23226_ (.A1(_14918_),
    .A2(_14905_),
    .B(_00909_),
    .Y(_14939_));
 NAND2x2_ASAP7_75t_SL _23227_ (.A(_14939_),
    .B(_14938_),
    .Y(_01186_));
 AOI21x1_ASAP7_75t_SL _23228_ (.A1(_14921_),
    .A2(_14928_),
    .B(_00911_),
    .Y(_14940_));
 AOI21x1_ASAP7_75t_SL _23229_ (.A1(_14931_),
    .A2(_14935_),
    .B(_14929_),
    .Y(_14941_));
 NOR2x2_ASAP7_75t_SL _23230_ (.A(_14940_),
    .B(_14941_),
    .Y(_14942_));
 NOR2x1_ASAP7_75t_SL _23233_ (.A(_00574_),
    .B(_00522_),
    .Y(_14944_));
 XOR2x2_ASAP7_75t_SL _23234_ (.A(_00657_),
    .B(_00662_),
    .Y(_14945_));
 XNOR2x2_ASAP7_75t_SL _23235_ (.A(_12146_),
    .B(_14945_),
    .Y(_14946_));
 XNOR2x2_ASAP7_75t_SL _23236_ (.A(_00594_),
    .B(_12145_),
    .Y(_14947_));
 XOR2x2_ASAP7_75t_SL _23237_ (.A(_14946_),
    .B(_14947_),
    .Y(_14948_));
 NOR2x1_ASAP7_75t_SL _23238_ (.A(_10675_),
    .B(_14948_),
    .Y(_14949_));
 OAI21x1_ASAP7_75t_SL _23239_ (.A1(_14944_),
    .A2(_14949_),
    .B(_00912_),
    .Y(_14950_));
 XNOR2x1_ASAP7_75t_SL _23240_ (.B(_14946_),
    .Y(_14951_),
    .A(_14947_));
 NAND2x1_ASAP7_75t_SL _23241_ (.A(_00574_),
    .B(_14951_),
    .Y(_14952_));
 INVx1_ASAP7_75t_R _23242_ (.A(_00912_),
    .Y(_14953_));
 INVx1_ASAP7_75t_SL _23243_ (.A(_14944_),
    .Y(_14954_));
 NAND3x1_ASAP7_75t_SL _23244_ (.A(_14952_),
    .B(_14953_),
    .C(_14954_),
    .Y(_14955_));
 NAND2x1_ASAP7_75t_SL _23245_ (.A(_14950_),
    .B(_14955_),
    .Y(_14956_));
 INVx1_ASAP7_75t_R _23248_ (.A(_01190_),
    .Y(_14959_));
 OAI21x1_ASAP7_75t_SL _23249_ (.A1(_14930_),
    .A2(_14936_),
    .B(_14959_),
    .Y(_14960_));
 AND2x2_ASAP7_75t_R _23250_ (.A(_10675_),
    .B(_00521_),
    .Y(_14961_));
 XOR2x2_ASAP7_75t_R _23251_ (.A(_00595_),
    .B(_00659_),
    .Y(_14962_));
 XOR2x2_ASAP7_75t_SL _23252_ (.A(_12158_),
    .B(_14962_),
    .Y(_14963_));
 XOR2x2_ASAP7_75t_R _23253_ (.A(_00658_),
    .B(_00662_),
    .Y(_14964_));
 INVx1_ASAP7_75t_R _23254_ (.A(_00691_),
    .Y(_14965_));
 XOR2x2_ASAP7_75t_SL _23255_ (.A(_14964_),
    .B(_14965_),
    .Y(_14966_));
 XOR2x2_ASAP7_75t_SL _23256_ (.A(_14963_),
    .B(_14966_),
    .Y(_14967_));
 NOR2x1_ASAP7_75t_R _23257_ (.A(_10675_),
    .B(_14967_),
    .Y(_14968_));
 OAI21x1_ASAP7_75t_SL _23258_ (.A1(_14961_),
    .A2(_14968_),
    .B(_00914_),
    .Y(_14969_));
 NOR2x1_ASAP7_75t_R _23259_ (.A(_00574_),
    .B(_00521_),
    .Y(_14970_));
 XNOR2x2_ASAP7_75t_SL _23260_ (.A(_14966_),
    .B(_14963_),
    .Y(_14971_));
 NOR2x1_ASAP7_75t_R _23261_ (.A(_10675_),
    .B(_14971_),
    .Y(_14972_));
 INVx1_ASAP7_75t_R _23262_ (.A(_00914_),
    .Y(_14973_));
 OAI21x1_ASAP7_75t_SL _23263_ (.A1(_14970_),
    .A2(_14972_),
    .B(_14973_),
    .Y(_14974_));
 NAND2x1_ASAP7_75t_SL _23264_ (.A(_14969_),
    .B(_14974_),
    .Y(_14975_));
 OA21x2_ASAP7_75t_SL _23266_ (.A1(_14956_),
    .A2(_14960_),
    .B(_14975_),
    .Y(_14977_));
 XNOR2x2_ASAP7_75t_SL _23267_ (.A(_14902_),
    .B(_00910_),
    .Y(_01187_));
 NOR2x2_ASAP7_75t_SL _23268_ (.A(_01187_),
    .B(_01193_),
    .Y(_14978_));
 NAND2x2_ASAP7_75t_L _23269_ (.A(_14942_),
    .B(_14978_),
    .Y(_14979_));
 OAI21x1_ASAP7_75t_R _23270_ (.A1(_14944_),
    .A2(_14949_),
    .B(_14953_),
    .Y(_14980_));
 NAND3x1_ASAP7_75t_R _23271_ (.A(_14952_),
    .B(_00912_),
    .C(_14954_),
    .Y(_14981_));
 NAND2x1_ASAP7_75t_SL _23272_ (.A(_14980_),
    .B(_14981_),
    .Y(_14982_));
 INVx1_ASAP7_75t_SL _23274_ (.A(_01195_),
    .Y(_14984_));
 NOR2x2_ASAP7_75t_SL _23275_ (.A(_14984_),
    .B(_14942_),
    .Y(_14985_));
 NOR2x1_ASAP7_75t_SL _23276_ (.A(_14982_),
    .B(_14985_),
    .Y(_14986_));
 NAND2x1_ASAP7_75t_SL _23277_ (.A(_14979_),
    .B(_14986_),
    .Y(_14987_));
 NAND2x1_ASAP7_75t_SL _23278_ (.A(_14977_),
    .B(_14987_),
    .Y(_14988_));
 NOR2x1_ASAP7_75t_SL _23279_ (.A(_14960_),
    .B(_14982_),
    .Y(_14989_));
 NOR2x1_ASAP7_75t_SL _23280_ (.A(_14975_),
    .B(_14989_),
    .Y(_14990_));
 AOI21x1_ASAP7_75t_R _23281_ (.A1(_14925_),
    .A2(_14934_),
    .B(_10675_),
    .Y(_14991_));
 OAI21x1_ASAP7_75t_R _23282_ (.A1(_14920_),
    .A2(_14991_),
    .B(_14929_),
    .Y(_14992_));
 NAND3x1_ASAP7_75t_R _23283_ (.A(_14928_),
    .B(_00911_),
    .C(_14921_),
    .Y(_14993_));
 AOI21x1_ASAP7_75t_R _23284_ (.A1(_14992_),
    .A2(_14993_),
    .B(_01194_),
    .Y(_14994_));
 NOR2x1_ASAP7_75t_R _23285_ (.A(_14994_),
    .B(_14956_),
    .Y(_14995_));
 NAND2x1_ASAP7_75t_SL _23286_ (.A(_14995_),
    .B(_14979_),
    .Y(_14996_));
 XOR2x2_ASAP7_75t_L _23287_ (.A(_00661_),
    .B(_00693_),
    .Y(_14997_));
 XOR2x2_ASAP7_75t_R _23288_ (.A(_12190_),
    .B(_00597_),
    .Y(_14998_));
 XNOR2x2_ASAP7_75t_R _23289_ (.A(_14997_),
    .B(_14998_),
    .Y(_14999_));
 NOR2x1_ASAP7_75t_R _23290_ (.A(_00574_),
    .B(_00519_),
    .Y(_15000_));
 AO21x1_ASAP7_75t_SL _23291_ (.A1(_14999_),
    .A2(_00574_),
    .B(_15000_),
    .Y(_15001_));
 XOR2x2_ASAP7_75t_SL _23292_ (.A(_15001_),
    .B(_00916_),
    .Y(_15002_));
 INVx1_ASAP7_75t_SL _23293_ (.A(_15002_),
    .Y(_15003_));
 AOI21x1_ASAP7_75t_SL _23295_ (.A1(_14990_),
    .A2(_14996_),
    .B(_15003_),
    .Y(_15005_));
 XOR2x2_ASAP7_75t_SL _23296_ (.A(_00659_),
    .B(_00660_),
    .Y(_15006_));
 INVx1_ASAP7_75t_R _23297_ (.A(_00692_),
    .Y(_15007_));
 XOR2x2_ASAP7_75t_R _23298_ (.A(_15006_),
    .B(_15007_),
    .Y(_15008_));
 XNOR2x2_ASAP7_75t_R _23299_ (.A(_00596_),
    .B(_00627_),
    .Y(_15009_));
 XOR2x2_ASAP7_75t_SL _23300_ (.A(_15008_),
    .B(_15009_),
    .Y(_15010_));
 OR2x2_ASAP7_75t_R _23302_ (.A(_00574_),
    .B(_00520_),
    .Y(_15012_));
 OA21x2_ASAP7_75t_R _23303_ (.A1(_15010_),
    .A2(_10675_),
    .B(_15012_),
    .Y(_15013_));
 NOR2x1_ASAP7_75t_R _23304_ (.A(_00915_),
    .B(_15013_),
    .Y(_15014_));
 AND2x2_ASAP7_75t_SL _23305_ (.A(_15013_),
    .B(_00915_),
    .Y(_15015_));
 NOR2x1_ASAP7_75t_SL _23306_ (.A(_15014_),
    .B(_15015_),
    .Y(_15016_));
 INVx1_ASAP7_75t_SL _23307_ (.A(_15016_),
    .Y(_15017_));
 AOI21x1_ASAP7_75t_SL _23309_ (.A1(_14988_),
    .A2(_15005_),
    .B(_15017_),
    .Y(_15019_));
 OAI21x1_ASAP7_75t_SL _23311_ (.A1(_14930_),
    .A2(_14936_),
    .B(_01192_),
    .Y(_15021_));
 NAND2x1_ASAP7_75t_SL _23312_ (.A(_15021_),
    .B(_14956_),
    .Y(_15022_));
 OAI21x1_ASAP7_75t_SL _23313_ (.A1(_14940_),
    .A2(_14941_),
    .B(_01188_),
    .Y(_15023_));
 AO21x1_ASAP7_75t_SL _23315_ (.A1(_15023_),
    .A2(_14960_),
    .B(_14956_),
    .Y(_15025_));
 AOI21x1_ASAP7_75t_SL _23317_ (.A1(_15022_),
    .A2(_15025_),
    .B(_14975_),
    .Y(_15027_));
 NAND2x1_ASAP7_75t_SL _23318_ (.A(_01187_),
    .B(_14942_),
    .Y(_15028_));
 OAI21x1_ASAP7_75t_SL _23319_ (.A1(_14940_),
    .A2(_14941_),
    .B(_01189_),
    .Y(_15029_));
 AO21x1_ASAP7_75t_SL _23320_ (.A1(_15028_),
    .A2(_15029_),
    .B(_14956_),
    .Y(_15030_));
 NAND2x1_ASAP7_75t_SL _23321_ (.A(_01194_),
    .B(_14937_),
    .Y(_15031_));
 NAND2x2_ASAP7_75t_SL _23322_ (.A(_01193_),
    .B(_14942_),
    .Y(_15032_));
 AO21x1_ASAP7_75t_SL _23324_ (.A1(_15031_),
    .A2(_15032_),
    .B(_14982_),
    .Y(_15034_));
 INVx1_ASAP7_75t_SL _23325_ (.A(_14975_),
    .Y(_15035_));
 AOI21x1_ASAP7_75t_SL _23328_ (.A1(_15030_),
    .A2(_15034_),
    .B(_15035_),
    .Y(_15038_));
 OAI21x1_ASAP7_75t_SL _23329_ (.A1(_15027_),
    .A2(_15038_),
    .B(_15003_),
    .Y(_15039_));
 NAND2x1_ASAP7_75t_SL _23330_ (.A(_15019_),
    .B(_15039_),
    .Y(_15040_));
 NOR2x2_ASAP7_75t_SL _23332_ (.A(_01192_),
    .B(_14942_),
    .Y(_15042_));
 AOI21x1_ASAP7_75t_SL _23333_ (.A1(_14982_),
    .A2(_15042_),
    .B(_14975_),
    .Y(_15043_));
 OAI21x1_ASAP7_75t_SL _23334_ (.A1(_14930_),
    .A2(_14936_),
    .B(_14984_),
    .Y(_15044_));
 NOR2x1_ASAP7_75t_SL _23336_ (.A(_15044_),
    .B(_14956_),
    .Y(_15046_));
 OAI21x1_ASAP7_75t_SL _23337_ (.A1(_14930_),
    .A2(_14936_),
    .B(_01189_),
    .Y(_15047_));
 NAND2x2_ASAP7_75t_SL _23338_ (.A(_14956_),
    .B(_15047_),
    .Y(_15048_));
 INVx3_ASAP7_75t_SL _23339_ (.A(_15048_),
    .Y(_15049_));
 NOR2x1_ASAP7_75t_SL _23340_ (.A(_15046_),
    .B(_15049_),
    .Y(_15050_));
 AOI21x1_ASAP7_75t_SL _23341_ (.A1(_15043_),
    .A2(_15050_),
    .B(_15002_),
    .Y(_15051_));
 NAND2x2_ASAP7_75t_SL _23342_ (.A(_01193_),
    .B(_14937_),
    .Y(_15052_));
 INVx3_ASAP7_75t_SL _23343_ (.A(_15052_),
    .Y(_15053_));
 AOI21x1_ASAP7_75t_SL _23345_ (.A1(_14903_),
    .A2(_01193_),
    .B(_14937_),
    .Y(_15055_));
 OAI21x1_ASAP7_75t_SL _23347_ (.A1(_15053_),
    .A2(_15055_),
    .B(_14956_),
    .Y(_15057_));
 INVx1_ASAP7_75t_SL _23348_ (.A(_15042_),
    .Y(_15058_));
 OA21x2_ASAP7_75t_SL _23349_ (.A1(_15058_),
    .A2(_14956_),
    .B(_14975_),
    .Y(_15059_));
 NAND2x1_ASAP7_75t_SL _23350_ (.A(_15057_),
    .B(_15059_),
    .Y(_15060_));
 NAND2x1_ASAP7_75t_SL _23351_ (.A(_15051_),
    .B(_15060_),
    .Y(_15061_));
 AO21x1_ASAP7_75t_SL _23352_ (.A1(_14955_),
    .A2(_14950_),
    .B(_01202_),
    .Y(_15062_));
 INVx1_ASAP7_75t_SL _23354_ (.A(_01189_),
    .Y(_15064_));
 OAI21x1_ASAP7_75t_SL _23355_ (.A1(_14940_),
    .A2(_14941_),
    .B(_15064_),
    .Y(_15065_));
 INVx2_ASAP7_75t_SL _23356_ (.A(_15065_),
    .Y(_15066_));
 AOI21x1_ASAP7_75t_SL _23357_ (.A1(_15066_),
    .A2(_14982_),
    .B(_14975_),
    .Y(_15067_));
 AOI21x1_ASAP7_75t_SL _23358_ (.A1(_15067_),
    .A2(_15062_),
    .B(_15003_),
    .Y(_15068_));
 NOR2x1_ASAP7_75t_SL _23359_ (.A(_14937_),
    .B(_14978_),
    .Y(_15069_));
 OAI21x1_ASAP7_75t_SL _23361_ (.A1(_15042_),
    .A2(_15069_),
    .B(_14982_),
    .Y(_15071_));
 OAI21x1_ASAP7_75t_SL _23363_ (.A1(_14930_),
    .A2(_14936_),
    .B(_01188_),
    .Y(_15073_));
 NAND2x1_ASAP7_75t_SL _23364_ (.A(_15073_),
    .B(_15052_),
    .Y(_15074_));
 OAI21x1_ASAP7_75t_R _23365_ (.A1(_14940_),
    .A2(_14941_),
    .B(_14959_),
    .Y(_15075_));
 OAI21x1_ASAP7_75t_SL _23366_ (.A1(_15075_),
    .A2(_14956_),
    .B(_14975_),
    .Y(_15076_));
 AOI21x1_ASAP7_75t_SL _23367_ (.A1(_14956_),
    .A2(_15074_),
    .B(_15076_),
    .Y(_15077_));
 NAND2x1_ASAP7_75t_SL _23368_ (.A(_15071_),
    .B(_15077_),
    .Y(_15078_));
 AOI21x1_ASAP7_75t_SL _23370_ (.A1(_15078_),
    .A2(_15068_),
    .B(_15016_),
    .Y(_15080_));
 XNOR2x2_ASAP7_75t_R _23371_ (.A(_00598_),
    .B(_00629_),
    .Y(_15081_));
 XOR2x2_ASAP7_75t_R _23372_ (.A(_00661_),
    .B(_00662_),
    .Y(_15082_));
 XOR2x2_ASAP7_75t_R _23373_ (.A(_15082_),
    .B(_12268_),
    .Y(_15083_));
 XNOR2x2_ASAP7_75t_R _23374_ (.A(_15081_),
    .B(_15083_),
    .Y(_15084_));
 NOR2x1_ASAP7_75t_R _23375_ (.A(_00574_),
    .B(_00518_),
    .Y(_15085_));
 AO21x1_ASAP7_75t_SL _23376_ (.A1(_15084_),
    .A2(_00574_),
    .B(_15085_),
    .Y(_15086_));
 XOR2x2_ASAP7_75t_SL _23377_ (.A(_15086_),
    .B(_00917_),
    .Y(_15087_));
 AOI21x1_ASAP7_75t_SL _23379_ (.A1(_15080_),
    .A2(_15061_),
    .B(_15087_),
    .Y(_15089_));
 NAND2x1_ASAP7_75t_SL _23380_ (.A(_15089_),
    .B(_15040_),
    .Y(_15090_));
 NAND2x1_ASAP7_75t_SL _23381_ (.A(_14903_),
    .B(_01186_),
    .Y(_15091_));
 AO21x1_ASAP7_75t_SL _23382_ (.A1(_15052_),
    .A2(_15091_),
    .B(_14956_),
    .Y(_15092_));
 NAND2x1_ASAP7_75t_SL _23384_ (.A(_01187_),
    .B(_01186_),
    .Y(_15094_));
 AOI21x1_ASAP7_75t_SL _23385_ (.A1(_15094_),
    .A2(_15032_),
    .B(_14982_),
    .Y(_15095_));
 NOR2x1_ASAP7_75t_SL _23386_ (.A(_14975_),
    .B(_15095_),
    .Y(_15096_));
 NAND2x1_ASAP7_75t_SL _23387_ (.A(_15092_),
    .B(_15096_),
    .Y(_15097_));
 NOR2x1_ASAP7_75t_SL _23388_ (.A(_01187_),
    .B(_01186_),
    .Y(_15098_));
 NAND2x1_ASAP7_75t_SL _23389_ (.A(_14937_),
    .B(_15098_),
    .Y(_15099_));
 NAND2x1_ASAP7_75t_SL _23390_ (.A(_14982_),
    .B(_15047_),
    .Y(_15100_));
 INVx2_ASAP7_75t_SL _23391_ (.A(_15100_),
    .Y(_15101_));
 NAND2x1_ASAP7_75t_SL _23392_ (.A(_15099_),
    .B(_15101_),
    .Y(_15102_));
 INVx1_ASAP7_75t_SL _23394_ (.A(_01194_),
    .Y(_15104_));
 OAI21x1_ASAP7_75t_SL _23395_ (.A1(_15104_),
    .A2(_14937_),
    .B(_15023_),
    .Y(_15105_));
 AOI21x1_ASAP7_75t_SL _23397_ (.A1(_14956_),
    .A2(_15105_),
    .B(_15035_),
    .Y(_15107_));
 AOI21x1_ASAP7_75t_SL _23398_ (.A1(_15102_),
    .A2(_15107_),
    .B(_15017_),
    .Y(_15108_));
 NAND2x1_ASAP7_75t_SL _23399_ (.A(_15097_),
    .B(_15108_),
    .Y(_15109_));
 NAND2x2_ASAP7_75t_SL _23400_ (.A(_01187_),
    .B(_14937_),
    .Y(_15110_));
 AOI21x1_ASAP7_75t_SL _23402_ (.A1(_15047_),
    .A2(_15110_),
    .B(_14956_),
    .Y(_15112_));
 AO21x1_ASAP7_75t_SL _23403_ (.A1(_14956_),
    .A2(_15029_),
    .B(_14975_),
    .Y(_15113_));
 NOR2x1_ASAP7_75t_SL _23404_ (.A(_15112_),
    .B(_15113_),
    .Y(_15114_));
 OAI21x1_ASAP7_75t_SL _23405_ (.A1(_14930_),
    .A2(_14936_),
    .B(_15064_),
    .Y(_15115_));
 AO21x1_ASAP7_75t_SL _23406_ (.A1(_15023_),
    .A2(_15115_),
    .B(_14982_),
    .Y(_15116_));
 OAI21x1_ASAP7_75t_R _23407_ (.A1(_14920_),
    .A2(_14991_),
    .B(_00911_),
    .Y(_15117_));
 NAND3x1_ASAP7_75t_R _23408_ (.A(_14928_),
    .B(_14929_),
    .C(_14921_),
    .Y(_15118_));
 INVx1_ASAP7_75t_R _23409_ (.A(_01188_),
    .Y(_15119_));
 AOI21x1_ASAP7_75t_SL _23410_ (.A1(_15117_),
    .A2(_15118_),
    .B(_15119_),
    .Y(_15120_));
 NOR2x1_ASAP7_75t_SL _23411_ (.A(_15104_),
    .B(_14942_),
    .Y(_15121_));
 OAI21x1_ASAP7_75t_SL _23412_ (.A1(_15120_),
    .A2(_15121_),
    .B(_14982_),
    .Y(_15122_));
 AOI21x1_ASAP7_75t_SL _23413_ (.A1(_15116_),
    .A2(_15122_),
    .B(_15035_),
    .Y(_15123_));
 OAI21x1_ASAP7_75t_SL _23414_ (.A1(_15114_),
    .A2(_15123_),
    .B(_15017_),
    .Y(_15124_));
 NAND3x1_ASAP7_75t_SL _23416_ (.A(_15109_),
    .B(_15124_),
    .C(_15002_),
    .Y(_15126_));
 OAI21x1_ASAP7_75t_R _23417_ (.A1(_14903_),
    .A2(_14942_),
    .B(_01186_),
    .Y(_15127_));
 NAND2x1_ASAP7_75t_SL _23418_ (.A(_14982_),
    .B(_15127_),
    .Y(_15128_));
 INVx2_ASAP7_75t_SL _23419_ (.A(_01197_),
    .Y(_15129_));
 NOR2x1_ASAP7_75t_SL _23420_ (.A(_15129_),
    .B(_14942_),
    .Y(_15130_));
 INVx1_ASAP7_75t_SL _23421_ (.A(_15130_),
    .Y(_15131_));
 AOI21x1_ASAP7_75t_SL _23423_ (.A1(_15131_),
    .A2(_15049_),
    .B(_14975_),
    .Y(_15133_));
 NAND2x1_ASAP7_75t_SL _23424_ (.A(_15128_),
    .B(_15133_),
    .Y(_15134_));
 NAND2x1_ASAP7_75t_SL _23426_ (.A(_01186_),
    .B(_14937_),
    .Y(_15136_));
 AOI21x1_ASAP7_75t_SL _23428_ (.A1(_14982_),
    .A2(_15136_),
    .B(_15035_),
    .Y(_15138_));
 NAND2x1_ASAP7_75t_SL _23429_ (.A(_14937_),
    .B(_14978_),
    .Y(_15139_));
 INVx2_ASAP7_75t_R _23430_ (.A(_15022_),
    .Y(_15140_));
 NAND2x1_ASAP7_75t_SL _23431_ (.A(_15139_),
    .B(_15140_),
    .Y(_15141_));
 AOI21x1_ASAP7_75t_SL _23433_ (.A1(_15138_),
    .A2(_15141_),
    .B(_15017_),
    .Y(_15143_));
 AOI21x1_ASAP7_75t_SL _23434_ (.A1(_15134_),
    .A2(_15143_),
    .B(_15002_),
    .Y(_15144_));
 AO21x1_ASAP7_75t_SL _23435_ (.A1(_15110_),
    .A2(_14960_),
    .B(_14956_),
    .Y(_15145_));
 NAND3x1_ASAP7_75t_SL _23436_ (.A(_15057_),
    .B(_15145_),
    .C(_14975_),
    .Y(_15146_));
 NOR2x2_ASAP7_75t_SL _23437_ (.A(_14903_),
    .B(_14937_),
    .Y(_15147_));
 NOR2x1_ASAP7_75t_SL _23438_ (.A(_14956_),
    .B(_15147_),
    .Y(_15148_));
 AOI21x1_ASAP7_75t_SL _23439_ (.A1(_15139_),
    .A2(_15148_),
    .B(_14975_),
    .Y(_15149_));
 NOR2x2_ASAP7_75t_SL _23440_ (.A(_01193_),
    .B(_14942_),
    .Y(_15150_));
 NOR2x1_ASAP7_75t_SL _23441_ (.A(_15129_),
    .B(_14937_),
    .Y(_15151_));
 OR3x1_ASAP7_75t_SL _23442_ (.A(_15150_),
    .B(_15151_),
    .C(_14982_),
    .Y(_15152_));
 AOI21x1_ASAP7_75t_SL _23444_ (.A1(_15149_),
    .A2(_15152_),
    .B(_15016_),
    .Y(_15154_));
 NAND2x1_ASAP7_75t_SL _23445_ (.A(_15146_),
    .B(_15154_),
    .Y(_15155_));
 INVx1_ASAP7_75t_SL _23446_ (.A(_15087_),
    .Y(_15156_));
 AOI21x1_ASAP7_75t_SL _23447_ (.A1(_15144_),
    .A2(_15155_),
    .B(_15156_),
    .Y(_15157_));
 NAND2x1_ASAP7_75t_SL _23448_ (.A(_15126_),
    .B(_15157_),
    .Y(_15158_));
 NAND2x1_ASAP7_75t_SL _23449_ (.A(_15158_),
    .B(_15090_),
    .Y(_00080_));
 NAND2x1_ASAP7_75t_SL _23450_ (.A(_15021_),
    .B(_14982_),
    .Y(_15159_));
 NOR2x1_ASAP7_75t_R _23451_ (.A(_15053_),
    .B(_15159_),
    .Y(_15160_));
 NOR2x1_ASAP7_75t_L _23452_ (.A(_15150_),
    .B(_15048_),
    .Y(_15161_));
 OAI21x1_ASAP7_75t_R _23454_ (.A1(_15160_),
    .A2(_15161_),
    .B(_15035_),
    .Y(_15163_));
 NAND2x1_ASAP7_75t_SL _23455_ (.A(_14937_),
    .B(_14956_),
    .Y(_15164_));
 NOR2x1_ASAP7_75t_SL _23456_ (.A(_14978_),
    .B(_15164_),
    .Y(_15165_));
 NOR2x2_ASAP7_75t_SL _23457_ (.A(_01187_),
    .B(_14937_),
    .Y(_15166_));
 NOR2x1_ASAP7_75t_SL _23458_ (.A(_14903_),
    .B(_01193_),
    .Y(_15167_));
 NOR3x1_ASAP7_75t_R _23460_ (.A(_15166_),
    .B(_15167_),
    .C(_14956_),
    .Y(_15169_));
 OAI21x1_ASAP7_75t_R _23462_ (.A1(_15165_),
    .A2(_15169_),
    .B(_14975_),
    .Y(_15171_));
 AOI21x1_ASAP7_75t_R _23464_ (.A1(_15163_),
    .A2(_15171_),
    .B(_15017_),
    .Y(_15173_));
 NAND2x1_ASAP7_75t_L _23465_ (.A(_15029_),
    .B(_14956_),
    .Y(_15174_));
 OAI21x1_ASAP7_75t_R _23467_ (.A1(_15151_),
    .A2(_15174_),
    .B(_14975_),
    .Y(_15176_));
 NAND2x1_ASAP7_75t_R _23468_ (.A(_14942_),
    .B(_15091_),
    .Y(_15177_));
 AOI21x1_ASAP7_75t_R _23469_ (.A1(_15058_),
    .A2(_15177_),
    .B(_14956_),
    .Y(_15178_));
 NOR2x1_ASAP7_75t_R _23470_ (.A(_15176_),
    .B(_15178_),
    .Y(_15179_));
 INVx1_ASAP7_75t_R _23471_ (.A(_15043_),
    .Y(_15180_));
 NAND2x1_ASAP7_75t_SL _23472_ (.A(_14903_),
    .B(_14937_),
    .Y(_15181_));
 AO21x1_ASAP7_75t_R _23473_ (.A1(_15181_),
    .A2(_14956_),
    .B(_15147_),
    .Y(_15182_));
 OAI21x1_ASAP7_75t_R _23474_ (.A1(_15180_),
    .A2(_15182_),
    .B(_15017_),
    .Y(_15183_));
 OAI21x1_ASAP7_75t_R _23475_ (.A1(_15179_),
    .A2(_15183_),
    .B(_15002_),
    .Y(_15184_));
 OAI21x1_ASAP7_75t_R _23476_ (.A1(_15173_),
    .A2(_15184_),
    .B(_15156_),
    .Y(_15185_));
 NAND3x1_ASAP7_75t_R _23478_ (.A(_15052_),
    .B(_14982_),
    .C(_15073_),
    .Y(_15187_));
 NAND2x1p5_ASAP7_75t_L _23479_ (.A(_15058_),
    .B(_15049_),
    .Y(_15188_));
 AOI21x1_ASAP7_75t_R _23480_ (.A1(_15187_),
    .A2(_15188_),
    .B(_14975_),
    .Y(_15189_));
 NOR2x2_ASAP7_75t_SL _23481_ (.A(_01193_),
    .B(_14937_),
    .Y(_15190_));
 NAND2x1p5_ASAP7_75t_SL _23482_ (.A(_14982_),
    .B(_15065_),
    .Y(_15191_));
 OAI21x1_ASAP7_75t_R _23483_ (.A1(_15190_),
    .A2(_15191_),
    .B(_14975_),
    .Y(_15192_));
 OA21x2_ASAP7_75t_R _23484_ (.A1(_15190_),
    .A2(_15098_),
    .B(_14956_),
    .Y(_15193_));
 OAI21x1_ASAP7_75t_SL _23485_ (.A1(_15193_),
    .A2(_15192_),
    .B(_15017_),
    .Y(_15194_));
 OAI21x1_ASAP7_75t_SL _23487_ (.A1(_15194_),
    .A2(_15189_),
    .B(_15003_),
    .Y(_15196_));
 NAND2x1_ASAP7_75t_R _23488_ (.A(_14982_),
    .B(_15055_),
    .Y(_15197_));
 NOR2x1_ASAP7_75t_R _23489_ (.A(_14982_),
    .B(_15130_),
    .Y(_15198_));
 AOI21x1_ASAP7_75t_SL _23490_ (.A1(_15028_),
    .A2(_15198_),
    .B(_14975_),
    .Y(_15199_));
 INVx1_ASAP7_75t_R _23491_ (.A(_01192_),
    .Y(_15200_));
 NAND2x1_ASAP7_75t_R _23492_ (.A(_15200_),
    .B(_14942_),
    .Y(_15201_));
 OAI21x1_ASAP7_75t_R _23493_ (.A1(_14956_),
    .A2(_15201_),
    .B(_14975_),
    .Y(_15202_));
 NAND2x2_ASAP7_75t_SL _23494_ (.A(_14903_),
    .B(_01193_),
    .Y(_15203_));
 NAND2x1_ASAP7_75t_R _23495_ (.A(_14937_),
    .B(_15203_),
    .Y(_15204_));
 AOI21x1_ASAP7_75t_R _23496_ (.A1(_15047_),
    .A2(_15204_),
    .B(_14982_),
    .Y(_15205_));
 OAI21x1_ASAP7_75t_R _23497_ (.A1(_15202_),
    .A2(_15205_),
    .B(_15016_),
    .Y(_15206_));
 AOI21x1_ASAP7_75t_R _23498_ (.A1(_15197_),
    .A2(_15199_),
    .B(_15206_),
    .Y(_15207_));
 NOR2x1_ASAP7_75t_L _23499_ (.A(_15207_),
    .B(_15196_),
    .Y(_15208_));
 NOR2x1_ASAP7_75t_R _23500_ (.A(_14903_),
    .B(_14942_),
    .Y(_15209_));
 OAI21x1_ASAP7_75t_R _23501_ (.A1(_15209_),
    .A2(_15022_),
    .B(_14975_),
    .Y(_15210_));
 NAND2x1_ASAP7_75t_SL _23502_ (.A(_15119_),
    .B(_14937_),
    .Y(_15211_));
 AND3x1_ASAP7_75t_R _23503_ (.A(_15032_),
    .B(_15211_),
    .C(_14982_),
    .Y(_15212_));
 OAI21x1_ASAP7_75t_R _23504_ (.A1(_15210_),
    .A2(_15212_),
    .B(_15016_),
    .Y(_15213_));
 NAND2x1_ASAP7_75t_R _23505_ (.A(_14960_),
    .B(_15052_),
    .Y(_15214_));
 NOR2x1_ASAP7_75t_R _23506_ (.A(_15073_),
    .B(_14982_),
    .Y(_15215_));
 AOI21x1_ASAP7_75t_R _23507_ (.A1(_14982_),
    .A2(_15214_),
    .B(_15215_),
    .Y(_15216_));
 OA21x2_ASAP7_75t_SL _23508_ (.A1(_15065_),
    .A2(_14982_),
    .B(_15035_),
    .Y(_15217_));
 AND2x2_ASAP7_75t_SL _23509_ (.A(_15216_),
    .B(_15217_),
    .Y(_15218_));
 NOR2x1_ASAP7_75t_SL _23510_ (.A(_15213_),
    .B(_15218_),
    .Y(_15219_));
 NAND2x1_ASAP7_75t_R _23511_ (.A(_14975_),
    .B(_15048_),
    .Y(_15220_));
 NOR2x1_ASAP7_75t_R _23512_ (.A(_14937_),
    .B(_15203_),
    .Y(_15221_));
 NAND2x1_ASAP7_75t_SL _23513_ (.A(_14982_),
    .B(_15136_),
    .Y(_15222_));
 NOR2x1_ASAP7_75t_R _23514_ (.A(_15221_),
    .B(_15222_),
    .Y(_15223_));
 OAI21x1_ASAP7_75t_SL _23515_ (.A1(_15220_),
    .A2(_15223_),
    .B(_15017_),
    .Y(_15224_));
 NOR2x1_ASAP7_75t_R _23516_ (.A(_14959_),
    .B(_14942_),
    .Y(_15225_));
 NAND2x1_ASAP7_75t_SL _23517_ (.A(_01197_),
    .B(_14942_),
    .Y(_15226_));
 NAND2x1_ASAP7_75t_L _23518_ (.A(_14982_),
    .B(_15226_),
    .Y(_15227_));
 OAI21x1_ASAP7_75t_R _23519_ (.A1(_15225_),
    .A2(_15227_),
    .B(_15035_),
    .Y(_15228_));
 NOR2x1_ASAP7_75t_R _23520_ (.A(_15205_),
    .B(_15228_),
    .Y(_15229_));
 OAI21x1_ASAP7_75t_R _23521_ (.A1(_15224_),
    .A2(_15229_),
    .B(_15003_),
    .Y(_15230_));
 OAI21x1_ASAP7_75t_SL _23522_ (.A1(_15230_),
    .A2(_15219_),
    .B(_15087_),
    .Y(_15231_));
 NOR2x1_ASAP7_75t_SL _23523_ (.A(_14956_),
    .B(_15190_),
    .Y(_15232_));
 AOI21x1_ASAP7_75t_R _23524_ (.A1(_15211_),
    .A2(_15232_),
    .B(_15017_),
    .Y(_15233_));
 NAND2x1_ASAP7_75t_SL _23525_ (.A(_14942_),
    .B(_15098_),
    .Y(_15234_));
 NAND3x1_ASAP7_75t_R _23526_ (.A(_15139_),
    .B(_15234_),
    .C(_14956_),
    .Y(_15235_));
 AOI21x1_ASAP7_75t_R _23527_ (.A1(_15233_),
    .A2(_15235_),
    .B(_14975_),
    .Y(_15236_));
 NAND2x1_ASAP7_75t_SL _23528_ (.A(_01186_),
    .B(_14942_),
    .Y(_15237_));
 AO21x1_ASAP7_75t_SL _23529_ (.A1(_15110_),
    .A2(_15237_),
    .B(_14956_),
    .Y(_15238_));
 NAND2x1_ASAP7_75t_SL _23530_ (.A(_15110_),
    .B(_15140_),
    .Y(_15239_));
 NAND3x1_ASAP7_75t_R _23531_ (.A(_15238_),
    .B(_15239_),
    .C(_15017_),
    .Y(_15240_));
 OAI21x1_ASAP7_75t_R _23532_ (.A1(_15014_),
    .A2(_15015_),
    .B(_01204_),
    .Y(_15241_));
 NOR2x1_ASAP7_75t_R _23533_ (.A(_14982_),
    .B(_15241_),
    .Y(_15242_));
 AOI21x1_ASAP7_75t_R _23534_ (.A1(_15234_),
    .A2(_14995_),
    .B(_15242_),
    .Y(_15243_));
 OAI21x1_ASAP7_75t_R _23535_ (.A1(_15035_),
    .A2(_15243_),
    .B(_15002_),
    .Y(_15244_));
 AOI21x1_ASAP7_75t_R _23536_ (.A1(_15236_),
    .A2(_15240_),
    .B(_15244_),
    .Y(_15245_));
 OAI22x1_ASAP7_75t_SL _23537_ (.A1(_15185_),
    .A2(_15208_),
    .B1(_15231_),
    .B2(_15245_),
    .Y(_00081_));
 AOI21x1_ASAP7_75t_R _23538_ (.A1(_15044_),
    .A2(_15110_),
    .B(_14982_),
    .Y(_15246_));
 NAND2x1_ASAP7_75t_SL _23539_ (.A(_15129_),
    .B(_14937_),
    .Y(_15247_));
 AOI21x1_ASAP7_75t_R _23540_ (.A1(_15247_),
    .A2(_15032_),
    .B(_14956_),
    .Y(_15248_));
 OAI21x1_ASAP7_75t_R _23541_ (.A1(_15246_),
    .A2(_15248_),
    .B(_15035_),
    .Y(_15249_));
 NOR2x1p5_ASAP7_75t_L _23542_ (.A(_15066_),
    .B(_15048_),
    .Y(_15250_));
 NOR2x1_ASAP7_75t_SL _23543_ (.A(_01186_),
    .B(_14937_),
    .Y(_15251_));
 NOR2x1_ASAP7_75t_SL _23544_ (.A(_01195_),
    .B(_14942_),
    .Y(_15252_));
 OA21x2_ASAP7_75t_SL _23545_ (.A1(_15251_),
    .A2(_15252_),
    .B(_14982_),
    .Y(_15253_));
 OAI21x1_ASAP7_75t_R _23546_ (.A1(_15253_),
    .A2(_15250_),
    .B(_14975_),
    .Y(_15254_));
 AOI21x1_ASAP7_75t_SL _23547_ (.A1(_15254_),
    .A2(_15249_),
    .B(_15017_),
    .Y(_15255_));
 AOI21x1_ASAP7_75t_R _23548_ (.A1(_15044_),
    .A2(_15247_),
    .B(_14956_),
    .Y(_15256_));
 AOI21x1_ASAP7_75t_R _23549_ (.A1(_15032_),
    .A2(_15058_),
    .B(_14982_),
    .Y(_15257_));
 OAI21x1_ASAP7_75t_R _23550_ (.A1(_15256_),
    .A2(_15257_),
    .B(_15035_),
    .Y(_15258_));
 AOI21x1_ASAP7_75t_R _23551_ (.A1(_15044_),
    .A2(_15058_),
    .B(_14956_),
    .Y(_15259_));
 NAND2x2_ASAP7_75t_SL _23552_ (.A(_14903_),
    .B(_14942_),
    .Y(_15260_));
 AOI21x1_ASAP7_75t_R _23553_ (.A1(_15260_),
    .A2(_15058_),
    .B(_14982_),
    .Y(_15261_));
 OAI21x1_ASAP7_75t_R _23554_ (.A1(_15259_),
    .A2(_15261_),
    .B(_14975_),
    .Y(_15262_));
 AOI21x1_ASAP7_75t_R _23555_ (.A1(_15258_),
    .A2(_15262_),
    .B(_15016_),
    .Y(_15263_));
 NOR3x1_ASAP7_75t_SL _23556_ (.A(_15255_),
    .B(_15263_),
    .C(_15002_),
    .Y(_15264_));
 INVx1_ASAP7_75t_R _23557_ (.A(_15159_),
    .Y(_15265_));
 NAND2x1_ASAP7_75t_SL _23558_ (.A(_15131_),
    .B(_15265_),
    .Y(_15266_));
 NAND3x1_ASAP7_75t_R _23559_ (.A(_15260_),
    .B(_15091_),
    .C(_14956_),
    .Y(_15267_));
 AO21x1_ASAP7_75t_R _23560_ (.A1(_15266_),
    .A2(_15267_),
    .B(_14975_),
    .Y(_15268_));
 AOI21x1_ASAP7_75t_SL _23561_ (.A1(_14942_),
    .A2(_15091_),
    .B(_15042_),
    .Y(_15269_));
 AOI21x1_ASAP7_75t_SL _23562_ (.A1(_14956_),
    .A2(_15269_),
    .B(_15035_),
    .Y(_15270_));
 NAND2x1_ASAP7_75t_SL _23563_ (.A(_15030_),
    .B(_15270_),
    .Y(_15271_));
 AOI21x1_ASAP7_75t_R _23564_ (.A1(_15268_),
    .A2(_15271_),
    .B(_15016_),
    .Y(_15272_));
 INVx2_ASAP7_75t_SL _23565_ (.A(_15115_),
    .Y(_15273_));
 NOR2x1p5_ASAP7_75t_SL _23566_ (.A(_14956_),
    .B(_15273_),
    .Y(_15274_));
 NAND2x1p5_ASAP7_75t_SL _23567_ (.A(_15274_),
    .B(_15110_),
    .Y(_15275_));
 INVx1_ASAP7_75t_R _23568_ (.A(_15075_),
    .Y(_15276_));
 OR3x1_ASAP7_75t_L _23569_ (.A(_15251_),
    .B(_15276_),
    .C(_14982_),
    .Y(_15277_));
 AOI21x1_ASAP7_75t_SL _23570_ (.A1(_15277_),
    .A2(_15275_),
    .B(_14975_),
    .Y(_15278_));
 OAI21x1_ASAP7_75t_SL _23571_ (.A1(_14942_),
    .A2(_15091_),
    .B(_14982_),
    .Y(_15279_));
 NAND2x1_ASAP7_75t_R _23572_ (.A(_14975_),
    .B(_15279_),
    .Y(_15280_));
 AO21x1_ASAP7_75t_SL _23573_ (.A1(_15098_),
    .A2(_14937_),
    .B(_14982_),
    .Y(_15281_));
 NOR2x1_ASAP7_75t_R _23574_ (.A(_15151_),
    .B(_15281_),
    .Y(_15282_));
 OAI21x1_ASAP7_75t_SL _23575_ (.A1(_15280_),
    .A2(_15282_),
    .B(_15016_),
    .Y(_15283_));
 OAI21x1_ASAP7_75t_SL _23576_ (.A1(_15283_),
    .A2(_15278_),
    .B(_15002_),
    .Y(_15284_));
 OAI21x1_ASAP7_75t_SL _23577_ (.A1(_15284_),
    .A2(_15272_),
    .B(_15087_),
    .Y(_15285_));
 NAND2x1_ASAP7_75t_R _23578_ (.A(_01204_),
    .B(_14982_),
    .Y(_15286_));
 NAND3x1_ASAP7_75t_L _23579_ (.A(_15260_),
    .B(_15094_),
    .C(_14956_),
    .Y(_15287_));
 AOI21x1_ASAP7_75t_R _23580_ (.A1(_15286_),
    .A2(_15287_),
    .B(_15035_),
    .Y(_15288_));
 NAND2x1_ASAP7_75t_SL _23581_ (.A(_01194_),
    .B(_14942_),
    .Y(_15289_));
 AO21x1_ASAP7_75t_SL _23582_ (.A1(_15065_),
    .A2(_15289_),
    .B(_14982_),
    .Y(_15290_));
 AO21x1_ASAP7_75t_R _23584_ (.A1(_15260_),
    .A2(_15023_),
    .B(_14956_),
    .Y(_15292_));
 AOI21x1_ASAP7_75t_SL _23585_ (.A1(_15292_),
    .A2(_15290_),
    .B(_14975_),
    .Y(_15293_));
 OAI21x1_ASAP7_75t_SL _23586_ (.A1(_15293_),
    .A2(_15288_),
    .B(_15017_),
    .Y(_15294_));
 OA21x2_ASAP7_75t_R _23587_ (.A1(_14956_),
    .A2(_01202_),
    .B(_14975_),
    .Y(_15295_));
 INVx1_ASAP7_75t_R _23588_ (.A(_15174_),
    .Y(_15296_));
 NAND2x1_ASAP7_75t_R _23589_ (.A(_14979_),
    .B(_15296_),
    .Y(_15297_));
 AOI21x1_ASAP7_75t_R _23590_ (.A1(_15295_),
    .A2(_15297_),
    .B(_15017_),
    .Y(_15298_));
 AO21x1_ASAP7_75t_SL _23591_ (.A1(_15181_),
    .A2(_15032_),
    .B(_14982_),
    .Y(_15299_));
 NOR2x1_ASAP7_75t_SL _23592_ (.A(_14956_),
    .B(_15166_),
    .Y(_15300_));
 AOI21x1_ASAP7_75t_SL _23593_ (.A1(_15300_),
    .A2(_15065_),
    .B(_14975_),
    .Y(_15301_));
 NAND2x1_ASAP7_75t_R _23594_ (.A(_15299_),
    .B(_15301_),
    .Y(_15302_));
 AOI21x1_ASAP7_75t_R _23595_ (.A1(_15298_),
    .A2(_15302_),
    .B(_15002_),
    .Y(_15303_));
 NAND2x1_ASAP7_75t_SL _23596_ (.A(_15303_),
    .B(_15294_),
    .Y(_15304_));
 NAND2x1_ASAP7_75t_SL _23597_ (.A(_01201_),
    .B(_14956_),
    .Y(_15305_));
 AOI21x1_ASAP7_75t_R _23598_ (.A1(_15305_),
    .A2(_15279_),
    .B(_15035_),
    .Y(_15306_));
 AO21x1_ASAP7_75t_R _23599_ (.A1(_14981_),
    .A2(_14980_),
    .B(_01206_),
    .Y(_15307_));
 AOI21x1_ASAP7_75t_R _23600_ (.A1(_15307_),
    .A2(_15267_),
    .B(_14975_),
    .Y(_15308_));
 OAI21x1_ASAP7_75t_R _23601_ (.A1(_15306_),
    .A2(_15308_),
    .B(_15017_),
    .Y(_15309_));
 OAI21x1_ASAP7_75t_R _23602_ (.A1(_15273_),
    .A2(_15042_),
    .B(_14956_),
    .Y(_15310_));
 NOR2x1_ASAP7_75t_SL _23603_ (.A(_15073_),
    .B(_14956_),
    .Y(_15311_));
 NOR2x1_ASAP7_75t_R _23604_ (.A(_15035_),
    .B(_15311_),
    .Y(_15312_));
 AOI21x1_ASAP7_75t_SL _23605_ (.A1(_15312_),
    .A2(_15310_),
    .B(_15017_),
    .Y(_15313_));
 AOI21x1_ASAP7_75t_R _23606_ (.A1(_14995_),
    .A2(_15234_),
    .B(_14975_),
    .Y(_15314_));
 AND2x2_ASAP7_75t_R _23607_ (.A(_01190_),
    .B(_01192_),
    .Y(_15315_));
 NOR2x2_ASAP7_75t_SL _23608_ (.A(_15315_),
    .B(_14937_),
    .Y(_15316_));
 NOR2x1_ASAP7_75t_SL _23609_ (.A(_14942_),
    .B(_15098_),
    .Y(_15317_));
 OAI21x1_ASAP7_75t_R _23610_ (.A1(_15316_),
    .A2(_15317_),
    .B(_14956_),
    .Y(_15318_));
 NAND2x1_ASAP7_75t_SL _23611_ (.A(_15314_),
    .B(_15318_),
    .Y(_15319_));
 AOI21x1_ASAP7_75t_R _23612_ (.A1(_15319_),
    .A2(_15313_),
    .B(_15003_),
    .Y(_15320_));
 AOI21x1_ASAP7_75t_SL _23613_ (.A1(_15320_),
    .A2(_15309_),
    .B(_15087_),
    .Y(_15321_));
 NAND2x1_ASAP7_75t_SL _23614_ (.A(_15304_),
    .B(_15321_),
    .Y(_15322_));
 OAI21x1_ASAP7_75t_SL _23615_ (.A1(_15264_),
    .A2(_15285_),
    .B(_15322_),
    .Y(_00082_));
 OAI21x1_ASAP7_75t_SL _23616_ (.A1(_15252_),
    .A2(_15316_),
    .B(_14956_),
    .Y(_15323_));
 NAND2x1_ASAP7_75t_SL _23617_ (.A(_14995_),
    .B(_15234_),
    .Y(_15324_));
 AOI21x1_ASAP7_75t_SL _23618_ (.A1(_15323_),
    .A2(_15324_),
    .B(_15035_),
    .Y(_15325_));
 NAND2x1_ASAP7_75t_SL _23619_ (.A(_14982_),
    .B(_15247_),
    .Y(_15326_));
 OAI21x1_ASAP7_75t_SL _23620_ (.A1(_15251_),
    .A2(_15326_),
    .B(_15035_),
    .Y(_15327_));
 NAND2x1_ASAP7_75t_SL _23621_ (.A(_15017_),
    .B(_15327_),
    .Y(_15328_));
 OAI21x1_ASAP7_75t_SL _23622_ (.A1(_15325_),
    .A2(_15328_),
    .B(_15003_),
    .Y(_15329_));
 NOR2x1_ASAP7_75t_SL _23623_ (.A(_15044_),
    .B(_14982_),
    .Y(_15330_));
 NOR2x1_ASAP7_75t_SL _23624_ (.A(_15330_),
    .B(_15101_),
    .Y(_15331_));
 OA21x2_ASAP7_75t_SL _23625_ (.A1(_15136_),
    .A2(_14982_),
    .B(_15035_),
    .Y(_15332_));
 OAI21x1_ASAP7_75t_SL _23626_ (.A1(_15130_),
    .A2(_15331_),
    .B(_15332_),
    .Y(_15333_));
 AO21x1_ASAP7_75t_SL _23627_ (.A1(_15052_),
    .A2(_15073_),
    .B(_14982_),
    .Y(_15334_));
 AOI21x1_ASAP7_75t_SL _23628_ (.A1(_15094_),
    .A2(_15300_),
    .B(_15035_),
    .Y(_15335_));
 NAND2x1_ASAP7_75t_SL _23629_ (.A(_15334_),
    .B(_15335_),
    .Y(_15336_));
 AOI21x1_ASAP7_75t_SL _23630_ (.A1(_15333_),
    .A2(_15336_),
    .B(_15017_),
    .Y(_15337_));
 NOR2x1_ASAP7_75t_SL _23631_ (.A(_15329_),
    .B(_15337_),
    .Y(_15338_));
 INVx1_ASAP7_75t_SL _23632_ (.A(_15047_),
    .Y(_15339_));
 NAND2x1_ASAP7_75t_SL _23633_ (.A(_14982_),
    .B(_15339_),
    .Y(_15340_));
 OAI21x1_ASAP7_75t_SL _23634_ (.A1(_15017_),
    .A2(_15340_),
    .B(_14990_),
    .Y(_15341_));
 INVx2_ASAP7_75t_R _23635_ (.A(_15029_),
    .Y(_15342_));
 NAND2x1_ASAP7_75t_SL _23636_ (.A(_14956_),
    .B(_15342_),
    .Y(_15343_));
 NAND2x1_ASAP7_75t_SL _23637_ (.A(_15260_),
    .B(_14995_),
    .Y(_15344_));
 AOI21x1_ASAP7_75t_SL _23639_ (.A1(_15343_),
    .A2(_15344_),
    .B(_15016_),
    .Y(_15346_));
 OAI21x1_ASAP7_75t_SL _23640_ (.A1(_15341_),
    .A2(_15346_),
    .B(_15002_),
    .Y(_15347_));
 INVx1_ASAP7_75t_SL _23641_ (.A(_15247_),
    .Y(_15348_));
 OAI21x1_ASAP7_75t_SL _23642_ (.A1(_15316_),
    .A2(_15348_),
    .B(_14956_),
    .Y(_15349_));
 AO21x1_ASAP7_75t_SL _23643_ (.A1(_15115_),
    .A2(_15052_),
    .B(_14956_),
    .Y(_15350_));
 AOI21x1_ASAP7_75t_SL _23644_ (.A1(_15349_),
    .A2(_15350_),
    .B(_15016_),
    .Y(_15351_));
 NOR2x1_ASAP7_75t_L _23645_ (.A(_14956_),
    .B(_14985_),
    .Y(_15352_));
 AOI21x1_ASAP7_75t_SL _23646_ (.A1(_15237_),
    .A2(_15352_),
    .B(_15330_),
    .Y(_15353_));
 OAI21x1_ASAP7_75t_SL _23647_ (.A1(_15017_),
    .A2(_15353_),
    .B(_14975_),
    .Y(_15354_));
 NOR2x1_ASAP7_75t_SL _23648_ (.A(_15351_),
    .B(_15354_),
    .Y(_15355_));
 OAI21x1_ASAP7_75t_SL _23649_ (.A1(_15347_),
    .A2(_15355_),
    .B(_15087_),
    .Y(_15356_));
 NOR2x1_ASAP7_75t_SL _23650_ (.A(_15338_),
    .B(_15356_),
    .Y(_15357_));
 OAI21x1_ASAP7_75t_SL _23651_ (.A1(_15120_),
    .A2(_15174_),
    .B(_15035_),
    .Y(_15358_));
 NAND2x1_ASAP7_75t_SL _23652_ (.A(_15289_),
    .B(_15052_),
    .Y(_15359_));
 NOR2x1_ASAP7_75t_SL _23653_ (.A(_14956_),
    .B(_15359_),
    .Y(_15360_));
 NOR2x1_ASAP7_75t_SL _23654_ (.A(_15358_),
    .B(_15360_),
    .Y(_15361_));
 NOR2x1_ASAP7_75t_SL _23655_ (.A(_01197_),
    .B(_14937_),
    .Y(_15362_));
 OAI21x1_ASAP7_75t_SL _23656_ (.A1(_15042_),
    .A2(_15362_),
    .B(_14956_),
    .Y(_15363_));
 AOI21x1_ASAP7_75t_SL _23657_ (.A1(_15363_),
    .A2(_15275_),
    .B(_15035_),
    .Y(_15364_));
 OAI21x1_ASAP7_75t_SL _23658_ (.A1(_15364_),
    .A2(_15361_),
    .B(_15016_),
    .Y(_15365_));
 AO21x1_ASAP7_75t_SL _23659_ (.A1(_15110_),
    .A2(_15232_),
    .B(_15113_),
    .Y(_15366_));
 AO21x1_ASAP7_75t_SL _23660_ (.A1(_15052_),
    .A2(_15094_),
    .B(_14956_),
    .Y(_15367_));
 AOI21x1_ASAP7_75t_SL _23661_ (.A1(_15049_),
    .A2(_15110_),
    .B(_15035_),
    .Y(_15368_));
 AOI21x1_ASAP7_75t_SL _23662_ (.A1(_15368_),
    .A2(_15367_),
    .B(_15016_),
    .Y(_15369_));
 NAND2x1_ASAP7_75t_SL _23663_ (.A(_15366_),
    .B(_15369_),
    .Y(_15370_));
 AOI21x1_ASAP7_75t_SL _23664_ (.A1(_15370_),
    .A2(_15365_),
    .B(_15003_),
    .Y(_15371_));
 OAI21x1_ASAP7_75t_SL _23665_ (.A1(_15055_),
    .A2(_15191_),
    .B(_14975_),
    .Y(_15372_));
 NAND2x1_ASAP7_75t_SL _23666_ (.A(_14956_),
    .B(_15110_),
    .Y(_15373_));
 NOR2x1_ASAP7_75t_SL _23667_ (.A(_15373_),
    .B(_15359_),
    .Y(_15374_));
 NOR2x1_ASAP7_75t_SL _23668_ (.A(_15372_),
    .B(_15374_),
    .Y(_15375_));
 OAI21x1_ASAP7_75t_SL _23669_ (.A1(_15121_),
    .A2(_15100_),
    .B(_15035_),
    .Y(_15376_));
 OAI21x1_ASAP7_75t_SL _23670_ (.A1(_15095_),
    .A2(_15376_),
    .B(_15016_),
    .Y(_15377_));
 OAI21x1_ASAP7_75t_SL _23671_ (.A1(_15375_),
    .A2(_15377_),
    .B(_15003_),
    .Y(_15378_));
 OAI21x1_ASAP7_75t_R _23672_ (.A1(_14903_),
    .A2(_01193_),
    .B(_14975_),
    .Y(_15379_));
 NOR2x1_ASAP7_75t_SL _23673_ (.A(_15053_),
    .B(_15379_),
    .Y(_15380_));
 OAI21x1_ASAP7_75t_SL _23674_ (.A1(_14937_),
    .A2(_14982_),
    .B(_15380_),
    .Y(_15381_));
 OR3x1_ASAP7_75t_SL _23675_ (.A(_14985_),
    .B(_14956_),
    .C(_15273_),
    .Y(_15382_));
 NAND2x1_ASAP7_75t_SL _23676_ (.A(_15382_),
    .B(_15199_),
    .Y(_15383_));
 AOI21x1_ASAP7_75t_SL _23677_ (.A1(_15381_),
    .A2(_15383_),
    .B(_15016_),
    .Y(_15384_));
 OAI21x1_ASAP7_75t_SL _23678_ (.A1(_15384_),
    .A2(_15378_),
    .B(_15156_),
    .Y(_15385_));
 NOR2x1_ASAP7_75t_SL _23679_ (.A(_15371_),
    .B(_15385_),
    .Y(_15386_));
 NOR2x1_ASAP7_75t_SL _23680_ (.A(_15357_),
    .B(_15386_),
    .Y(_00083_));
 AOI21x1_ASAP7_75t_SL _23681_ (.A1(_15287_),
    .A2(_15238_),
    .B(_15035_),
    .Y(_15387_));
 AO21x1_ASAP7_75t_SL _23682_ (.A1(_15260_),
    .A2(_15023_),
    .B(_14982_),
    .Y(_15388_));
 AO21x1_ASAP7_75t_SL _23683_ (.A1(_15110_),
    .A2(_15091_),
    .B(_14956_),
    .Y(_15389_));
 AOI21x1_ASAP7_75t_SL _23684_ (.A1(_15388_),
    .A2(_15389_),
    .B(_14975_),
    .Y(_15390_));
 OAI21x1_ASAP7_75t_SL _23685_ (.A1(_15387_),
    .A2(_15390_),
    .B(_15017_),
    .Y(_15391_));
 NAND2x1_ASAP7_75t_SL _23686_ (.A(_14960_),
    .B(_15035_),
    .Y(_15392_));
 OA21x2_ASAP7_75t_SL _23687_ (.A1(_14986_),
    .A2(_15392_),
    .B(_15016_),
    .Y(_15393_));
 NAND2x1_ASAP7_75t_SL _23688_ (.A(_14956_),
    .B(_15181_),
    .Y(_15394_));
 AOI21x1_ASAP7_75t_SL _23689_ (.A1(_15211_),
    .A2(_15232_),
    .B(_15035_),
    .Y(_15395_));
 OAI21x1_ASAP7_75t_SL _23690_ (.A1(_15190_),
    .A2(_15394_),
    .B(_15395_),
    .Y(_15396_));
 AOI21x1_ASAP7_75t_SL _23691_ (.A1(_15393_),
    .A2(_15396_),
    .B(_15002_),
    .Y(_15397_));
 NAND2x1_ASAP7_75t_SL _23692_ (.A(_15391_),
    .B(_15397_),
    .Y(_15398_));
 OA21x2_ASAP7_75t_SL _23693_ (.A1(_15065_),
    .A2(_14982_),
    .B(_15044_),
    .Y(_15399_));
 AOI21x1_ASAP7_75t_SL _23694_ (.A1(_15043_),
    .A2(_15399_),
    .B(_15017_),
    .Y(_15400_));
 OAI21x1_ASAP7_75t_SL _23695_ (.A1(_01197_),
    .A2(_14937_),
    .B(_15065_),
    .Y(_15401_));
 AOI21x1_ASAP7_75t_SL _23696_ (.A1(_14982_),
    .A2(_15401_),
    .B(_15035_),
    .Y(_15402_));
 NAND2x1_ASAP7_75t_SL _23697_ (.A(_14987_),
    .B(_15402_),
    .Y(_15403_));
 AOI21x1_ASAP7_75t_SL _23698_ (.A1(_15400_),
    .A2(_15403_),
    .B(_15003_),
    .Y(_15404_));
 AO21x1_ASAP7_75t_R _23699_ (.A1(_14956_),
    .A2(_15120_),
    .B(_15035_),
    .Y(_15405_));
 AND3x1_ASAP7_75t_R _23700_ (.A(_14956_),
    .B(_14903_),
    .C(_14937_),
    .Y(_15406_));
 NOR2x1_ASAP7_75t_SL _23701_ (.A(_15405_),
    .B(_15406_),
    .Y(_15407_));
 NAND2x1_ASAP7_75t_SL _23702_ (.A(_15071_),
    .B(_15407_),
    .Y(_15408_));
 INVx1_ASAP7_75t_R _23703_ (.A(_15181_),
    .Y(_15409_));
 OAI21x1_ASAP7_75t_SL _23704_ (.A1(_15409_),
    .A2(_15069_),
    .B(_14956_),
    .Y(_15410_));
 OA21x2_ASAP7_75t_SL _23705_ (.A1(_15159_),
    .A2(_15130_),
    .B(_15035_),
    .Y(_15411_));
 AOI21x1_ASAP7_75t_SL _23706_ (.A1(_15410_),
    .A2(_15411_),
    .B(_15016_),
    .Y(_15412_));
 NAND2x1_ASAP7_75t_SL _23707_ (.A(_15408_),
    .B(_15412_),
    .Y(_15413_));
 AOI21x1_ASAP7_75t_SL _23708_ (.A1(_15404_),
    .A2(_15413_),
    .B(_15087_),
    .Y(_15414_));
 NAND2x1_ASAP7_75t_SL _23709_ (.A(_15398_),
    .B(_15414_),
    .Y(_15415_));
 NOR2x1_ASAP7_75t_SL _23710_ (.A(_15066_),
    .B(_15159_),
    .Y(_15416_));
 NAND2x1_ASAP7_75t_SL _23711_ (.A(_14975_),
    .B(_15057_),
    .Y(_15417_));
 OA21x2_ASAP7_75t_SL _23712_ (.A1(_15225_),
    .A2(_14956_),
    .B(_15035_),
    .Y(_15418_));
 AOI21x1_ASAP7_75t_SL _23713_ (.A1(_15281_),
    .A2(_15418_),
    .B(_15017_),
    .Y(_15419_));
 OAI21x1_ASAP7_75t_SL _23714_ (.A1(_15416_),
    .A2(_15417_),
    .B(_15419_),
    .Y(_15420_));
 OA21x2_ASAP7_75t_SL _23715_ (.A1(_15110_),
    .A2(_14956_),
    .B(_15035_),
    .Y(_15421_));
 AOI21x1_ASAP7_75t_SL _23716_ (.A1(_15110_),
    .A2(_15140_),
    .B(_15311_),
    .Y(_15422_));
 NAND2x1_ASAP7_75t_SL _23717_ (.A(_15421_),
    .B(_15422_),
    .Y(_15423_));
 AND2x2_ASAP7_75t_SL _23718_ (.A(_15164_),
    .B(_14975_),
    .Y(_15424_));
 AO21x1_ASAP7_75t_SL _23719_ (.A1(_15237_),
    .A2(_15247_),
    .B(_14956_),
    .Y(_15425_));
 AOI21x1_ASAP7_75t_SL _23720_ (.A1(_15424_),
    .A2(_15425_),
    .B(_15016_),
    .Y(_15426_));
 AOI21x1_ASAP7_75t_SL _23721_ (.A1(_15423_),
    .A2(_15426_),
    .B(_15002_),
    .Y(_15427_));
 AOI21x1_ASAP7_75t_SL _23722_ (.A1(_15420_),
    .A2(_15427_),
    .B(_15156_),
    .Y(_15428_));
 OR3x1_ASAP7_75t_SL _23723_ (.A(_15190_),
    .B(_15252_),
    .C(_14982_),
    .Y(_15429_));
 AOI21x1_ASAP7_75t_SL _23724_ (.A1(_15389_),
    .A2(_15429_),
    .B(_14975_),
    .Y(_15430_));
 NOR2x1_ASAP7_75t_SL _23725_ (.A(_15035_),
    .B(_15095_),
    .Y(_15431_));
 AO21x1_ASAP7_75t_SL _23726_ (.A1(_15431_),
    .A2(_15025_),
    .B(_15016_),
    .Y(_15432_));
 AO21x1_ASAP7_75t_SL _23727_ (.A1(_14982_),
    .A2(_01196_),
    .B(_15035_),
    .Y(_15433_));
 NOR2x1_ASAP7_75t_SL _23728_ (.A(_14982_),
    .B(_15066_),
    .Y(_15434_));
 OA21x2_ASAP7_75t_SL _23729_ (.A1(_15433_),
    .A2(_15434_),
    .B(_15016_),
    .Y(_15435_));
 NAND2x1_ASAP7_75t_SL _23730_ (.A(_14982_),
    .B(_15069_),
    .Y(_15436_));
 OAI21x1_ASAP7_75t_SL _23731_ (.A1(_15252_),
    .A2(_15166_),
    .B(_14956_),
    .Y(_15437_));
 NAND3x1_ASAP7_75t_SL _23732_ (.A(_15436_),
    .B(_15035_),
    .C(_15437_),
    .Y(_15438_));
 AOI21x1_ASAP7_75t_SL _23733_ (.A1(_15435_),
    .A2(_15438_),
    .B(_15003_),
    .Y(_15439_));
 OAI21x1_ASAP7_75t_SL _23734_ (.A1(_15430_),
    .A2(_15432_),
    .B(_15439_),
    .Y(_15440_));
 NAND2x1_ASAP7_75t_SL _23735_ (.A(_15428_),
    .B(_15440_),
    .Y(_15441_));
 NAND2x1_ASAP7_75t_SL _23736_ (.A(_15415_),
    .B(_15441_),
    .Y(_00084_));
 NOR2x1_ASAP7_75t_SL _23737_ (.A(_14956_),
    .B(_15032_),
    .Y(_15442_));
 OAI21x1_ASAP7_75t_R _23738_ (.A1(_15348_),
    .A2(_15055_),
    .B(_14982_),
    .Y(_15443_));
 OA21x2_ASAP7_75t_R _23739_ (.A1(_15031_),
    .A2(_14982_),
    .B(_15035_),
    .Y(_15444_));
 AOI21x1_ASAP7_75t_R _23740_ (.A1(_15443_),
    .A2(_15444_),
    .B(_15016_),
    .Y(_15445_));
 OA21x2_ASAP7_75t_SL _23741_ (.A1(_15060_),
    .A2(_15442_),
    .B(_15445_),
    .Y(_15446_));
 OA21x2_ASAP7_75t_R _23742_ (.A1(_14982_),
    .A2(_01186_),
    .B(_14975_),
    .Y(_15447_));
 AO21x1_ASAP7_75t_R _23743_ (.A1(_15092_),
    .A2(_15447_),
    .B(_15017_),
    .Y(_15448_));
 NAND2x1_ASAP7_75t_SL _23744_ (.A(_15028_),
    .B(_15352_),
    .Y(_15449_));
 NAND2x1_ASAP7_75t_L _23745_ (.A(_15139_),
    .B(_15049_),
    .Y(_15450_));
 AND3x1_ASAP7_75t_SL _23746_ (.A(_15449_),
    .B(_15450_),
    .C(_15035_),
    .Y(_15451_));
 OAI21x1_ASAP7_75t_R _23747_ (.A1(_15448_),
    .A2(_15451_),
    .B(_15003_),
    .Y(_15452_));
 NAND2x1_ASAP7_75t_R _23748_ (.A(_15315_),
    .B(_14942_),
    .Y(_15453_));
 AOI21x1_ASAP7_75t_R _23749_ (.A1(_14956_),
    .A2(_15453_),
    .B(_15035_),
    .Y(_15454_));
 OAI21x1_ASAP7_75t_R _23750_ (.A1(_15279_),
    .A2(_15221_),
    .B(_15454_),
    .Y(_15455_));
 INVx1_ASAP7_75t_SL _23751_ (.A(_15198_),
    .Y(_15456_));
 AOI21x1_ASAP7_75t_R _23752_ (.A1(_15043_),
    .A2(_15456_),
    .B(_15017_),
    .Y(_15457_));
 AOI21x1_ASAP7_75t_R _23753_ (.A1(_15455_),
    .A2(_15457_),
    .B(_15003_),
    .Y(_15458_));
 NOR2x1_ASAP7_75t_R _23754_ (.A(_14994_),
    .B(_15048_),
    .Y(_15459_));
 AO21x1_ASAP7_75t_SL _23755_ (.A1(_15131_),
    .A2(_15274_),
    .B(_14975_),
    .Y(_15460_));
 OA21x2_ASAP7_75t_R _23756_ (.A1(_14982_),
    .A2(_15104_),
    .B(_14975_),
    .Y(_15461_));
 AO21x1_ASAP7_75t_R _23757_ (.A1(_15098_),
    .A2(_14942_),
    .B(_14956_),
    .Y(_15462_));
 AOI21x1_ASAP7_75t_R _23758_ (.A1(_15461_),
    .A2(_15462_),
    .B(_15016_),
    .Y(_15463_));
 OAI21x1_ASAP7_75t_SL _23759_ (.A1(_15460_),
    .A2(_15459_),
    .B(_15463_),
    .Y(_15464_));
 AOI21x1_ASAP7_75t_SL _23760_ (.A1(_15464_),
    .A2(_15458_),
    .B(_15156_),
    .Y(_15465_));
 OAI21x1_ASAP7_75t_SL _23761_ (.A1(_15446_),
    .A2(_15452_),
    .B(_15465_),
    .Y(_15466_));
 NOR2x1_ASAP7_75t_R _23762_ (.A(_14956_),
    .B(_15150_),
    .Y(_15467_));
 NOR2x1_ASAP7_75t_SL _23763_ (.A(_15121_),
    .B(_15055_),
    .Y(_15468_));
 AOI22x1_ASAP7_75t_SL _23764_ (.A1(_15203_),
    .A2(_15467_),
    .B1(_15468_),
    .B2(_14956_),
    .Y(_15469_));
 OA21x2_ASAP7_75t_R _23765_ (.A1(_14982_),
    .A2(_01187_),
    .B(_14975_),
    .Y(_15470_));
 AOI21x1_ASAP7_75t_R _23766_ (.A1(_15470_),
    .A2(_15389_),
    .B(_15003_),
    .Y(_15471_));
 OAI21x1_ASAP7_75t_SL _23767_ (.A1(_14975_),
    .A2(_15469_),
    .B(_15471_),
    .Y(_15472_));
 NAND2x1_ASAP7_75t_R _23768_ (.A(_01192_),
    .B(_14960_),
    .Y(_15473_));
 AOI21x1_ASAP7_75t_R _23769_ (.A1(_14956_),
    .A2(_15473_),
    .B(_14975_),
    .Y(_15474_));
 NAND2x1_ASAP7_75t_R _23770_ (.A(_14979_),
    .B(_15352_),
    .Y(_15475_));
 AOI21x1_ASAP7_75t_R _23771_ (.A1(_15474_),
    .A2(_15475_),
    .B(_15002_),
    .Y(_15476_));
 NAND2x1_ASAP7_75t_SL _23772_ (.A(_15131_),
    .B(_15140_),
    .Y(_15477_));
 NAND3x1_ASAP7_75t_R _23773_ (.A(_15145_),
    .B(_15477_),
    .C(_14975_),
    .Y(_15478_));
 AOI21x1_ASAP7_75t_R _23774_ (.A1(_15476_),
    .A2(_15478_),
    .B(_15017_),
    .Y(_15479_));
 NAND2x1_ASAP7_75t_R _23775_ (.A(_15472_),
    .B(_15479_),
    .Y(_15480_));
 AO21x1_ASAP7_75t_R _23776_ (.A1(_15028_),
    .A2(_15075_),
    .B(_14956_),
    .Y(_15481_));
 AOI21x1_ASAP7_75t_SL _23777_ (.A1(_15481_),
    .A2(_15217_),
    .B(_15003_),
    .Y(_15482_));
 NAND2x1p5_ASAP7_75t_SL _23778_ (.A(_15049_),
    .B(_15023_),
    .Y(_15483_));
 AO21x1_ASAP7_75t_SL _23779_ (.A1(_15326_),
    .A2(_15483_),
    .B(_15035_),
    .Y(_15484_));
 NAND2x1_ASAP7_75t_SL _23780_ (.A(_15484_),
    .B(_15482_),
    .Y(_15485_));
 AOI21x1_ASAP7_75t_SL _23781_ (.A1(_14956_),
    .A2(_15150_),
    .B(_15035_),
    .Y(_15486_));
 AOI21x1_ASAP7_75t_R _23782_ (.A1(_15486_),
    .A2(_15331_),
    .B(_15002_),
    .Y(_15487_));
 NOR2x1_ASAP7_75t_R _23783_ (.A(_14975_),
    .B(_15165_),
    .Y(_15488_));
 NAND2x1_ASAP7_75t_SL _23784_ (.A(_15159_),
    .B(_15488_),
    .Y(_15489_));
 AOI21x1_ASAP7_75t_R _23785_ (.A1(_15487_),
    .A2(_15489_),
    .B(_15016_),
    .Y(_15490_));
 AOI21x1_ASAP7_75t_SL _23786_ (.A1(_15490_),
    .A2(_15485_),
    .B(_15087_),
    .Y(_15491_));
 NAND2x1_ASAP7_75t_SL _23787_ (.A(_15491_),
    .B(_15480_),
    .Y(_15492_));
 NAND2x2_ASAP7_75t_SL _23788_ (.A(_15466_),
    .B(_15492_),
    .Y(_00085_));
 AOI21x1_ASAP7_75t_SL _23789_ (.A1(_14956_),
    .A2(_15181_),
    .B(_14975_),
    .Y(_15493_));
 AOI21x1_ASAP7_75t_SL _23790_ (.A1(_15128_),
    .A2(_15493_),
    .B(_15016_),
    .Y(_15494_));
 AOI21x1_ASAP7_75t_SL _23791_ (.A1(_14982_),
    .A2(_15273_),
    .B(_15330_),
    .Y(_15495_));
 NAND2x1_ASAP7_75t_SL _23792_ (.A(_15486_),
    .B(_15495_),
    .Y(_15496_));
 NAND2x1_ASAP7_75t_SL _23793_ (.A(_15494_),
    .B(_15496_),
    .Y(_15497_));
 NAND2x1_ASAP7_75t_SL _23794_ (.A(_14956_),
    .B(_15094_),
    .Y(_15498_));
 AOI21x1_ASAP7_75t_SL _23795_ (.A1(_15498_),
    .A2(_15227_),
    .B(_15053_),
    .Y(_15499_));
 NAND2x1_ASAP7_75t_SL _23796_ (.A(_01187_),
    .B(_14982_),
    .Y(_15500_));
 AOI21x1_ASAP7_75t_SL _23797_ (.A1(_15500_),
    .A2(_15380_),
    .B(_15017_),
    .Y(_15501_));
 OAI21x1_ASAP7_75t_SL _23798_ (.A1(_14975_),
    .A2(_15499_),
    .B(_15501_),
    .Y(_15502_));
 AOI21x1_ASAP7_75t_SL _23799_ (.A1(_15497_),
    .A2(_15502_),
    .B(_15002_),
    .Y(_15503_));
 OA21x2_ASAP7_75t_SL _23800_ (.A1(_15052_),
    .A2(_14956_),
    .B(_15035_),
    .Y(_15504_));
 OAI21x1_ASAP7_75t_SL _23801_ (.A1(_15273_),
    .A2(_15456_),
    .B(_15504_),
    .Y(_15505_));
 AOI21x1_ASAP7_75t_SL _23802_ (.A1(_01200_),
    .A2(_14956_),
    .B(_15035_),
    .Y(_15506_));
 AOI21x1_ASAP7_75t_SL _23803_ (.A1(_15506_),
    .A2(_15449_),
    .B(_15017_),
    .Y(_15507_));
 NAND2x1_ASAP7_75t_SL _23804_ (.A(_15505_),
    .B(_15507_),
    .Y(_15508_));
 INVx1_ASAP7_75t_SL _23805_ (.A(_14995_),
    .Y(_15509_));
 AOI21x1_ASAP7_75t_SL _23806_ (.A1(_15509_),
    .A2(_15437_),
    .B(_14975_),
    .Y(_15510_));
 OAI21x1_ASAP7_75t_SL _23807_ (.A1(_15510_),
    .A2(_15270_),
    .B(_15017_),
    .Y(_15511_));
 AOI21x1_ASAP7_75t_SL _23808_ (.A1(_15508_),
    .A2(_15511_),
    .B(_15003_),
    .Y(_15512_));
 OAI21x1_ASAP7_75t_SL _23809_ (.A1(_15503_),
    .A2(_15512_),
    .B(_15087_),
    .Y(_15513_));
 AND2x2_ASAP7_75t_SL _23810_ (.A(_01205_),
    .B(_01199_),
    .Y(_15514_));
 OA21x2_ASAP7_75t_SL _23811_ (.A1(_14956_),
    .A2(_15514_),
    .B(_14975_),
    .Y(_15515_));
 AO21x1_ASAP7_75t_SL _23812_ (.A1(_15028_),
    .A2(_15203_),
    .B(_14982_),
    .Y(_15516_));
 NAND2x1_ASAP7_75t_SL _23813_ (.A(_15515_),
    .B(_15516_),
    .Y(_15517_));
 NAND2x1_ASAP7_75t_SL _23814_ (.A(_15044_),
    .B(_15075_),
    .Y(_15518_));
 AO21x1_ASAP7_75t_SL _23815_ (.A1(_14982_),
    .A2(_15120_),
    .B(_14975_),
    .Y(_15519_));
 AO21x1_ASAP7_75t_SL _23816_ (.A1(_14956_),
    .A2(_15518_),
    .B(_15519_),
    .Y(_15520_));
 AOI21x1_ASAP7_75t_SL _23817_ (.A1(_15517_),
    .A2(_15520_),
    .B(_15017_),
    .Y(_15521_));
 NOR3x1_ASAP7_75t_SL _23818_ (.A(_15518_),
    .B(_14982_),
    .C(_15042_),
    .Y(_15522_));
 INVx1_ASAP7_75t_SL _23819_ (.A(_15442_),
    .Y(_15523_));
 NAND2x1_ASAP7_75t_SL _23820_ (.A(_15523_),
    .B(_15067_),
    .Y(_15524_));
 OAI21x1_ASAP7_75t_SL _23821_ (.A1(_15522_),
    .A2(_15524_),
    .B(_15017_),
    .Y(_15525_));
 NAND2x1_ASAP7_75t_SL _23822_ (.A(_14956_),
    .B(_15317_),
    .Y(_15526_));
 AOI21x1_ASAP7_75t_SL _23823_ (.A1(_15226_),
    .A2(_15352_),
    .B(_14989_),
    .Y(_15527_));
 AOI21x1_ASAP7_75t_SL _23824_ (.A1(_15526_),
    .A2(_15527_),
    .B(_15035_),
    .Y(_15528_));
 NOR2x1_ASAP7_75t_SL _23825_ (.A(_15525_),
    .B(_15528_),
    .Y(_15529_));
 OAI21x1_ASAP7_75t_SL _23826_ (.A1(_15529_),
    .A2(_15521_),
    .B(_15003_),
    .Y(_15530_));
 AO21x1_ASAP7_75t_SL _23827_ (.A1(_15339_),
    .A2(_14982_),
    .B(_14975_),
    .Y(_15531_));
 AOI21x1_ASAP7_75t_SL _23828_ (.A1(_15279_),
    .A2(_15305_),
    .B(_15531_),
    .Y(_15532_));
 AO21x1_ASAP7_75t_SL _23829_ (.A1(_15047_),
    .A2(_15075_),
    .B(_14956_),
    .Y(_15533_));
 NOR2x1_ASAP7_75t_SL _23830_ (.A(_14982_),
    .B(_15147_),
    .Y(_15534_));
 NAND2x1_ASAP7_75t_SL _23831_ (.A(_15139_),
    .B(_15534_),
    .Y(_15535_));
 AOI21x1_ASAP7_75t_SL _23832_ (.A1(_15533_),
    .A2(_15535_),
    .B(_15035_),
    .Y(_15536_));
 OAI21x1_ASAP7_75t_SL _23833_ (.A1(_15532_),
    .A2(_15536_),
    .B(_15016_),
    .Y(_15537_));
 OAI21x1_ASAP7_75t_SL _23834_ (.A1(_15342_),
    .A2(_15316_),
    .B(_14982_),
    .Y(_15538_));
 OAI21x1_ASAP7_75t_SL _23835_ (.A1(_15167_),
    .A2(_15251_),
    .B(_14956_),
    .Y(_15539_));
 NAND3x1_ASAP7_75t_SL _23836_ (.A(_15538_),
    .B(_15486_),
    .C(_15539_),
    .Y(_15540_));
 AO21x1_ASAP7_75t_SL _23837_ (.A1(_15032_),
    .A2(_14903_),
    .B(_14982_),
    .Y(_15541_));
 OA21x2_ASAP7_75t_SL _23838_ (.A1(_15031_),
    .A2(_14956_),
    .B(_15035_),
    .Y(_15542_));
 AOI21x1_ASAP7_75t_SL _23839_ (.A1(_15541_),
    .A2(_15542_),
    .B(_15016_),
    .Y(_15543_));
 AOI21x1_ASAP7_75t_SL _23840_ (.A1(_15540_),
    .A2(_15543_),
    .B(_15003_),
    .Y(_15544_));
 AOI21x1_ASAP7_75t_SL _23841_ (.A1(_15537_),
    .A2(_15544_),
    .B(_15087_),
    .Y(_15545_));
 NAND2x1_ASAP7_75t_SL _23842_ (.A(_15545_),
    .B(_15530_),
    .Y(_15546_));
 NAND2x1_ASAP7_75t_SL _23843_ (.A(_15513_),
    .B(_15546_),
    .Y(_00086_));
 NAND2x1_ASAP7_75t_SL _23844_ (.A(_14956_),
    .B(_15401_),
    .Y(_15547_));
 AOI21x1_ASAP7_75t_SL _23845_ (.A1(_15547_),
    .A2(_15350_),
    .B(_14975_),
    .Y(_15548_));
 NAND2x1_ASAP7_75t_SL _23846_ (.A(_15226_),
    .B(_15352_),
    .Y(_15549_));
 AOI21x1_ASAP7_75t_SL _23847_ (.A1(_15299_),
    .A2(_15549_),
    .B(_15035_),
    .Y(_15550_));
 OAI21x1_ASAP7_75t_SL _23848_ (.A1(_15548_),
    .A2(_15550_),
    .B(_15017_),
    .Y(_15551_));
 AOI21x1_ASAP7_75t_SL _23849_ (.A1(_14979_),
    .A2(_15467_),
    .B(_14975_),
    .Y(_15552_));
 AO21x1_ASAP7_75t_SL _23850_ (.A1(_15204_),
    .A2(_15073_),
    .B(_14982_),
    .Y(_15553_));
 NAND2x1_ASAP7_75t_SL _23851_ (.A(_15552_),
    .B(_15553_),
    .Y(_15554_));
 AND2x2_ASAP7_75t_SL _23852_ (.A(_15227_),
    .B(_14975_),
    .Y(_15555_));
 AOI21x1_ASAP7_75t_SL _23853_ (.A1(_15437_),
    .A2(_15555_),
    .B(_15017_),
    .Y(_15556_));
 AOI21x1_ASAP7_75t_SL _23854_ (.A1(_15554_),
    .A2(_15556_),
    .B(_15002_),
    .Y(_15557_));
 NAND2x1_ASAP7_75t_SL _23855_ (.A(_15551_),
    .B(_15557_),
    .Y(_15558_));
 NAND2x1_ASAP7_75t_SL _23856_ (.A(_14956_),
    .B(_15055_),
    .Y(_15559_));
 OA21x2_ASAP7_75t_SL _23857_ (.A1(_14956_),
    .A2(_15047_),
    .B(_14975_),
    .Y(_15560_));
 AOI21x1_ASAP7_75t_SL _23858_ (.A1(_15559_),
    .A2(_15560_),
    .B(_15016_),
    .Y(_15561_));
 NAND2x1_ASAP7_75t_SL _23859_ (.A(_15274_),
    .B(_15099_),
    .Y(_15562_));
 AOI21x1_ASAP7_75t_SL _23860_ (.A1(_14956_),
    .A2(_14979_),
    .B(_14975_),
    .Y(_15563_));
 NAND2x1_ASAP7_75t_SL _23861_ (.A(_15562_),
    .B(_15563_),
    .Y(_15564_));
 AOI21x1_ASAP7_75t_SL _23862_ (.A1(_15561_),
    .A2(_15564_),
    .B(_15003_),
    .Y(_15565_));
 NAND2x1_ASAP7_75t_R _23863_ (.A(_01186_),
    .B(_14982_),
    .Y(_15566_));
 OAI21x1_ASAP7_75t_SL _23864_ (.A1(_15190_),
    .A2(_15394_),
    .B(_15566_),
    .Y(_15567_));
 NOR2x1_ASAP7_75t_SL _23865_ (.A(_14975_),
    .B(_15567_),
    .Y(_15568_));
 NAND2x1_ASAP7_75t_SL _23866_ (.A(_15099_),
    .B(_15148_),
    .Y(_15569_));
 AOI21x1_ASAP7_75t_SL _23867_ (.A1(_15287_),
    .A2(_15569_),
    .B(_15035_),
    .Y(_15570_));
 OAI21x1_ASAP7_75t_SL _23868_ (.A1(_15568_),
    .A2(_15570_),
    .B(_15016_),
    .Y(_15571_));
 AOI21x1_ASAP7_75t_SL _23869_ (.A1(_15565_),
    .A2(_15571_),
    .B(_15156_),
    .Y(_15572_));
 NAND2x1_ASAP7_75t_SL _23870_ (.A(_15558_),
    .B(_15572_),
    .Y(_01548_));
 OA21x2_ASAP7_75t_SL _23871_ (.A1(_15174_),
    .A2(_15273_),
    .B(_15035_),
    .Y(_01549_));
 OAI21x1_ASAP7_75t_SL _23872_ (.A1(_15222_),
    .A2(_15147_),
    .B(_01549_),
    .Y(_01550_));
 NAND2x1_ASAP7_75t_SL _23873_ (.A(_14982_),
    .B(_15342_),
    .Y(_01551_));
 INVx1_ASAP7_75t_R _23874_ (.A(_01205_),
    .Y(_01552_));
 AOI211x1_ASAP7_75t_SL _23875_ (.A1(_01552_),
    .A2(_14956_),
    .B(_15046_),
    .C(_15035_),
    .Y(_01553_));
 AOI21x1_ASAP7_75t_SL _23876_ (.A1(_01551_),
    .A2(_01553_),
    .B(_15016_),
    .Y(_01554_));
 NAND2x1_ASAP7_75t_SL _23877_ (.A(_01550_),
    .B(_01554_),
    .Y(_01555_));
 AND3x1_ASAP7_75t_SL _23878_ (.A(_14981_),
    .B(_01196_),
    .C(_14980_),
    .Y(_01556_));
 OA21x2_ASAP7_75t_SL _23879_ (.A1(_15076_),
    .A2(_01556_),
    .B(_15016_),
    .Y(_01557_));
 AO21x1_ASAP7_75t_SL _23880_ (.A1(_15032_),
    .A2(_14903_),
    .B(_14956_),
    .Y(_01558_));
 NAND3x1_ASAP7_75t_SL _23881_ (.A(_01558_),
    .B(_15239_),
    .C(_15035_),
    .Y(_01559_));
 AOI21x1_ASAP7_75t_SL _23882_ (.A1(_01557_),
    .A2(_01559_),
    .B(_15003_),
    .Y(_01560_));
 NAND2x1_ASAP7_75t_SL _23883_ (.A(_01555_),
    .B(_01560_),
    .Y(_01561_));
 AO21x1_ASAP7_75t_SL _23884_ (.A1(_15110_),
    .A2(_15073_),
    .B(_14982_),
    .Y(_01562_));
 NOR2x1_ASAP7_75t_SL _23885_ (.A(_15311_),
    .B(_15076_),
    .Y(_01563_));
 NAND2x1_ASAP7_75t_SL _23886_ (.A(_01562_),
    .B(_01563_),
    .Y(_01564_));
 OA21x2_ASAP7_75t_SL _23887_ (.A1(_14956_),
    .A2(_01192_),
    .B(_15035_),
    .Y(_01565_));
 AOI21x1_ASAP7_75t_SL _23888_ (.A1(_01565_),
    .A2(_15516_),
    .B(_15016_),
    .Y(_01566_));
 AOI21x1_ASAP7_75t_SL _23889_ (.A1(_01564_),
    .A2(_01566_),
    .B(_15002_),
    .Y(_01567_));
 AO21x1_ASAP7_75t_SL _23890_ (.A1(_15136_),
    .A2(_14903_),
    .B(_14956_),
    .Y(_01568_));
 AOI21x1_ASAP7_75t_SL _23891_ (.A1(_15323_),
    .A2(_01568_),
    .B(_14975_),
    .Y(_01569_));
 NOR2x1_ASAP7_75t_SL _23892_ (.A(_15121_),
    .B(_15048_),
    .Y(_01570_));
 NAND2x1_ASAP7_75t_SL _23893_ (.A(_15073_),
    .B(_15110_),
    .Y(_01571_));
 OAI21x1_ASAP7_75t_SL _23894_ (.A1(_15222_),
    .A2(_01571_),
    .B(_14975_),
    .Y(_01572_));
 NOR2x1_ASAP7_75t_SL _23895_ (.A(_01570_),
    .B(_01572_),
    .Y(_01573_));
 OAI21x1_ASAP7_75t_SL _23896_ (.A1(_01569_),
    .A2(_01573_),
    .B(_15016_),
    .Y(_01574_));
 AOI21x1_ASAP7_75t_SL _23897_ (.A1(_01567_),
    .A2(_01574_),
    .B(_15087_),
    .Y(_01575_));
 NAND2x1_ASAP7_75t_SL _23898_ (.A(_01561_),
    .B(_01575_),
    .Y(_01576_));
 NAND2x1_ASAP7_75t_SL _23899_ (.A(_01548_),
    .B(_01576_),
    .Y(_00087_));
 NOR2x1_ASAP7_75t_R _23900_ (.A(_00574_),
    .B(_00465_),
    .Y(_01577_));
 INVx1_ASAP7_75t_R _23901_ (.A(_00600_),
    .Y(_01578_));
 XOR2x2_ASAP7_75t_R _23902_ (.A(_12766_),
    .B(_01578_),
    .Y(_01579_));
 XNOR2x2_ASAP7_75t_L _23903_ (.A(_00663_),
    .B(_00670_),
    .Y(_01580_));
 XOR2x1_ASAP7_75t_SL _23904_ (.A(_00664_),
    .Y(_01581_),
    .B(_00696_));
 XOR2x2_ASAP7_75t_SL _23905_ (.A(_01580_),
    .B(_01581_),
    .Y(_01582_));
 NAND2x1_ASAP7_75t_SL _23906_ (.A(_01579_),
    .B(_01582_),
    .Y(_01583_));
 XOR2x2_ASAP7_75t_R _23907_ (.A(_12766_),
    .B(_00600_),
    .Y(_01584_));
 XOR2x2_ASAP7_75t_SL _23908_ (.A(_00663_),
    .B(_00670_),
    .Y(_01585_));
 XOR2x2_ASAP7_75t_L _23909_ (.A(_01585_),
    .B(_01581_),
    .Y(_01586_));
 NAND2x1_ASAP7_75t_SL _23910_ (.A(_01584_),
    .B(_01586_),
    .Y(_01587_));
 AOI21x1_ASAP7_75t_SL _23911_ (.A1(_01583_),
    .A2(_01587_),
    .B(_10675_),
    .Y(_01588_));
 OAI21x1_ASAP7_75t_R _23912_ (.A1(_01577_),
    .A2(_01588_),
    .B(_00942_),
    .Y(_01589_));
 AND2x2_ASAP7_75t_R _23913_ (.A(_10675_),
    .B(_00465_),
    .Y(_01590_));
 NAND2x1_ASAP7_75t_L _23914_ (.A(_01584_),
    .B(_01582_),
    .Y(_01591_));
 NAND2x1_ASAP7_75t_L _23915_ (.A(_01579_),
    .B(_01586_),
    .Y(_01592_));
 AOI21x1_ASAP7_75t_SL _23916_ (.A1(_01591_),
    .A2(_01592_),
    .B(_10675_),
    .Y(_01593_));
 OAI21x1_ASAP7_75t_SL _23917_ (.A1(_01590_),
    .A2(_01593_),
    .B(_08047_),
    .Y(_01594_));
 NAND2x1p5_ASAP7_75t_SL _23918_ (.A(_01594_),
    .B(_01589_),
    .Y(_01595_));
 NOR2x1_ASAP7_75t_SL _23920_ (.A(_00574_),
    .B(_00466_),
    .Y(_01596_));
 INVx1_ASAP7_75t_SL _23921_ (.A(_01596_),
    .Y(_01597_));
 XOR2x2_ASAP7_75t_L _23922_ (.A(_00599_),
    .B(_00638_),
    .Y(_01598_));
 NAND2x1p5_ASAP7_75t_L _23923_ (.A(_01598_),
    .B(_12786_),
    .Y(_01599_));
 XNOR2x2_ASAP7_75t_L _23924_ (.A(_00599_),
    .B(_00638_),
    .Y(_01600_));
 NAND2x1_ASAP7_75t_L _23925_ (.A(_00695_),
    .B(_01600_),
    .Y(_01601_));
 AOI21x1_ASAP7_75t_SL _23926_ (.A1(_01601_),
    .A2(_01599_),
    .B(_01580_),
    .Y(_01602_));
 XOR2x2_ASAP7_75t_L _23927_ (.A(_00638_),
    .B(_00695_),
    .Y(_01603_));
 NAND2x1_ASAP7_75t_L _23928_ (.A(_00599_),
    .B(_01603_),
    .Y(_01604_));
 INVx1_ASAP7_75t_R _23929_ (.A(_00599_),
    .Y(_01605_));
 XNOR2x2_ASAP7_75t_L _23930_ (.A(_00638_),
    .B(_00695_),
    .Y(_01606_));
 NAND2x1_ASAP7_75t_L _23931_ (.A(_01605_),
    .B(_01606_),
    .Y(_01607_));
 AOI21x1_ASAP7_75t_SL _23932_ (.A1(_01607_),
    .A2(_01604_),
    .B(_01585_),
    .Y(_01608_));
 OAI21x1_ASAP7_75t_SL _23933_ (.A1(_01602_),
    .A2(_01608_),
    .B(_00574_),
    .Y(_01609_));
 NAND2x1_ASAP7_75t_SL _23934_ (.A(_01597_),
    .B(_01609_),
    .Y(_01610_));
 XOR2x2_ASAP7_75t_SL _23935_ (.A(_01610_),
    .B(_08040_),
    .Y(_01611_));
 OR2x2_ASAP7_75t_R _23937_ (.A(_00574_),
    .B(_00467_),
    .Y(_01612_));
 NAND2x1_ASAP7_75t_R _23938_ (.A(_00665_),
    .B(_00697_),
    .Y(_01613_));
 NOR2x1_ASAP7_75t_SL _23939_ (.A(_00665_),
    .B(_00697_),
    .Y(_01614_));
 INVx1_ASAP7_75t_SL _23940_ (.A(_01614_),
    .Y(_01615_));
 INVx1_ASAP7_75t_R _23941_ (.A(_00601_),
    .Y(_01616_));
 AOI21x1_ASAP7_75t_R _23942_ (.A1(_01613_),
    .A2(_01615_),
    .B(_01616_),
    .Y(_01617_));
 NOR2x1_ASAP7_75t_SL _23943_ (.A(_00601_),
    .B(_12809_),
    .Y(_01618_));
 OAI21x1_ASAP7_75t_SL _23944_ (.A1(_01617_),
    .A2(_01618_),
    .B(_12769_),
    .Y(_01619_));
 INVx1_ASAP7_75t_SL _23945_ (.A(_01619_),
    .Y(_01620_));
 NOR3x1_ASAP7_75t_R _23946_ (.A(_01618_),
    .B(_01617_),
    .C(_12769_),
    .Y(_01621_));
 OAI21x1_ASAP7_75t_SL _23947_ (.A1(_01620_),
    .A2(_01621_),
    .B(_00574_),
    .Y(_01622_));
 INVx1_ASAP7_75t_R _23948_ (.A(_00943_),
    .Y(_01623_));
 AOI21x1_ASAP7_75t_SL _23949_ (.A1(_01612_),
    .A2(_01622_),
    .B(_01623_),
    .Y(_01624_));
 NAND2x1_ASAP7_75t_R _23950_ (.A(_00467_),
    .B(_10675_),
    .Y(_01625_));
 NAND2x1_ASAP7_75t_R _23951_ (.A(_01616_),
    .B(_12813_),
    .Y(_01626_));
 AND2x2_ASAP7_75t_R _23952_ (.A(_00665_),
    .B(_00697_),
    .Y(_01627_));
 OAI21x1_ASAP7_75t_R _23953_ (.A1(_01614_),
    .A2(_01627_),
    .B(_00601_),
    .Y(_01628_));
 INVx1_ASAP7_75t_R _23954_ (.A(_12769_),
    .Y(_01629_));
 NAND3x1_ASAP7_75t_SL _23955_ (.A(_01626_),
    .B(_01628_),
    .C(_01629_),
    .Y(_01630_));
 NAND3x1_ASAP7_75t_SL _23956_ (.A(_01630_),
    .B(_00574_),
    .C(_01619_),
    .Y(_01631_));
 AOI21x1_ASAP7_75t_SL _23957_ (.A1(_01625_),
    .A2(_01631_),
    .B(_00943_),
    .Y(_01632_));
 NOR2x2_ASAP7_75t_SL _23958_ (.A(_01624_),
    .B(_01632_),
    .Y(_01633_));
 XOR2x2_ASAP7_75t_SL _23961_ (.A(_00941_),
    .B(_01610_),
    .Y(_01635_));
 AOI21x1_ASAP7_75t_SL _23963_ (.A1(_01612_),
    .A2(_01622_),
    .B(_00943_),
    .Y(_01636_));
 AOI21x1_ASAP7_75t_SL _23964_ (.A1(_01625_),
    .A2(_01631_),
    .B(_01623_),
    .Y(_01637_));
 NOR2x2_ASAP7_75t_SL _23965_ (.A(_01636_),
    .B(_01637_),
    .Y(_01638_));
 NOR2x1_ASAP7_75t_SL _23968_ (.A(_01611_),
    .B(_01595_),
    .Y(_01640_));
 INVx1_ASAP7_75t_SL _23969_ (.A(_01640_),
    .Y(_01641_));
 NAND2x1_ASAP7_75t_SL _23970_ (.A(_01638_),
    .B(_01611_),
    .Y(_01642_));
 NOR2x1_ASAP7_75t_R _23972_ (.A(_00574_),
    .B(_00544_),
    .Y(_01644_));
 XOR2x2_ASAP7_75t_R _23973_ (.A(_12831_),
    .B(_00602_),
    .Y(_01645_));
 XOR2x2_ASAP7_75t_L _23974_ (.A(_00665_),
    .B(_00670_),
    .Y(_01646_));
 XNOR2x2_ASAP7_75t_L _23975_ (.A(_01646_),
    .B(_12830_),
    .Y(_01647_));
 NAND2x1_ASAP7_75t_SL _23976_ (.A(_01645_),
    .B(_01647_),
    .Y(_01648_));
 INVx1_ASAP7_75t_R _23977_ (.A(_00602_),
    .Y(_01649_));
 XOR2x2_ASAP7_75t_R _23978_ (.A(_12831_),
    .B(_01649_),
    .Y(_01650_));
 XOR2x2_ASAP7_75t_L _23979_ (.A(_12830_),
    .B(_01646_),
    .Y(_01651_));
 NAND2x1_ASAP7_75t_R _23980_ (.A(_01650_),
    .B(_01651_),
    .Y(_01652_));
 AOI21x1_ASAP7_75t_R _23981_ (.A1(_01648_),
    .A2(_01652_),
    .B(_10675_),
    .Y(_01653_));
 OAI21x1_ASAP7_75t_SL _23982_ (.A1(_01644_),
    .A2(_01653_),
    .B(_08031_),
    .Y(_01654_));
 NOR2x1_ASAP7_75t_R _23983_ (.A(_01650_),
    .B(_01651_),
    .Y(_01655_));
 NOR2x1_ASAP7_75t_SL _23984_ (.A(_01645_),
    .B(_01647_),
    .Y(_01656_));
 OAI21x1_ASAP7_75t_SL _23985_ (.A1(_01655_),
    .A2(_01656_),
    .B(_00574_),
    .Y(_01657_));
 INVx1_ASAP7_75t_SL _23986_ (.A(_01644_),
    .Y(_01658_));
 NAND3x1_ASAP7_75t_SL _23987_ (.A(_01657_),
    .B(_00944_),
    .C(_01658_),
    .Y(_01659_));
 NAND2x1_ASAP7_75t_SL _23988_ (.A(_01654_),
    .B(_01659_),
    .Y(_01660_));
 AO21x1_ASAP7_75t_SL _23990_ (.A1(_01641_),
    .A2(_01642_),
    .B(_01660_),
    .Y(_01662_));
 AND2x2_ASAP7_75t_R _23991_ (.A(_10675_),
    .B(_00543_),
    .Y(_01663_));
 XOR2x2_ASAP7_75t_L _23992_ (.A(_00666_),
    .B(_00670_),
    .Y(_01664_));
 INVx1_ASAP7_75t_R _23993_ (.A(_00699_),
    .Y(_01665_));
 XOR2x2_ASAP7_75t_R _23994_ (.A(_01664_),
    .B(_01665_),
    .Y(_01666_));
 XOR2x2_ASAP7_75t_L _23995_ (.A(_00634_),
    .B(_00638_),
    .Y(_01667_));
 XOR2x2_ASAP7_75t_L _23996_ (.A(_00603_),
    .B(_00667_),
    .Y(_01668_));
 XOR2x2_ASAP7_75t_R _23997_ (.A(_01667_),
    .B(_01668_),
    .Y(_01669_));
 NAND2x1_ASAP7_75t_SL _23998_ (.A(_01666_),
    .B(_01669_),
    .Y(_01670_));
 XOR2x2_ASAP7_75t_R _23999_ (.A(_01664_),
    .B(_00699_),
    .Y(_01671_));
 XOR2x2_ASAP7_75t_R _24000_ (.A(_12847_),
    .B(_01668_),
    .Y(_01672_));
 NAND2x1_ASAP7_75t_R _24001_ (.A(_01671_),
    .B(_01672_),
    .Y(_01673_));
 AOI21x1_ASAP7_75t_R _24002_ (.A1(_01670_),
    .A2(_01673_),
    .B(_10675_),
    .Y(_01674_));
 OAI21x1_ASAP7_75t_SL _24003_ (.A1(_01663_),
    .A2(_01674_),
    .B(_00946_),
    .Y(_01675_));
 NOR2x1_ASAP7_75t_R _24004_ (.A(_00574_),
    .B(_00543_),
    .Y(_01676_));
 XOR2x2_ASAP7_75t_R _24005_ (.A(_01667_),
    .B(_00603_),
    .Y(_01677_));
 XOR2x2_ASAP7_75t_R _24006_ (.A(_12848_),
    .B(_01664_),
    .Y(_01678_));
 NAND2x1_ASAP7_75t_SL _24007_ (.A(_01677_),
    .B(_01678_),
    .Y(_01679_));
 XNOR2x2_ASAP7_75t_R _24008_ (.A(_00603_),
    .B(_01667_),
    .Y(_01680_));
 XNOR2x2_ASAP7_75t_R _24009_ (.A(_12848_),
    .B(_01664_),
    .Y(_01681_));
 NAND2x1_ASAP7_75t_R _24010_ (.A(_01680_),
    .B(_01681_),
    .Y(_01682_));
 AOI21x1_ASAP7_75t_R _24011_ (.A1(_01679_),
    .A2(_01682_),
    .B(_10675_),
    .Y(_01683_));
 INVx1_ASAP7_75t_R _24012_ (.A(_00946_),
    .Y(_01684_));
 OAI21x1_ASAP7_75t_SL _24013_ (.A1(_01676_),
    .A2(_01683_),
    .B(_01684_),
    .Y(_01685_));
 NAND2x2_ASAP7_75t_SL _24014_ (.A(_01675_),
    .B(_01685_),
    .Y(_01686_));
 INVx2_ASAP7_75t_SL _24015_ (.A(_01686_),
    .Y(_01687_));
 NAND2x1_ASAP7_75t_SL _24018_ (.A(_01635_),
    .B(_01595_),
    .Y(_01690_));
 NAND2x1_ASAP7_75t_L _24019_ (.A(_01633_),
    .B(_01611_),
    .Y(_01691_));
 OAI21x1_ASAP7_75t_R _24020_ (.A1(_01644_),
    .A2(_01653_),
    .B(_00944_),
    .Y(_01692_));
 NAND3x1_ASAP7_75t_SL _24021_ (.A(_01657_),
    .B(_08031_),
    .C(_01658_),
    .Y(_01693_));
 NAND2x2_ASAP7_75t_SL _24022_ (.A(_01692_),
    .B(_01693_),
    .Y(_01694_));
 AO21x1_ASAP7_75t_SL _24024_ (.A1(_01690_),
    .A2(_01691_),
    .B(_01694_),
    .Y(_01696_));
 NAND3x1_ASAP7_75t_SL _24025_ (.A(_01662_),
    .B(_01687_),
    .C(_01696_),
    .Y(_01697_));
 OAI21x1_ASAP7_75t_SL _24026_ (.A1(_01624_),
    .A2(_01632_),
    .B(_01210_),
    .Y(_01698_));
 AND2x2_ASAP7_75t_SL _24028_ (.A(_01660_),
    .B(_01698_),
    .Y(_01700_));
 OAI21x1_ASAP7_75t_SL _24029_ (.A1(_01577_),
    .A2(_01588_),
    .B(_08047_),
    .Y(_01701_));
 OAI21x1_ASAP7_75t_SL _24030_ (.A1(_01590_),
    .A2(_01593_),
    .B(_00942_),
    .Y(_01702_));
 NAND2x2_ASAP7_75t_SL _24031_ (.A(_01702_),
    .B(_01701_),
    .Y(_01208_));
 NOR2x1_ASAP7_75t_SL _24032_ (.A(_01635_),
    .B(_01208_),
    .Y(_01703_));
 NAND2x1_ASAP7_75t_SL _24033_ (.A(_01633_),
    .B(_01703_),
    .Y(_01704_));
 NAND2x1_ASAP7_75t_SL _24034_ (.A(_01700_),
    .B(_01704_),
    .Y(_01705_));
 NAND2x1_ASAP7_75t_SL _24037_ (.A(_01209_),
    .B(_01633_),
    .Y(_01708_));
 NAND2x1_ASAP7_75t_SL _24038_ (.A(_01215_),
    .B(_01638_),
    .Y(_01709_));
 NAND2x1_ASAP7_75t_SL _24039_ (.A(_01708_),
    .B(_01709_),
    .Y(_01710_));
 AOI21x1_ASAP7_75t_SL _24040_ (.A1(_01694_),
    .A2(_01710_),
    .B(_01687_),
    .Y(_01711_));
 XOR2x2_ASAP7_75t_SL _24041_ (.A(_00667_),
    .B(_00668_),
    .Y(_01712_));
 INVx1_ASAP7_75t_R _24042_ (.A(_00700_),
    .Y(_01713_));
 XOR2x2_ASAP7_75t_R _24043_ (.A(_01712_),
    .B(_01713_),
    .Y(_01714_));
 XNOR2x2_ASAP7_75t_R _24044_ (.A(_00604_),
    .B(_00635_),
    .Y(_01715_));
 XOR2x2_ASAP7_75t_SL _24045_ (.A(_01714_),
    .B(_01715_),
    .Y(_01716_));
 NOR2x1_ASAP7_75t_R _24046_ (.A(_00574_),
    .B(_00542_),
    .Y(_01717_));
 INVx1_ASAP7_75t_R _24047_ (.A(_01717_),
    .Y(_01718_));
 OA21x2_ASAP7_75t_R _24048_ (.A1(_01716_),
    .A2(_10675_),
    .B(_01718_),
    .Y(_01719_));
 XOR2x2_ASAP7_75t_R _24049_ (.A(_01719_),
    .B(_08023_),
    .Y(_01720_));
 AOI21x1_ASAP7_75t_SL _24052_ (.A1(_01705_),
    .A2(_01711_),
    .B(_01720_),
    .Y(_01723_));
 INVx1_ASAP7_75t_SL _24053_ (.A(_01210_),
    .Y(_01724_));
 NOR2x1p5_ASAP7_75t_SL _24054_ (.A(_01638_),
    .B(_01724_),
    .Y(_01725_));
 AO21x1_ASAP7_75t_SL _24056_ (.A1(_01725_),
    .A2(_01694_),
    .B(_01686_),
    .Y(_01727_));
 NOR2x1p5_ASAP7_75t_SL _24058_ (.A(_01694_),
    .B(_01698_),
    .Y(_01729_));
 NAND2x2_ASAP7_75t_SL _24060_ (.A(_01633_),
    .B(_01208_),
    .Y(_01731_));
 NAND2x1_ASAP7_75t_SL _24061_ (.A(_01660_),
    .B(_01731_),
    .Y(_01732_));
 NOR2x1_ASAP7_75t_SL _24062_ (.A(_01729_),
    .B(_01732_),
    .Y(_01733_));
 OAI21x1_ASAP7_75t_SL _24063_ (.A1(_01727_),
    .A2(_01733_),
    .B(_01720_),
    .Y(_01734_));
 INVx1_ASAP7_75t_SL _24064_ (.A(_01209_),
    .Y(_01735_));
 NOR2x1_ASAP7_75t_R _24065_ (.A(_01735_),
    .B(_01633_),
    .Y(_01736_));
 NAND2x1_ASAP7_75t_SL _24066_ (.A(_01660_),
    .B(_01736_),
    .Y(_01737_));
 AND2x2_ASAP7_75t_SL _24068_ (.A(_01737_),
    .B(_01686_),
    .Y(_01739_));
 NAND2x1_ASAP7_75t_SL _24069_ (.A(_01735_),
    .B(_01633_),
    .Y(_01740_));
 NAND2x1p5_ASAP7_75t_SL _24070_ (.A(_01698_),
    .B(_01694_),
    .Y(_01741_));
 INVx3_ASAP7_75t_SL _24071_ (.A(_01741_),
    .Y(_01742_));
 OAI21x1_ASAP7_75t_R _24072_ (.A1(_01636_),
    .A2(_01637_),
    .B(_01215_),
    .Y(_01743_));
 NOR2x1_ASAP7_75t_SL _24073_ (.A(_01694_),
    .B(_01743_),
    .Y(_01744_));
 AOI21x1_ASAP7_75t_SL _24074_ (.A1(_01742_),
    .A2(_01740_),
    .B(_01744_),
    .Y(_01745_));
 AND2x2_ASAP7_75t_SL _24075_ (.A(_01739_),
    .B(_01745_),
    .Y(_01746_));
 NOR2x1_ASAP7_75t_SL _24076_ (.A(_01734_),
    .B(_01746_),
    .Y(_01747_));
 XOR2x2_ASAP7_75t_R _24077_ (.A(_00669_),
    .B(_00701_),
    .Y(_01748_));
 XOR2x2_ASAP7_75t_R _24078_ (.A(_12870_),
    .B(_00605_),
    .Y(_01749_));
 XNOR2x2_ASAP7_75t_R _24079_ (.A(_01748_),
    .B(_01749_),
    .Y(_01750_));
 NOR2x1_ASAP7_75t_R _24080_ (.A(_00574_),
    .B(_00541_),
    .Y(_01751_));
 AO21x1_ASAP7_75t_SL _24081_ (.A1(_01750_),
    .A2(_00574_),
    .B(_01751_),
    .Y(_01752_));
 XOR2x2_ASAP7_75t_SL _24082_ (.A(_01752_),
    .B(_00948_),
    .Y(_01753_));
 INVx1_ASAP7_75t_SL _24083_ (.A(_01753_),
    .Y(_01754_));
 AOI211x1_ASAP7_75t_SL _24085_ (.A1(_01697_),
    .A2(_01723_),
    .B(_01754_),
    .C(_01747_),
    .Y(_01756_));
 NOR2x1_ASAP7_75t_SL _24086_ (.A(_01638_),
    .B(_01635_),
    .Y(_01757_));
 AOI21x1_ASAP7_75t_SL _24087_ (.A1(_01611_),
    .A2(_01595_),
    .B(_01633_),
    .Y(_01758_));
 OAI21x1_ASAP7_75t_SL _24089_ (.A1(_01757_),
    .A2(_01758_),
    .B(_01694_),
    .Y(_01760_));
 INVx1_ASAP7_75t_SL _24090_ (.A(_01211_),
    .Y(_01761_));
 NAND2x1_ASAP7_75t_SL _24091_ (.A(_01761_),
    .B(_01638_),
    .Y(_01762_));
 AO21x1_ASAP7_75t_SL _24092_ (.A1(_01731_),
    .A2(_01762_),
    .B(_01694_),
    .Y(_01763_));
 NAND2x1_ASAP7_75t_SL _24093_ (.A(_01760_),
    .B(_01763_),
    .Y(_01764_));
 OAI21x1_ASAP7_75t_SL _24094_ (.A1(_01687_),
    .A2(_01764_),
    .B(_01720_),
    .Y(_01765_));
 NAND2x1_ASAP7_75t_R _24095_ (.A(_01208_),
    .B(_01660_),
    .Y(_01766_));
 NAND2x1_ASAP7_75t_SL _24096_ (.A(_01633_),
    .B(_01635_),
    .Y(_01767_));
 NAND2x1_ASAP7_75t_R _24097_ (.A(_01660_),
    .B(_01767_),
    .Y(_01768_));
 NAND2x1_ASAP7_75t_SL _24098_ (.A(_01766_),
    .B(_01768_),
    .Y(_01769_));
 NAND2x1_ASAP7_75t_SL _24099_ (.A(_01638_),
    .B(_01208_),
    .Y(_01770_));
 NAND2x1_ASAP7_75t_SL _24101_ (.A(_01218_),
    .B(_01638_),
    .Y(_01772_));
 AND3x1_ASAP7_75t_SL _24103_ (.A(_01767_),
    .B(_01772_),
    .C(_01694_),
    .Y(_01774_));
 AOI211x1_ASAP7_75t_SL _24104_ (.A1(_01769_),
    .A2(_01770_),
    .B(_01686_),
    .C(_01774_),
    .Y(_01775_));
 NOR2x1_ASAP7_75t_SL _24105_ (.A(_01765_),
    .B(_01775_),
    .Y(_01776_));
 INVx2_ASAP7_75t_R _24106_ (.A(_01213_),
    .Y(_01777_));
 NOR2x1_ASAP7_75t_SL _24107_ (.A(_01777_),
    .B(_01633_),
    .Y(_01778_));
 NOR2x1_ASAP7_75t_SL _24108_ (.A(_01660_),
    .B(_01778_),
    .Y(_01779_));
 NAND3x1_ASAP7_75t_SL _24109_ (.A(_01595_),
    .B(_01635_),
    .C(_01633_),
    .Y(_01780_));
 NOR2x1_ASAP7_75t_SL _24110_ (.A(_01638_),
    .B(_01611_),
    .Y(_01781_));
 NOR2x1_ASAP7_75t_L _24111_ (.A(_01694_),
    .B(_01781_),
    .Y(_01782_));
 AOI211x1_ASAP7_75t_SL _24112_ (.A1(_01779_),
    .A2(_01780_),
    .B(_01687_),
    .C(_01782_),
    .Y(_01783_));
 INVx1_ASAP7_75t_R _24113_ (.A(_01218_),
    .Y(_01784_));
 NOR2x1_ASAP7_75t_SL _24114_ (.A(_01784_),
    .B(_01638_),
    .Y(_01785_));
 OA21x2_ASAP7_75t_SL _24116_ (.A1(_01785_),
    .A2(_01741_),
    .B(_01687_),
    .Y(_01787_));
 OAI21x1_ASAP7_75t_SL _24119_ (.A1(_01638_),
    .A2(_01595_),
    .B(_01635_),
    .Y(_01790_));
 NAND2x1_ASAP7_75t_SL _24120_ (.A(_01660_),
    .B(_01790_),
    .Y(_01791_));
 AO21x1_ASAP7_75t_SL _24122_ (.A1(_01787_),
    .A2(_01791_),
    .B(_01720_),
    .Y(_01793_));
 OAI21x1_ASAP7_75t_SL _24123_ (.A1(_01783_),
    .A2(_01793_),
    .B(_01754_),
    .Y(_01794_));
 XOR2x2_ASAP7_75t_R _24124_ (.A(_00606_),
    .B(_00637_),
    .Y(_01795_));
 XOR2x2_ASAP7_75t_SL _24125_ (.A(_00569_),
    .B(_00669_),
    .Y(_01796_));
 XOR2x2_ASAP7_75t_R _24126_ (.A(_01796_),
    .B(_00670_),
    .Y(_01797_));
 XNOR2x2_ASAP7_75t_L _24127_ (.A(_01795_),
    .B(_01797_),
    .Y(_01798_));
 NOR2x1_ASAP7_75t_R _24128_ (.A(_00574_),
    .B(_00540_),
    .Y(_01799_));
 AO21x1_ASAP7_75t_SL _24129_ (.A1(_01798_),
    .A2(_00574_),
    .B(_01799_),
    .Y(_01800_));
 XOR2x2_ASAP7_75t_SL _24130_ (.A(_01800_),
    .B(_00949_),
    .Y(_01801_));
 OAI21x1_ASAP7_75t_SL _24132_ (.A1(_01794_),
    .A2(_01776_),
    .B(_01801_),
    .Y(_01803_));
 AO21x1_ASAP7_75t_SL _24134_ (.A1(_01762_),
    .A2(_01708_),
    .B(_01694_),
    .Y(_01805_));
 INVx1_ASAP7_75t_SL _24135_ (.A(_01779_),
    .Y(_01806_));
 AO21x1_ASAP7_75t_SL _24136_ (.A1(_01805_),
    .A2(_01806_),
    .B(_01686_),
    .Y(_01807_));
 NAND2x1p5_ASAP7_75t_SL _24137_ (.A(_01633_),
    .B(_01724_),
    .Y(_01808_));
 NOR2x1_ASAP7_75t_SL _24138_ (.A(_01633_),
    .B(_01208_),
    .Y(_01809_));
 NOR2x1_ASAP7_75t_SL _24139_ (.A(_01694_),
    .B(_01809_),
    .Y(_01810_));
 NAND2x1_ASAP7_75t_SL _24140_ (.A(_01808_),
    .B(_01810_),
    .Y(_01811_));
 AO21x1_ASAP7_75t_SL _24142_ (.A1(_01642_),
    .A2(_01743_),
    .B(_01660_),
    .Y(_01813_));
 AO21x1_ASAP7_75t_SL _24143_ (.A1(_01811_),
    .A2(_01813_),
    .B(_01687_),
    .Y(_01814_));
 AOI21x1_ASAP7_75t_SL _24145_ (.A1(_01807_),
    .A2(_01814_),
    .B(_01753_),
    .Y(_01816_));
 INVx1_ASAP7_75t_R _24146_ (.A(_01215_),
    .Y(_01817_));
 AOI21x1_ASAP7_75t_SL _24147_ (.A1(_01817_),
    .A2(_01633_),
    .B(_01694_),
    .Y(_01818_));
 NAND2x1_ASAP7_75t_SL _24148_ (.A(_01635_),
    .B(_01809_),
    .Y(_01819_));
 NAND2x1_ASAP7_75t_SL _24149_ (.A(_01818_),
    .B(_01819_),
    .Y(_01820_));
 NOR2x1_ASAP7_75t_SL _24151_ (.A(_01660_),
    .B(_01762_),
    .Y(_01822_));
 NOR2x1_ASAP7_75t_SL _24152_ (.A(_01686_),
    .B(_01822_),
    .Y(_01823_));
 AO21x1_ASAP7_75t_SL _24153_ (.A1(_01820_),
    .A2(_01823_),
    .B(_01754_),
    .Y(_01824_));
 NAND2x1_ASAP7_75t_SL _24154_ (.A(_01216_),
    .B(_01633_),
    .Y(_01825_));
 NAND3x1_ASAP7_75t_SL _24155_ (.A(_01819_),
    .B(_01694_),
    .C(_01825_),
    .Y(_01826_));
 OA21x2_ASAP7_75t_SL _24156_ (.A1(_01762_),
    .A2(_01694_),
    .B(_01686_),
    .Y(_01827_));
 AND2x2_ASAP7_75t_SL _24157_ (.A(_01826_),
    .B(_01827_),
    .Y(_01828_));
 XOR2x2_ASAP7_75t_SL _24158_ (.A(_01719_),
    .B(_00947_),
    .Y(_01829_));
 OAI21x1_ASAP7_75t_SL _24161_ (.A1(_01824_),
    .A2(_01828_),
    .B(_01829_),
    .Y(_01832_));
 AOI21x1_ASAP7_75t_SL _24162_ (.A1(_01694_),
    .A2(_01698_),
    .B(_01686_),
    .Y(_01833_));
 INVx1_ASAP7_75t_R _24163_ (.A(_01216_),
    .Y(_01834_));
 OAI21x1_ASAP7_75t_R _24164_ (.A1(_01624_),
    .A2(_01632_),
    .B(_01834_),
    .Y(_01835_));
 INVx2_ASAP7_75t_SL _24165_ (.A(_01835_),
    .Y(_01836_));
 NOR2x1_ASAP7_75t_SL _24166_ (.A(_01213_),
    .B(_01638_),
    .Y(_01837_));
 OAI21x1_ASAP7_75t_SL _24167_ (.A1(_01836_),
    .A2(_01837_),
    .B(_01660_),
    .Y(_01838_));
 AOI21x1_ASAP7_75t_SL _24168_ (.A1(_01833_),
    .A2(_01838_),
    .B(_01753_),
    .Y(_01839_));
 AOI21x1_ASAP7_75t_SL _24170_ (.A1(_01660_),
    .A2(_01837_),
    .B(_01687_),
    .Y(_01841_));
 NAND2x1_ASAP7_75t_SL _24171_ (.A(_01841_),
    .B(_01760_),
    .Y(_01842_));
 AOI21x1_ASAP7_75t_SL _24172_ (.A1(_01839_),
    .A2(_01842_),
    .B(_01829_),
    .Y(_01843_));
 AOI21x1_ASAP7_75t_SL _24173_ (.A1(_01635_),
    .A2(_01595_),
    .B(_01633_),
    .Y(_01844_));
 OAI21x1_ASAP7_75t_SL _24174_ (.A1(_01837_),
    .A2(_01844_),
    .B(_01660_),
    .Y(_01845_));
 INVx1_ASAP7_75t_SL _24175_ (.A(_01845_),
    .Y(_01846_));
 OAI21x1_ASAP7_75t_SL _24176_ (.A1(_01636_),
    .A2(_01637_),
    .B(_01761_),
    .Y(_01847_));
 NOR2x1_ASAP7_75t_SL _24177_ (.A(_01694_),
    .B(_01847_),
    .Y(_01848_));
 NOR2x1_ASAP7_75t_SL _24178_ (.A(_01687_),
    .B(_01848_),
    .Y(_01849_));
 NAND2x1_ASAP7_75t_SL _24179_ (.A(_01209_),
    .B(_01638_),
    .Y(_01850_));
 AO21x1_ASAP7_75t_SL _24180_ (.A1(_01691_),
    .A2(_01850_),
    .B(_01660_),
    .Y(_01851_));
 NAND2x1_ASAP7_75t_SL _24181_ (.A(_01849_),
    .B(_01851_),
    .Y(_01852_));
 AO21x1_ASAP7_75t_SL _24182_ (.A1(_01693_),
    .A2(_01692_),
    .B(_01223_),
    .Y(_01853_));
 NOR2x1_ASAP7_75t_SL _24183_ (.A(_01210_),
    .B(_01638_),
    .Y(_01854_));
 AOI21x1_ASAP7_75t_SL _24184_ (.A1(_01660_),
    .A2(_01854_),
    .B(_01686_),
    .Y(_01855_));
 AOI21x1_ASAP7_75t_SL _24185_ (.A1(_01853_),
    .A2(_01855_),
    .B(_01754_),
    .Y(_01856_));
 OAI21x1_ASAP7_75t_SL _24186_ (.A1(_01846_),
    .A2(_01852_),
    .B(_01856_),
    .Y(_01857_));
 AOI21x1_ASAP7_75t_SL _24187_ (.A1(_01843_),
    .A2(_01857_),
    .B(_01801_),
    .Y(_01858_));
 OAI21x1_ASAP7_75t_SL _24188_ (.A1(_01816_),
    .A2(_01832_),
    .B(_01858_),
    .Y(_01859_));
 OAI21x1_ASAP7_75t_SL _24189_ (.A1(_01756_),
    .A2(_01803_),
    .B(_01859_),
    .Y(_00088_));
 NAND2x1_ASAP7_75t_SL _24190_ (.A(_01660_),
    .B(_01758_),
    .Y(_01860_));
 NOR2x1_ASAP7_75t_SL _24191_ (.A(_01660_),
    .B(_01785_),
    .Y(_01861_));
 AOI21x1_ASAP7_75t_SL _24192_ (.A1(_01770_),
    .A2(_01861_),
    .B(_01686_),
    .Y(_01862_));
 NAND2x1_ASAP7_75t_SL _24193_ (.A(_01860_),
    .B(_01862_),
    .Y(_01863_));
 NAND2x1_ASAP7_75t_SL _24195_ (.A(_01777_),
    .B(_01638_),
    .Y(_01865_));
 OA21x2_ASAP7_75t_SL _24196_ (.A1(_01865_),
    .A2(_01694_),
    .B(_01686_),
    .Y(_01866_));
 INVx2_ASAP7_75t_SL _24197_ (.A(_01698_),
    .Y(_01867_));
 NOR2x1_ASAP7_75t_R _24198_ (.A(_01638_),
    .B(_01703_),
    .Y(_01868_));
 OAI21x1_ASAP7_75t_SL _24200_ (.A1(_01867_),
    .A2(_01868_),
    .B(_01694_),
    .Y(_01870_));
 AOI21x1_ASAP7_75t_SL _24201_ (.A1(_01866_),
    .A2(_01870_),
    .B(_01720_),
    .Y(_01871_));
 AOI21x1_ASAP7_75t_SL _24202_ (.A1(_01863_),
    .A2(_01871_),
    .B(_01801_),
    .Y(_01872_));
 NAND2x1_ASAP7_75t_R _24203_ (.A(_01611_),
    .B(_01595_),
    .Y(_01873_));
 NAND2x1_ASAP7_75t_SL _24204_ (.A(_01638_),
    .B(_01635_),
    .Y(_01874_));
 AO21x1_ASAP7_75t_SL _24205_ (.A1(_01873_),
    .A2(_01874_),
    .B(_01660_),
    .Y(_01875_));
 INVx2_ASAP7_75t_SL _24206_ (.A(_01725_),
    .Y(_01876_));
 AO21x1_ASAP7_75t_SL _24207_ (.A1(_01876_),
    .A2(_01642_),
    .B(_01694_),
    .Y(_01877_));
 AOI21x1_ASAP7_75t_SL _24208_ (.A1(_01875_),
    .A2(_01877_),
    .B(_01687_),
    .Y(_01878_));
 NAND2x1_ASAP7_75t_SL _24209_ (.A(_01777_),
    .B(_01633_),
    .Y(_01879_));
 NAND2x1_ASAP7_75t_SL _24210_ (.A(_01850_),
    .B(_01691_),
    .Y(_01880_));
 OAI21x1_ASAP7_75t_SL _24212_ (.A1(_01694_),
    .A2(_01880_),
    .B(_01687_),
    .Y(_01882_));
 AOI21x1_ASAP7_75t_SL _24213_ (.A1(_01879_),
    .A2(_01742_),
    .B(_01882_),
    .Y(_01883_));
 OAI21x1_ASAP7_75t_SL _24214_ (.A1(_01878_),
    .A2(_01883_),
    .B(_01720_),
    .Y(_01884_));
 NAND2x1_ASAP7_75t_SL _24215_ (.A(_01872_),
    .B(_01884_),
    .Y(_01885_));
 AO21x1_ASAP7_75t_SL _24216_ (.A1(_01850_),
    .A2(_01808_),
    .B(_01660_),
    .Y(_01886_));
 AO21x1_ASAP7_75t_SL _24218_ (.A1(_01691_),
    .A2(_01762_),
    .B(_01694_),
    .Y(_01888_));
 AOI21x1_ASAP7_75t_SL _24220_ (.A1(_01886_),
    .A2(_01888_),
    .B(_01686_),
    .Y(_01890_));
 AO21x1_ASAP7_75t_SL _24221_ (.A1(_01874_),
    .A2(_01708_),
    .B(_01694_),
    .Y(_01891_));
 NAND2x1_ASAP7_75t_SL _24222_ (.A(_01633_),
    .B(_01595_),
    .Y(_01892_));
 AO21x1_ASAP7_75t_SL _24223_ (.A1(_01892_),
    .A2(_01865_),
    .B(_01660_),
    .Y(_01893_));
 AOI21x1_ASAP7_75t_SL _24225_ (.A1(_01891_),
    .A2(_01893_),
    .B(_01687_),
    .Y(_01895_));
 OAI21x1_ASAP7_75t_SL _24226_ (.A1(_01890_),
    .A2(_01895_),
    .B(_01829_),
    .Y(_01896_));
 NAND2x1_ASAP7_75t_SL _24227_ (.A(_01784_),
    .B(_01638_),
    .Y(_01897_));
 NAND2x1_ASAP7_75t_SL _24228_ (.A(_01847_),
    .B(_01897_),
    .Y(_01898_));
 AOI21x1_ASAP7_75t_SL _24229_ (.A1(_01660_),
    .A2(_01898_),
    .B(_01686_),
    .Y(_01899_));
 NAND2x1_ASAP7_75t_SL _24230_ (.A(_01899_),
    .B(_01870_),
    .Y(_01900_));
 AND2x2_ASAP7_75t_SL _24231_ (.A(_01741_),
    .B(_01686_),
    .Y(_01901_));
 NOR2x1_ASAP7_75t_SL _24232_ (.A(_01633_),
    .B(_01635_),
    .Y(_01902_));
 NAND2x1_ASAP7_75t_SL _24233_ (.A(_01595_),
    .B(_01902_),
    .Y(_01903_));
 NAND2x1_ASAP7_75t_SL _24234_ (.A(_01903_),
    .B(_01782_),
    .Y(_01904_));
 AOI21x1_ASAP7_75t_SL _24236_ (.A1(_01901_),
    .A2(_01904_),
    .B(_01829_),
    .Y(_01906_));
 INVx1_ASAP7_75t_SL _24237_ (.A(_01801_),
    .Y(_01907_));
 AOI21x1_ASAP7_75t_SL _24238_ (.A1(_01900_),
    .A2(_01906_),
    .B(_01907_),
    .Y(_01908_));
 AOI21x1_ASAP7_75t_SL _24239_ (.A1(_01896_),
    .A2(_01908_),
    .B(_01753_),
    .Y(_01909_));
 NAND2x1_ASAP7_75t_SL _24240_ (.A(_01885_),
    .B(_01909_),
    .Y(_01910_));
 AOI21x1_ASAP7_75t_SL _24241_ (.A1(_01731_),
    .A2(_01779_),
    .B(_01686_),
    .Y(_01911_));
 NOR2x1_ASAP7_75t_R _24242_ (.A(_01694_),
    .B(_01902_),
    .Y(_01912_));
 AOI21x1_ASAP7_75t_SL _24243_ (.A1(_01892_),
    .A2(_01912_),
    .B(_01829_),
    .Y(_01913_));
 NAND2x1_ASAP7_75t_SL _24244_ (.A(_01911_),
    .B(_01913_),
    .Y(_01914_));
 NAND2x1_ASAP7_75t_SL _24245_ (.A(_01818_),
    .B(_01903_),
    .Y(_01915_));
 NAND2x1_ASAP7_75t_R _24246_ (.A(_01225_),
    .B(_01694_),
    .Y(_01916_));
 OA21x2_ASAP7_75t_SL _24247_ (.A1(_01916_),
    .A2(_01829_),
    .B(_01686_),
    .Y(_01917_));
 AOI21x1_ASAP7_75t_SL _24248_ (.A1(_01915_),
    .A2(_01917_),
    .B(_01907_),
    .Y(_01918_));
 NAND2x1_ASAP7_75t_SL _24249_ (.A(_01914_),
    .B(_01918_),
    .Y(_01919_));
 AO21x1_ASAP7_75t_SL _24250_ (.A1(_01642_),
    .A2(_01708_),
    .B(_01694_),
    .Y(_01920_));
 NAND2x1_ASAP7_75t_SL _24251_ (.A(_01687_),
    .B(_01829_),
    .Y(_01921_));
 INVx1_ASAP7_75t_SL _24252_ (.A(_01921_),
    .Y(_01922_));
 NOR2x1_ASAP7_75t_SL _24253_ (.A(_01638_),
    .B(_01660_),
    .Y(_01923_));
 NAND2x1_ASAP7_75t_SL _24254_ (.A(_01690_),
    .B(_01923_),
    .Y(_01924_));
 NAND2x1_ASAP7_75t_SL _24255_ (.A(_01694_),
    .B(_01758_),
    .Y(_01925_));
 AND4x1_ASAP7_75t_SL _24256_ (.A(_01920_),
    .B(_01922_),
    .C(_01924_),
    .D(_01925_),
    .Y(_01926_));
 NOR2x1_ASAP7_75t_SL _24257_ (.A(_01919_),
    .B(_01926_),
    .Y(_01927_));
 NOR2x1p5_ASAP7_75t_SL _24258_ (.A(_01660_),
    .B(_01725_),
    .Y(_01928_));
 AOI21x1_ASAP7_75t_SL _24259_ (.A1(_01772_),
    .A2(_01928_),
    .B(_01687_),
    .Y(_01929_));
 NAND2x1_ASAP7_75t_SL _24260_ (.A(_01845_),
    .B(_01929_),
    .Y(_01930_));
 INVx1_ASAP7_75t_SL _24261_ (.A(_01770_),
    .Y(_01931_));
 AOI21x1_ASAP7_75t_SL _24262_ (.A1(_01694_),
    .A2(_01892_),
    .B(_01931_),
    .Y(_01932_));
 OA21x2_ASAP7_75t_SL _24263_ (.A1(_01879_),
    .A2(_01694_),
    .B(_01687_),
    .Y(_01933_));
 AOI21x1_ASAP7_75t_SL _24264_ (.A1(_01932_),
    .A2(_01933_),
    .B(_01829_),
    .Y(_01934_));
 NAND2x1_ASAP7_75t_SL _24265_ (.A(_01930_),
    .B(_01934_),
    .Y(_01935_));
 NAND2x1p5_ASAP7_75t_SL _24266_ (.A(_01767_),
    .B(_01742_),
    .Y(_01936_));
 AO21x1_ASAP7_75t_SL _24267_ (.A1(_01767_),
    .A2(_01865_),
    .B(_01694_),
    .Y(_01937_));
 AOI21x1_ASAP7_75t_SL _24268_ (.A1(_01937_),
    .A2(_01936_),
    .B(_01921_),
    .Y(_01938_));
 NAND2x1_ASAP7_75t_SL _24269_ (.A(_01641_),
    .B(_01810_),
    .Y(_01939_));
 NAND2x1_ASAP7_75t_SL _24270_ (.A(_01686_),
    .B(_01829_),
    .Y(_01940_));
 AOI21x1_ASAP7_75t_SL _24271_ (.A1(_01924_),
    .A2(_01939_),
    .B(_01940_),
    .Y(_01941_));
 NOR2x1_ASAP7_75t_SL _24272_ (.A(_01938_),
    .B(_01941_),
    .Y(_01942_));
 AOI21x1_ASAP7_75t_SL _24273_ (.A1(_01935_),
    .A2(_01942_),
    .B(_01801_),
    .Y(_01943_));
 OAI21x1_ASAP7_75t_SL _24274_ (.A1(_01927_),
    .A2(_01943_),
    .B(_01753_),
    .Y(_01944_));
 NAND2x1_ASAP7_75t_SL _24275_ (.A(_01910_),
    .B(_01944_),
    .Y(_00089_));
 OAI21x1_ASAP7_75t_R _24276_ (.A1(_01837_),
    .A2(_01844_),
    .B(_01694_),
    .Y(_01945_));
 NAND2x1_ASAP7_75t_SL _24277_ (.A(_01638_),
    .B(_01595_),
    .Y(_01946_));
 AO21x1_ASAP7_75t_R _24278_ (.A1(_01946_),
    .A2(_01808_),
    .B(_01694_),
    .Y(_01947_));
 AOI21x1_ASAP7_75t_SL _24279_ (.A1(_01945_),
    .A2(_01947_),
    .B(_01687_),
    .Y(_01948_));
 NAND2x1_ASAP7_75t_SL _24280_ (.A(_01784_),
    .B(_01633_),
    .Y(_01949_));
 AO21x1_ASAP7_75t_SL _24281_ (.A1(_01949_),
    .A2(_01865_),
    .B(_01694_),
    .Y(_01950_));
 NOR2x1_ASAP7_75t_R _24282_ (.A(_01611_),
    .B(_01208_),
    .Y(_01951_));
 OR3x1_ASAP7_75t_SL _24283_ (.A(_01951_),
    .B(_01809_),
    .C(_01660_),
    .Y(_01952_));
 AOI21x1_ASAP7_75t_SL _24284_ (.A1(_01950_),
    .A2(_01952_),
    .B(_01686_),
    .Y(_01953_));
 OAI21x1_ASAP7_75t_SL _24285_ (.A1(_01948_),
    .A2(_01953_),
    .B(_01720_),
    .Y(_01954_));
 NAND2x1_ASAP7_75t_SL _24287_ (.A(_01660_),
    .B(_01780_),
    .Y(_01956_));
 AO21x1_ASAP7_75t_R _24288_ (.A1(_01595_),
    .A2(_01611_),
    .B(_01638_),
    .Y(_01957_));
 AO21x1_ASAP7_75t_SL _24289_ (.A1(_01957_),
    .A2(_01897_),
    .B(_01660_),
    .Y(_01958_));
 AOI21x1_ASAP7_75t_SL _24290_ (.A1(_01956_),
    .A2(_01958_),
    .B(_01940_),
    .Y(_01959_));
 AND3x1_ASAP7_75t_SL _24291_ (.A(_01642_),
    .B(_01694_),
    .C(_01847_),
    .Y(_01960_));
 NAND2x1_ASAP7_75t_SL _24292_ (.A(_01892_),
    .B(_01698_),
    .Y(_01961_));
 AO21x1_ASAP7_75t_SL _24293_ (.A1(_01961_),
    .A2(_01660_),
    .B(_01921_),
    .Y(_01962_));
 OAI21x1_ASAP7_75t_SL _24294_ (.A1(_01960_),
    .A2(_01962_),
    .B(_01753_),
    .Y(_01963_));
 NOR2x1_ASAP7_75t_SL _24295_ (.A(_01959_),
    .B(_01963_),
    .Y(_01964_));
 NAND2x1_ASAP7_75t_SL _24296_ (.A(_01954_),
    .B(_01964_),
    .Y(_01965_));
 NAND2x1p5_ASAP7_75t_SL _24297_ (.A(_01808_),
    .B(_01742_),
    .Y(_01966_));
 NAND2x1_ASAP7_75t_SL _24298_ (.A(_01834_),
    .B(_01633_),
    .Y(_01967_));
 AO21x1_ASAP7_75t_SL _24299_ (.A1(_01642_),
    .A2(_01967_),
    .B(_01694_),
    .Y(_01968_));
 AOI21x1_ASAP7_75t_SL _24300_ (.A1(_01968_),
    .A2(_01966_),
    .B(_01940_),
    .Y(_01969_));
 NAND2x1_ASAP7_75t_SL _24301_ (.A(_01660_),
    .B(_01949_),
    .Y(_01970_));
 OAI21x1_ASAP7_75t_SL _24302_ (.A1(_01902_),
    .A2(_01970_),
    .B(_01687_),
    .Y(_01971_));
 NAND2x1_ASAP7_75t_R _24303_ (.A(_01694_),
    .B(_01731_),
    .Y(_01972_));
 OAI21x1_ASAP7_75t_SL _24304_ (.A1(_01836_),
    .A2(_01972_),
    .B(_01829_),
    .Y(_01973_));
 OAI21x1_ASAP7_75t_SL _24305_ (.A1(_01971_),
    .A2(_01973_),
    .B(_01754_),
    .Y(_01974_));
 NOR2x1_ASAP7_75t_SL _24306_ (.A(_01969_),
    .B(_01974_),
    .Y(_01975_));
 AO21x1_ASAP7_75t_SL _24307_ (.A1(_01946_),
    .A2(_01879_),
    .B(_01660_),
    .Y(_01976_));
 AOI21x1_ASAP7_75t_SL _24308_ (.A1(_01838_),
    .A2(_01976_),
    .B(_01687_),
    .Y(_01977_));
 AO21x1_ASAP7_75t_SL _24309_ (.A1(_01949_),
    .A2(_01835_),
    .B(_01694_),
    .Y(_01978_));
 AO21x1_ASAP7_75t_SL _24310_ (.A1(_01642_),
    .A2(_01879_),
    .B(_01660_),
    .Y(_01979_));
 AOI21x1_ASAP7_75t_SL _24311_ (.A1(_01978_),
    .A2(_01979_),
    .B(_01686_),
    .Y(_01980_));
 OAI21x1_ASAP7_75t_SL _24312_ (.A1(_01977_),
    .A2(_01980_),
    .B(_01720_),
    .Y(_01981_));
 AOI21x1_ASAP7_75t_SL _24313_ (.A1(_01975_),
    .A2(_01981_),
    .B(_01907_),
    .Y(_01982_));
 NAND2x1_ASAP7_75t_SL _24314_ (.A(_01965_),
    .B(_01982_),
    .Y(_01983_));
 AND2x2_ASAP7_75t_L _24315_ (.A(_01211_),
    .B(_01213_),
    .Y(_01984_));
 NAND2x1_ASAP7_75t_SL _24316_ (.A(_01984_),
    .B(_01638_),
    .Y(_01985_));
 AND3x1_ASAP7_75t_SL _24317_ (.A(_01704_),
    .B(_01694_),
    .C(_01985_),
    .Y(_01986_));
 AO21x1_ASAP7_75t_SL _24318_ (.A1(_01903_),
    .A2(_01818_),
    .B(_01686_),
    .Y(_01987_));
 NAND2x1_ASAP7_75t_SL _24319_ (.A(_01213_),
    .B(_01633_),
    .Y(_01988_));
 NAND2x1_ASAP7_75t_SL _24320_ (.A(_01988_),
    .B(_01742_),
    .Y(_01989_));
 AOI21x1_ASAP7_75t_SL _24321_ (.A1(_01989_),
    .A2(_01739_),
    .B(_01720_),
    .Y(_01990_));
 OAI21x1_ASAP7_75t_SL _24322_ (.A1(_01986_),
    .A2(_01987_),
    .B(_01990_),
    .Y(_01991_));
 NAND2x1_ASAP7_75t_SL _24323_ (.A(_01222_),
    .B(_01694_),
    .Y(_01992_));
 NAND3x1_ASAP7_75t_SL _24324_ (.A(_01956_),
    .B(_01686_),
    .C(_01992_),
    .Y(_01993_));
 OA21x2_ASAP7_75t_SL _24325_ (.A1(_01694_),
    .A2(_01227_),
    .B(_01687_),
    .Y(_01994_));
 AOI21x1_ASAP7_75t_SL _24326_ (.A1(_01994_),
    .A2(_01952_),
    .B(_01829_),
    .Y(_01995_));
 AOI21x1_ASAP7_75t_SL _24327_ (.A1(_01993_),
    .A2(_01995_),
    .B(_01754_),
    .Y(_01996_));
 NAND2x1_ASAP7_75t_SL _24328_ (.A(_01991_),
    .B(_01996_),
    .Y(_01997_));
 AO21x1_ASAP7_75t_SL _24329_ (.A1(_01808_),
    .A2(_01709_),
    .B(_01660_),
    .Y(_01998_));
 AO21x1_ASAP7_75t_SL _24330_ (.A1(_01946_),
    .A2(_01708_),
    .B(_01694_),
    .Y(_01999_));
 AOI21x1_ASAP7_75t_SL _24331_ (.A1(_01998_),
    .A2(_01999_),
    .B(_01686_),
    .Y(_02000_));
 NAND2x1_ASAP7_75t_SL _24332_ (.A(_01225_),
    .B(_01660_),
    .Y(_02001_));
 NOR2x1_ASAP7_75t_R _24333_ (.A(_01660_),
    .B(_01640_),
    .Y(_02002_));
 NAND2x1_ASAP7_75t_SL _24334_ (.A(_01946_),
    .B(_02002_),
    .Y(_02003_));
 AOI21x1_ASAP7_75t_SL _24335_ (.A1(_02001_),
    .A2(_02003_),
    .B(_01687_),
    .Y(_02004_));
 OAI21x1_ASAP7_75t_SL _24336_ (.A1(_02000_),
    .A2(_02004_),
    .B(_01720_),
    .Y(_02005_));
 AO21x1_ASAP7_75t_SL _24337_ (.A1(_01892_),
    .A2(_01642_),
    .B(_01660_),
    .Y(_02006_));
 AOI21x1_ASAP7_75t_SL _24338_ (.A1(_01808_),
    .A2(_01810_),
    .B(_01686_),
    .Y(_02007_));
 NAND2x1_ASAP7_75t_SL _24339_ (.A(_02006_),
    .B(_02007_),
    .Y(_02008_));
 OA21x2_ASAP7_75t_SL _24340_ (.A1(_01694_),
    .A2(_01223_),
    .B(_01686_),
    .Y(_02009_));
 NAND2x1_ASAP7_75t_SL _24341_ (.A(_01928_),
    .B(_01819_),
    .Y(_02010_));
 AOI21x1_ASAP7_75t_SL _24342_ (.A1(_02009_),
    .A2(_02010_),
    .B(_01720_),
    .Y(_02011_));
 AOI21x1_ASAP7_75t_SL _24343_ (.A1(_02008_),
    .A2(_02011_),
    .B(_01753_),
    .Y(_02012_));
 AOI21x1_ASAP7_75t_SL _24344_ (.A1(_02005_),
    .A2(_02012_),
    .B(_01801_),
    .Y(_02013_));
 NAND2x1_ASAP7_75t_SL _24345_ (.A(_01997_),
    .B(_02013_),
    .Y(_02014_));
 NAND2x1_ASAP7_75t_SL _24346_ (.A(_01983_),
    .B(_02014_),
    .Y(_00090_));
 NAND2x1_ASAP7_75t_SL _24347_ (.A(_01638_),
    .B(_01694_),
    .Y(_02015_));
 OAI21x1_ASAP7_75t_R _24348_ (.A1(_01638_),
    .A2(_01635_),
    .B(_01686_),
    .Y(_02016_));
 NOR2x1_ASAP7_75t_SL _24349_ (.A(_01640_),
    .B(_02016_),
    .Y(_02017_));
 AOI21x1_ASAP7_75t_SL _24350_ (.A1(_02015_),
    .A2(_02017_),
    .B(_01829_),
    .Y(_02018_));
 AO21x1_ASAP7_75t_SL _24351_ (.A1(_01967_),
    .A2(_01698_),
    .B(_01694_),
    .Y(_02019_));
 NAND2x1_ASAP7_75t_SL _24352_ (.A(_02019_),
    .B(_01862_),
    .Y(_02020_));
 AOI21x1_ASAP7_75t_SL _24353_ (.A1(_02018_),
    .A2(_02020_),
    .B(_01801_),
    .Y(_02021_));
 NAND2x1_ASAP7_75t_R _24354_ (.A(_01709_),
    .B(_01691_),
    .Y(_02022_));
 NOR2x1_ASAP7_75t_SL _24355_ (.A(_01972_),
    .B(_02022_),
    .Y(_02023_));
 NAND2x1p5_ASAP7_75t_L _24356_ (.A(_01660_),
    .B(_01808_),
    .Y(_02024_));
 OAI21x1_ASAP7_75t_SL _24357_ (.A1(_01758_),
    .A2(_02024_),
    .B(_01686_),
    .Y(_02025_));
 NOR2x1_ASAP7_75t_SL _24358_ (.A(_02023_),
    .B(_02025_),
    .Y(_02026_));
 AO21x1_ASAP7_75t_SL _24359_ (.A1(_01743_),
    .A2(_01698_),
    .B(_01694_),
    .Y(_02027_));
 AO21x1_ASAP7_75t_SL _24360_ (.A1(_01690_),
    .A2(_01691_),
    .B(_01660_),
    .Y(_02028_));
 AOI21x1_ASAP7_75t_SL _24361_ (.A1(_02027_),
    .A2(_02028_),
    .B(_01686_),
    .Y(_02029_));
 OAI21x1_ASAP7_75t_SL _24362_ (.A1(_02026_),
    .A2(_02029_),
    .B(_01829_),
    .Y(_02030_));
 NAND2x1_ASAP7_75t_SL _24363_ (.A(_02021_),
    .B(_02030_),
    .Y(_02031_));
 NAND2x1_ASAP7_75t_SL _24364_ (.A(_01720_),
    .B(_01971_),
    .Y(_02032_));
 INVx1_ASAP7_75t_R _24365_ (.A(_01984_),
    .Y(_02033_));
 NAND2x1_ASAP7_75t_SL _24366_ (.A(_02033_),
    .B(_01638_),
    .Y(_02034_));
 AO21x1_ASAP7_75t_SL _24367_ (.A1(_01967_),
    .A2(_02034_),
    .B(_01660_),
    .Y(_02035_));
 AOI21x1_ASAP7_75t_SL _24368_ (.A1(_02035_),
    .A2(_01915_),
    .B(_01687_),
    .Y(_02036_));
 NOR2x1_ASAP7_75t_SL _24369_ (.A(_02032_),
    .B(_02036_),
    .Y(_02037_));
 AOI21x1_ASAP7_75t_SL _24370_ (.A1(_01694_),
    .A2(_01880_),
    .B(_01940_),
    .Y(_02038_));
 NAND2x1_ASAP7_75t_SL _24371_ (.A(_01939_),
    .B(_02038_),
    .Y(_02039_));
 OAI21x1_ASAP7_75t_R _24372_ (.A1(_01611_),
    .A2(_01638_),
    .B(_01835_),
    .Y(_02040_));
 NAND2x1_ASAP7_75t_SL _24373_ (.A(_01694_),
    .B(_02040_),
    .Y(_02041_));
 INVx1_ASAP7_75t_SL _24374_ (.A(_01785_),
    .Y(_02042_));
 AOI21x1_ASAP7_75t_SL _24375_ (.A1(_02042_),
    .A2(_01700_),
    .B(_01921_),
    .Y(_02043_));
 NAND2x1_ASAP7_75t_SL _24376_ (.A(_02041_),
    .B(_02043_),
    .Y(_02044_));
 NAND2x1_ASAP7_75t_SL _24377_ (.A(_02039_),
    .B(_02044_),
    .Y(_02045_));
 OAI21x1_ASAP7_75t_SL _24378_ (.A1(_02037_),
    .A2(_02045_),
    .B(_01801_),
    .Y(_02046_));
 AOI21x1_ASAP7_75t_SL _24379_ (.A1(_02031_),
    .A2(_02046_),
    .B(_01753_),
    .Y(_02047_));
 AO21x1_ASAP7_75t_SL _24380_ (.A1(_01879_),
    .A2(_01897_),
    .B(_01660_),
    .Y(_02048_));
 AOI21x1_ASAP7_75t_SL _24381_ (.A1(_01660_),
    .A2(_01961_),
    .B(_01720_),
    .Y(_02049_));
 NAND2x1_ASAP7_75t_SL _24382_ (.A(_02048_),
    .B(_02049_),
    .Y(_02050_));
 INVx1_ASAP7_75t_SL _24383_ (.A(_01731_),
    .Y(_02051_));
 AOI21x1_ASAP7_75t_SL _24384_ (.A1(_01690_),
    .A2(_01912_),
    .B(_01829_),
    .Y(_02052_));
 OAI21x1_ASAP7_75t_SL _24385_ (.A1(_01741_),
    .A2(_02051_),
    .B(_02052_),
    .Y(_02053_));
 AOI21x1_ASAP7_75t_SL _24386_ (.A1(_02050_),
    .A2(_02053_),
    .B(_01687_),
    .Y(_02054_));
 AND2x2_ASAP7_75t_SL _24387_ (.A(_01694_),
    .B(_01725_),
    .Y(_02055_));
 NOR2x1_ASAP7_75t_SL _24388_ (.A(_01921_),
    .B(_02055_),
    .Y(_02056_));
 AO21x1_ASAP7_75t_SL _24389_ (.A1(_01691_),
    .A2(_01709_),
    .B(_01694_),
    .Y(_02057_));
 OR3x1_ASAP7_75t_SL _24390_ (.A(_01660_),
    .B(_01735_),
    .C(_01633_),
    .Y(_02058_));
 NAND3x1_ASAP7_75t_SL _24391_ (.A(_02058_),
    .B(_02057_),
    .C(_02056_),
    .Y(_02059_));
 AO21x1_ASAP7_75t_SL _24392_ (.A1(_01892_),
    .A2(_01642_),
    .B(_01694_),
    .Y(_02060_));
 NOR3x1_ASAP7_75t_SL _24393_ (.A(_01928_),
    .B(_01686_),
    .C(_01829_),
    .Y(_02061_));
 AOI21x1_ASAP7_75t_SL _24394_ (.A1(_02060_),
    .A2(_02061_),
    .B(_01801_),
    .Y(_02062_));
 NAND2x1_ASAP7_75t_SL _24395_ (.A(_02059_),
    .B(_02062_),
    .Y(_02063_));
 NOR2x1_ASAP7_75t_SL _24396_ (.A(_02054_),
    .B(_02063_),
    .Y(_02064_));
 AO21x1_ASAP7_75t_SL _24397_ (.A1(_01946_),
    .A2(_01818_),
    .B(_02055_),
    .Y(_02065_));
 INVx1_ASAP7_75t_SL _24398_ (.A(_01729_),
    .Y(_02066_));
 OAI21x1_ASAP7_75t_SL _24399_ (.A1(_01720_),
    .A2(_02066_),
    .B(_01823_),
    .Y(_02067_));
 AOI21x1_ASAP7_75t_SL _24400_ (.A1(_01720_),
    .A2(_02065_),
    .B(_02067_),
    .Y(_02068_));
 AOI21x1_ASAP7_75t_SL _24401_ (.A1(_01694_),
    .A2(_01836_),
    .B(_01940_),
    .Y(_02069_));
 AOI21x1_ASAP7_75t_SL _24402_ (.A1(_01968_),
    .A2(_02069_),
    .B(_01907_),
    .Y(_02070_));
 OAI21x1_ASAP7_75t_SL _24403_ (.A1(_01624_),
    .A2(_01632_),
    .B(_01724_),
    .Y(_02071_));
 AO21x2_ASAP7_75t_SL _24404_ (.A1(_02071_),
    .A2(_01691_),
    .B(_01694_),
    .Y(_02072_));
 AO21x1_ASAP7_75t_SL _24405_ (.A1(_01949_),
    .A2(_02034_),
    .B(_01660_),
    .Y(_02073_));
 NOR2x1_ASAP7_75t_SL _24406_ (.A(_01687_),
    .B(_01829_),
    .Y(_02074_));
 NAND3x1_ASAP7_75t_SL _24407_ (.A(_02072_),
    .B(_02073_),
    .C(_02074_),
    .Y(_02075_));
 NAND2x1_ASAP7_75t_SL _24408_ (.A(_02070_),
    .B(_02075_),
    .Y(_02076_));
 OAI21x1_ASAP7_75t_SL _24409_ (.A1(_02068_),
    .A2(_02076_),
    .B(_01753_),
    .Y(_02077_));
 NOR2x1_ASAP7_75t_SL _24410_ (.A(_02064_),
    .B(_02077_),
    .Y(_02078_));
 NOR2x1_ASAP7_75t_SL _24411_ (.A(_02047_),
    .B(_02078_),
    .Y(_00091_));
 AND3x1_ASAP7_75t_SL _24412_ (.A(_01642_),
    .B(_01694_),
    .C(_01825_),
    .Y(_02079_));
 AO21x1_ASAP7_75t_SL _24413_ (.A1(_01873_),
    .A2(_01770_),
    .B(_01694_),
    .Y(_02080_));
 NAND2x1_ASAP7_75t_SL _24414_ (.A(_01687_),
    .B(_02080_),
    .Y(_02081_));
 OAI21x1_ASAP7_75t_SL _24415_ (.A1(_02079_),
    .A2(_02081_),
    .B(_01720_),
    .Y(_02082_));
 AND3x1_ASAP7_75t_SL _24416_ (.A(_01662_),
    .B(_01686_),
    .C(_01805_),
    .Y(_02083_));
 NAND2x1_ASAP7_75t_SL _24417_ (.A(_01660_),
    .B(_01844_),
    .Y(_02084_));
 NOR2x1_ASAP7_75t_SL _24418_ (.A(_01216_),
    .B(_01638_),
    .Y(_02085_));
 OAI21x1_ASAP7_75t_SL _24419_ (.A1(_02085_),
    .A2(_01809_),
    .B(_01694_),
    .Y(_02086_));
 AOI21x1_ASAP7_75t_SL _24420_ (.A1(_02084_),
    .A2(_02086_),
    .B(_01921_),
    .Y(_02087_));
 NAND2x1_ASAP7_75t_SL _24421_ (.A(_01694_),
    .B(_01854_),
    .Y(_02088_));
 AO21x1_ASAP7_75t_SL _24422_ (.A1(_01659_),
    .A2(_01654_),
    .B(_01217_),
    .Y(_02089_));
 INVx1_ASAP7_75t_SL _24423_ (.A(_01940_),
    .Y(_02090_));
 AO31x2_ASAP7_75t_SL _24424_ (.A1(_02088_),
    .A2(_02089_),
    .A3(_02090_),
    .B(_01754_),
    .Y(_02091_));
 NOR2x1_ASAP7_75t_SL _24425_ (.A(_02087_),
    .B(_02091_),
    .Y(_02092_));
 OAI21x1_ASAP7_75t_SL _24426_ (.A1(_02082_),
    .A2(_02083_),
    .B(_02092_),
    .Y(_02093_));
 NAND2x1_ASAP7_75t_SL _24427_ (.A(_01686_),
    .B(_01760_),
    .Y(_02094_));
 NOR2x1_ASAP7_75t_SL _24428_ (.A(_01778_),
    .B(_02024_),
    .Y(_02095_));
 AO21x1_ASAP7_75t_SL _24429_ (.A1(_01703_),
    .A2(_01633_),
    .B(_01660_),
    .Y(_02096_));
 NOR2x1_ASAP7_75t_SL _24430_ (.A(_01761_),
    .B(_01638_),
    .Y(_02097_));
 OA21x2_ASAP7_75t_SL _24431_ (.A1(_02097_),
    .A2(_01694_),
    .B(_01687_),
    .Y(_02098_));
 AOI21x1_ASAP7_75t_SL _24432_ (.A1(_02096_),
    .A2(_02098_),
    .B(_01720_),
    .Y(_02099_));
 OAI21x1_ASAP7_75t_SL _24433_ (.A1(_02094_),
    .A2(_02095_),
    .B(_02099_),
    .Y(_02100_));
 NOR2x1_ASAP7_75t_SL _24434_ (.A(_01687_),
    .B(_01923_),
    .Y(_02101_));
 AO21x1_ASAP7_75t_SL _24435_ (.A1(_01874_),
    .A2(_01949_),
    .B(_01694_),
    .Y(_02102_));
 AOI21x1_ASAP7_75t_SL _24436_ (.A1(_02101_),
    .A2(_02102_),
    .B(_01829_),
    .Y(_02103_));
 AO21x1_ASAP7_75t_SL _24437_ (.A1(_01731_),
    .A2(_01850_),
    .B(_01694_),
    .Y(_02104_));
 NAND2x1_ASAP7_75t_SL _24438_ (.A(_02104_),
    .B(_01911_),
    .Y(_02105_));
 AOI21x1_ASAP7_75t_SL _24439_ (.A1(_02103_),
    .A2(_02105_),
    .B(_01753_),
    .Y(_02106_));
 AOI21x1_ASAP7_75t_SL _24440_ (.A1(_02100_),
    .A2(_02106_),
    .B(_01907_),
    .Y(_02107_));
 NAND2x1_ASAP7_75t_SL _24441_ (.A(_02093_),
    .B(_02107_),
    .Y(_02108_));
 AO21x1_ASAP7_75t_SL _24442_ (.A1(_01731_),
    .A2(_01642_),
    .B(_01660_),
    .Y(_02109_));
 AOI21x1_ASAP7_75t_SL _24443_ (.A1(_01920_),
    .A2(_02109_),
    .B(_01940_),
    .Y(_02110_));
 NOR2x1_ASAP7_75t_SL _24444_ (.A(_01211_),
    .B(_01633_),
    .Y(_02111_));
 AO21x1_ASAP7_75t_SL _24445_ (.A1(_01825_),
    .A2(_01694_),
    .B(_02111_),
    .Y(_02112_));
 AO21x1_ASAP7_75t_SL _24446_ (.A1(_02112_),
    .A2(_01922_),
    .B(_01753_),
    .Y(_02113_));
 NOR2x1_ASAP7_75t_SL _24447_ (.A(_02110_),
    .B(_02113_),
    .Y(_02114_));
 AO21x1_ASAP7_75t_SL _24448_ (.A1(_01946_),
    .A2(_01708_),
    .B(_01660_),
    .Y(_02115_));
 AO21x1_ASAP7_75t_SL _24449_ (.A1(_01690_),
    .A2(_01731_),
    .B(_01694_),
    .Y(_02116_));
 AOI21x1_ASAP7_75t_SL _24450_ (.A1(_02115_),
    .A2(_02116_),
    .B(_01686_),
    .Y(_02117_));
 AO21x1_ASAP7_75t_SL _24451_ (.A1(_01731_),
    .A2(_01874_),
    .B(_01694_),
    .Y(_02118_));
 AOI21x1_ASAP7_75t_SL _24452_ (.A1(_02118_),
    .A2(_02003_),
    .B(_01687_),
    .Y(_02119_));
 OAI21x1_ASAP7_75t_SL _24453_ (.A1(_02117_),
    .A2(_02119_),
    .B(_01720_),
    .Y(_02120_));
 AOI21x1_ASAP7_75t_SL _24454_ (.A1(_02114_),
    .A2(_02120_),
    .B(_01801_),
    .Y(_02121_));
 AND3x1_ASAP7_75t_SL _24455_ (.A(_01819_),
    .B(_01694_),
    .C(_01731_),
    .Y(_02122_));
 NAND2x1_ASAP7_75t_SL _24456_ (.A(_01687_),
    .B(_01950_),
    .Y(_02123_));
 NAND2x1_ASAP7_75t_SL _24457_ (.A(_01850_),
    .B(_01892_),
    .Y(_02124_));
 AOI21x1_ASAP7_75t_SL _24458_ (.A1(_01694_),
    .A2(_02124_),
    .B(_01687_),
    .Y(_02125_));
 AOI21x1_ASAP7_75t_SL _24459_ (.A1(_01845_),
    .A2(_02125_),
    .B(_01829_),
    .Y(_02126_));
 OAI21x1_ASAP7_75t_SL _24460_ (.A1(_02122_),
    .A2(_02123_),
    .B(_02126_),
    .Y(_02127_));
 NAND2x1_ASAP7_75t_SL _24461_ (.A(_01660_),
    .B(_01772_),
    .Y(_02128_));
 OA21x2_ASAP7_75t_SL _24462_ (.A1(_02128_),
    .A2(_01725_),
    .B(_01686_),
    .Y(_02129_));
 NAND2x1_ASAP7_75t_SL _24463_ (.A(_01826_),
    .B(_02129_),
    .Y(_02130_));
 AO21x1_ASAP7_75t_SL _24464_ (.A1(_01837_),
    .A2(_01660_),
    .B(_01686_),
    .Y(_02131_));
 AO21x1_ASAP7_75t_SL _24465_ (.A1(_01854_),
    .A2(_01694_),
    .B(_01836_),
    .Y(_02132_));
 OA21x2_ASAP7_75t_SL _24466_ (.A1(_02131_),
    .A2(_02132_),
    .B(_01829_),
    .Y(_02133_));
 AOI21x1_ASAP7_75t_SL _24467_ (.A1(_02130_),
    .A2(_02133_),
    .B(_01754_),
    .Y(_02134_));
 NAND2x1_ASAP7_75t_SL _24468_ (.A(_02127_),
    .B(_02134_),
    .Y(_02135_));
 NAND2x1_ASAP7_75t_SL _24469_ (.A(_02121_),
    .B(_02135_),
    .Y(_02136_));
 NAND2x1_ASAP7_75t_SL _24470_ (.A(_02108_),
    .B(_02136_),
    .Y(_00092_));
 NOR2x1_ASAP7_75t_SL _24471_ (.A(_01694_),
    .B(_01642_),
    .Y(_02137_));
 OA21x2_ASAP7_75t_SL _24472_ (.A1(_01743_),
    .A2(_01660_),
    .B(_01687_),
    .Y(_02138_));
 NOR2x1_ASAP7_75t_SL _24473_ (.A(_01218_),
    .B(_01638_),
    .Y(_02139_));
 OAI21x1_ASAP7_75t_SL _24474_ (.A1(_02139_),
    .A2(_01758_),
    .B(_01660_),
    .Y(_02140_));
 AOI21x1_ASAP7_75t_SL _24475_ (.A1(_02138_),
    .A2(_02140_),
    .B(_01829_),
    .Y(_02141_));
 OAI21x1_ASAP7_75t_SL _24476_ (.A1(_01842_),
    .A2(_02137_),
    .B(_02141_),
    .Y(_02142_));
 OA21x2_ASAP7_75t_SL _24477_ (.A1(_01660_),
    .A2(_01635_),
    .B(_01686_),
    .Y(_02143_));
 AOI21x1_ASAP7_75t_SL _24478_ (.A1(_02143_),
    .A2(_01696_),
    .B(_01720_),
    .Y(_02144_));
 NAND2x1p5_ASAP7_75t_SL _24479_ (.A(_01742_),
    .B(_01780_),
    .Y(_02145_));
 OA21x2_ASAP7_75t_R _24480_ (.A1(_01834_),
    .A2(_01638_),
    .B(_01660_),
    .Y(_02146_));
 AOI21x1_ASAP7_75t_SL _24481_ (.A1(_01770_),
    .A2(_02146_),
    .B(_01686_),
    .Y(_02147_));
 NAND2x1_ASAP7_75t_SL _24482_ (.A(_02145_),
    .B(_02147_),
    .Y(_02148_));
 AOI21x1_ASAP7_75t_SL _24483_ (.A1(_02144_),
    .A2(_02148_),
    .B(_01753_),
    .Y(_02149_));
 AOI21x1_ASAP7_75t_SL _24484_ (.A1(_02142_),
    .A2(_02149_),
    .B(_01907_),
    .Y(_02150_));
 NAND2x1_ASAP7_75t_SL _24485_ (.A(_02071_),
    .B(_01660_),
    .Y(_02151_));
 AO21x1_ASAP7_75t_SL _24486_ (.A1(_02071_),
    .A2(_01743_),
    .B(_01660_),
    .Y(_02152_));
 OA21x2_ASAP7_75t_SL _24487_ (.A1(_01785_),
    .A2(_02151_),
    .B(_02152_),
    .Y(_02153_));
 AO21x1_ASAP7_75t_SL _24488_ (.A1(_01694_),
    .A2(_01215_),
    .B(_01687_),
    .Y(_02154_));
 OA21x2_ASAP7_75t_SL _24489_ (.A1(_01946_),
    .A2(_01635_),
    .B(_01660_),
    .Y(_02155_));
 OAI21x1_ASAP7_75t_SL _24490_ (.A1(_02154_),
    .A2(_02155_),
    .B(_01720_),
    .Y(_02156_));
 AO21x1_ASAP7_75t_SL _24491_ (.A1(_01687_),
    .A2(_02153_),
    .B(_02156_),
    .Y(_02157_));
 AO21x1_ASAP7_75t_SL _24492_ (.A1(_01985_),
    .A2(_01694_),
    .B(_01687_),
    .Y(_02158_));
 AO21x1_ASAP7_75t_SL _24493_ (.A1(_01769_),
    .A2(_01903_),
    .B(_02158_),
    .Y(_02159_));
 OA21x2_ASAP7_75t_SL _24494_ (.A1(_02131_),
    .A2(_01861_),
    .B(_01829_),
    .Y(_02160_));
 AOI21x1_ASAP7_75t_SL _24495_ (.A1(_02159_),
    .A2(_02160_),
    .B(_01754_),
    .Y(_02161_));
 NAND2x1_ASAP7_75t_SL _24496_ (.A(_02157_),
    .B(_02161_),
    .Y(_02162_));
 NAND2x1_ASAP7_75t_SL _24497_ (.A(_02150_),
    .B(_02162_),
    .Y(_02163_));
 NOR2x1_ASAP7_75t_SL _24498_ (.A(_01687_),
    .B(_01700_),
    .Y(_02164_));
 NAND2x1_ASAP7_75t_SL _24499_ (.A(_02041_),
    .B(_02164_),
    .Y(_02165_));
 OA21x2_ASAP7_75t_SL _24500_ (.A1(_01778_),
    .A2(_01694_),
    .B(_01687_),
    .Y(_02166_));
 AOI21x1_ASAP7_75t_SL _24501_ (.A1(_01924_),
    .A2(_02166_),
    .B(_01829_),
    .Y(_02167_));
 AOI21x1_ASAP7_75t_SL _24502_ (.A1(_02165_),
    .A2(_02167_),
    .B(_01753_),
    .Y(_02168_));
 AO21x1_ASAP7_75t_SL _24503_ (.A1(_01949_),
    .A2(_01865_),
    .B(_01660_),
    .Y(_02169_));
 AOI21x1_ASAP7_75t_SL _24504_ (.A1(_02169_),
    .A2(_01763_),
    .B(_01687_),
    .Y(_02170_));
 AO21x1_ASAP7_75t_SL _24505_ (.A1(_01762_),
    .A2(_01213_),
    .B(_01660_),
    .Y(_02171_));
 NAND2x1_ASAP7_75t_SL _24506_ (.A(_01819_),
    .B(_02146_),
    .Y(_02172_));
 AOI21x1_ASAP7_75t_SL _24507_ (.A1(_02171_),
    .A2(_02172_),
    .B(_01686_),
    .Y(_02173_));
 OAI21x1_ASAP7_75t_SL _24508_ (.A1(_02170_),
    .A2(_02173_),
    .B(_01829_),
    .Y(_02174_));
 AOI21x1_ASAP7_75t_SL _24509_ (.A1(_02168_),
    .A2(_02174_),
    .B(_01801_),
    .Y(_02175_));
 INVx1_ASAP7_75t_R _24510_ (.A(_01743_),
    .Y(_02176_));
 OAI21x1_ASAP7_75t_SL _24511_ (.A1(_02176_),
    .A2(_01758_),
    .B(_01694_),
    .Y(_02177_));
 AO21x1_ASAP7_75t_SL _24512_ (.A1(_01873_),
    .A2(_01767_),
    .B(_01694_),
    .Y(_02178_));
 AOI21x1_ASAP7_75t_SL _24513_ (.A1(_02177_),
    .A2(_02178_),
    .B(_01686_),
    .Y(_02179_));
 OA21x2_ASAP7_75t_SL _24514_ (.A1(_01660_),
    .A2(_01595_),
    .B(_01686_),
    .Y(_02180_));
 AO21x1_ASAP7_75t_SL _24515_ (.A1(_02080_),
    .A2(_02180_),
    .B(_01720_),
    .Y(_02181_));
 NOR2x1_ASAP7_75t_SL _24516_ (.A(_02179_),
    .B(_02181_),
    .Y(_02182_));
 INVx1_ASAP7_75t_R _24517_ (.A(_01847_),
    .Y(_02183_));
 OAI21x1_ASAP7_75t_SL _24518_ (.A1(_02183_),
    .A2(_01931_),
    .B(_01660_),
    .Y(_02184_));
 NAND3x1_ASAP7_75t_SL _24519_ (.A(_02184_),
    .B(_01687_),
    .C(_02088_),
    .Y(_02185_));
 NAND2x1p5_ASAP7_75t_SL _24520_ (.A(_01708_),
    .B(_01742_),
    .Y(_02186_));
 AO21x1_ASAP7_75t_SL _24521_ (.A1(_01970_),
    .A2(_02186_),
    .B(_01687_),
    .Y(_02187_));
 AOI21x1_ASAP7_75t_SL _24522_ (.A1(_02185_),
    .A2(_02187_),
    .B(_01829_),
    .Y(_02188_));
 OAI21x1_ASAP7_75t_SL _24523_ (.A1(_02188_),
    .A2(_02182_),
    .B(_01753_),
    .Y(_02189_));
 NAND2x1_ASAP7_75t_SL _24524_ (.A(_02175_),
    .B(_02189_),
    .Y(_02190_));
 NAND2x1_ASAP7_75t_SL _24525_ (.A(_02163_),
    .B(_02190_),
    .Y(_00093_));
 NOR2x1_ASAP7_75t_R _24526_ (.A(_01984_),
    .B(_01638_),
    .Y(_02191_));
 OA21x2_ASAP7_75t_R _24527_ (.A1(_02191_),
    .A2(_01836_),
    .B(_01694_),
    .Y(_02192_));
 NOR2x1_ASAP7_75t_SL _24528_ (.A(_01633_),
    .B(_01611_),
    .Y(_02193_));
 OA21x2_ASAP7_75t_SL _24529_ (.A1(_01725_),
    .A2(_02193_),
    .B(_01660_),
    .Y(_02194_));
 OAI21x1_ASAP7_75t_SL _24530_ (.A1(_02192_),
    .A2(_02194_),
    .B(_01687_),
    .Y(_02195_));
 AND3x1_ASAP7_75t_L _24531_ (.A(_01825_),
    .B(_01772_),
    .C(_01660_),
    .Y(_02196_));
 AOI21x1_ASAP7_75t_R _24532_ (.A1(_01762_),
    .A2(_01957_),
    .B(_01660_),
    .Y(_02197_));
 OAI21x1_ASAP7_75t_R _24533_ (.A1(_02196_),
    .A2(_02197_),
    .B(_01686_),
    .Y(_02198_));
 AOI21x1_ASAP7_75t_R _24534_ (.A1(_02195_),
    .A2(_02198_),
    .B(_01829_),
    .Y(_02199_));
 AO21x1_ASAP7_75t_R _24535_ (.A1(_01847_),
    .A2(_01835_),
    .B(_01660_),
    .Y(_02200_));
 AND3x1_ASAP7_75t_R _24536_ (.A(_02200_),
    .B(_01687_),
    .C(_01737_),
    .Y(_02201_));
 NAND2x1_ASAP7_75t_R _24537_ (.A(_01226_),
    .B(_01220_),
    .Y(_02202_));
 AO21x1_ASAP7_75t_R _24538_ (.A1(_01660_),
    .A2(_02202_),
    .B(_01687_),
    .Y(_02203_));
 AO21x1_ASAP7_75t_R _24539_ (.A1(_01873_),
    .A2(_01770_),
    .B(_01660_),
    .Y(_02204_));
 INVx1_ASAP7_75t_R _24540_ (.A(_02204_),
    .Y(_02205_));
 OAI21x1_ASAP7_75t_R _24541_ (.A1(_02203_),
    .A2(_02205_),
    .B(_01829_),
    .Y(_02206_));
 NOR2x1_ASAP7_75t_SL _24542_ (.A(_02201_),
    .B(_02206_),
    .Y(_02207_));
 NOR3x1_ASAP7_75t_L _24543_ (.A(_02199_),
    .B(_01753_),
    .C(_02207_),
    .Y(_02208_));
 INVx1_ASAP7_75t_R _24544_ (.A(_02034_),
    .Y(_02209_));
 OAI21x1_ASAP7_75t_R _24545_ (.A1(_01725_),
    .A2(_02209_),
    .B(_01660_),
    .Y(_02210_));
 OAI21x1_ASAP7_75t_R _24546_ (.A1(_01781_),
    .A2(_01844_),
    .B(_01694_),
    .Y(_02211_));
 NAND2x1_ASAP7_75t_R _24547_ (.A(_02210_),
    .B(_02211_),
    .Y(_02212_));
 OAI21x1_ASAP7_75t_SL _24548_ (.A1(_01633_),
    .A2(_01635_),
    .B(_01595_),
    .Y(_02213_));
 AOI21x1_ASAP7_75t_R _24549_ (.A1(_01694_),
    .A2(_02213_),
    .B(_01744_),
    .Y(_02214_));
 AOI21x1_ASAP7_75t_SL _24550_ (.A1(_01687_),
    .A2(_02214_),
    .B(_01829_),
    .Y(_02215_));
 OAI21x1_ASAP7_75t_SL _24551_ (.A1(_01687_),
    .A2(_02212_),
    .B(_02215_),
    .Y(_02216_));
 INVx1_ASAP7_75t_SL _24552_ (.A(_02071_),
    .Y(_02217_));
 AOI21x1_ASAP7_75t_R _24553_ (.A1(_01635_),
    .A2(_01595_),
    .B(_01638_),
    .Y(_02218_));
 OAI21x1_ASAP7_75t_SL _24554_ (.A1(_02218_),
    .A2(_02217_),
    .B(_01660_),
    .Y(_02219_));
 NAND3x1_ASAP7_75t_SL _24555_ (.A(_01992_),
    .B(_01687_),
    .C(_02219_),
    .Y(_02220_));
 AOI21x1_ASAP7_75t_R _24556_ (.A1(_01208_),
    .A2(_01638_),
    .B(_01660_),
    .Y(_02221_));
 AOI21x1_ASAP7_75t_SL _24557_ (.A1(_01698_),
    .A2(_01847_),
    .B(_01694_),
    .Y(_02222_));
 AOI21x1_ASAP7_75t_R _24558_ (.A1(_02221_),
    .A2(_01780_),
    .B(_02222_),
    .Y(_02223_));
 AOI21x1_ASAP7_75t_R _24559_ (.A1(_01686_),
    .A2(_02223_),
    .B(_01720_),
    .Y(_02224_));
 NAND2x1_ASAP7_75t_L _24560_ (.A(_02220_),
    .B(_02224_),
    .Y(_02225_));
 NAND2x1_ASAP7_75t_SL _24561_ (.A(_02216_),
    .B(_02225_),
    .Y(_02226_));
 OAI21x1_ASAP7_75t_R _24562_ (.A1(_01754_),
    .A2(_02226_),
    .B(_01907_),
    .Y(_02227_));
 AOI21x1_ASAP7_75t_R _24563_ (.A1(_01694_),
    .A2(_01892_),
    .B(_01686_),
    .Y(_02228_));
 AOI21x1_ASAP7_75t_R _24564_ (.A1(_02228_),
    .A2(_01791_),
    .B(_01829_),
    .Y(_02229_));
 NOR2x1_ASAP7_75t_SL _24565_ (.A(_01694_),
    .B(_02071_),
    .Y(_02230_));
 AOI21x1_ASAP7_75t_R _24566_ (.A1(_01694_),
    .A2(_02040_),
    .B(_02230_),
    .Y(_02231_));
 NAND2x1_ASAP7_75t_SL _24567_ (.A(_02231_),
    .B(_01686_),
    .Y(_02232_));
 NAND2x1_ASAP7_75t_L _24568_ (.A(_02229_),
    .B(_02232_),
    .Y(_02233_));
 INVx1_ASAP7_75t_R _24569_ (.A(_02002_),
    .Y(_02234_));
 AOI21x1_ASAP7_75t_R _24570_ (.A1(_02128_),
    .A2(_02234_),
    .B(_01757_),
    .Y(_02235_));
 AOI21x1_ASAP7_75t_R _24571_ (.A1(_01766_),
    .A2(_02017_),
    .B(_01720_),
    .Y(_02236_));
 OAI21x1_ASAP7_75t_R _24572_ (.A1(_01686_),
    .A2(_02235_),
    .B(_02236_),
    .Y(_02237_));
 AOI21x1_ASAP7_75t_R _24573_ (.A1(_02233_),
    .A2(_02237_),
    .B(_01753_),
    .Y(_02238_));
 OAI21x1_ASAP7_75t_R _24574_ (.A1(_01867_),
    .A2(_02139_),
    .B(_01694_),
    .Y(_02239_));
 AOI21x1_ASAP7_75t_R _24575_ (.A1(_01660_),
    .A2(_01757_),
    .B(_01686_),
    .Y(_02240_));
 NAND2x1_ASAP7_75t_SL _24576_ (.A(_02239_),
    .B(_02240_),
    .Y(_02241_));
 NAND2x1_ASAP7_75t_R _24577_ (.A(_01660_),
    .B(_01825_),
    .Y(_02242_));
 AOI21x1_ASAP7_75t_R _24578_ (.A1(_01221_),
    .A2(_01694_),
    .B(_01687_),
    .Y(_02243_));
 OAI21x1_ASAP7_75t_SL _24579_ (.A1(_01931_),
    .A2(_02242_),
    .B(_02243_),
    .Y(_02244_));
 NAND3x1_ASAP7_75t_L _24580_ (.A(_02241_),
    .B(_02244_),
    .C(_01829_),
    .Y(_02245_));
 OAI21x1_ASAP7_75t_R _24581_ (.A1(_01611_),
    .A2(_01946_),
    .B(_01988_),
    .Y(_02246_));
 AOI21x1_ASAP7_75t_R _24582_ (.A1(_01694_),
    .A2(_02246_),
    .B(_01687_),
    .Y(_02247_));
 INVx1_ASAP7_75t_R _24583_ (.A(_01818_),
    .Y(_02248_));
 AOI21x1_ASAP7_75t_R _24584_ (.A1(_02248_),
    .A2(_02086_),
    .B(_01686_),
    .Y(_02249_));
 OAI21x1_ASAP7_75t_R _24585_ (.A1(_02247_),
    .A2(_02249_),
    .B(_01720_),
    .Y(_02250_));
 AOI21x1_ASAP7_75t_R _24586_ (.A1(_02245_),
    .A2(_02250_),
    .B(_01754_),
    .Y(_02251_));
 OAI21x1_ASAP7_75t_SL _24587_ (.A1(_02251_),
    .A2(_02238_),
    .B(_01801_),
    .Y(_02252_));
 OAI21x1_ASAP7_75t_SL _24588_ (.A1(_02208_),
    .A2(_02227_),
    .B(_02252_),
    .Y(_00094_));
 AOI221x1_ASAP7_75t_R _24589_ (.A1(_02071_),
    .A2(_01928_),
    .B1(_01770_),
    .B2(_01782_),
    .C(_01686_),
    .Y(_02253_));
 AO21x1_ASAP7_75t_R _24590_ (.A1(_01876_),
    .A2(_01835_),
    .B(_01694_),
    .Y(_02254_));
 OA21x2_ASAP7_75t_R _24591_ (.A1(_01660_),
    .A2(_01226_),
    .B(_01686_),
    .Y(_02255_));
 AO21x1_ASAP7_75t_SL _24592_ (.A1(_02255_),
    .A2(_02254_),
    .B(_01829_),
    .Y(_02256_));
 NAND2x1_ASAP7_75t_R _24593_ (.A(_01217_),
    .B(_01694_),
    .Y(_02257_));
 AOI21x1_ASAP7_75t_R _24594_ (.A1(_02257_),
    .A2(_01849_),
    .B(_01720_),
    .Y(_02258_));
 NAND2x1_ASAP7_75t_R _24595_ (.A(_01660_),
    .B(_02213_),
    .Y(_02259_));
 NAND2x1_ASAP7_75t_SL _24596_ (.A(_02259_),
    .B(_01911_),
    .Y(_02260_));
 AOI21x1_ASAP7_75t_R _24597_ (.A1(_02258_),
    .A2(_02260_),
    .B(_01754_),
    .Y(_02261_));
 OAI21x1_ASAP7_75t_SL _24598_ (.A1(_02256_),
    .A2(_02253_),
    .B(_02261_),
    .Y(_02262_));
 AO21x1_ASAP7_75t_R _24599_ (.A1(_01767_),
    .A2(_01595_),
    .B(_01694_),
    .Y(_02263_));
 NAND2x1_ASAP7_75t_SL _24600_ (.A(_01967_),
    .B(_02034_),
    .Y(_02264_));
 AOI21x1_ASAP7_75t_R _24601_ (.A1(_01694_),
    .A2(_02264_),
    .B(_01720_),
    .Y(_02265_));
 NAND2x1_ASAP7_75t_R _24602_ (.A(_02263_),
    .B(_02265_),
    .Y(_02266_));
 OA21x2_ASAP7_75t_R _24603_ (.A1(_01213_),
    .A2(_01694_),
    .B(_01720_),
    .Y(_02267_));
 AOI21x1_ASAP7_75t_R _24604_ (.A1(_02267_),
    .A2(_02204_),
    .B(_01686_),
    .Y(_02268_));
 AOI21x1_ASAP7_75t_R _24605_ (.A1(_02266_),
    .A2(_02268_),
    .B(_01753_),
    .Y(_02269_));
 NOR2x1_ASAP7_75t_SL _24606_ (.A(_01736_),
    .B(_01868_),
    .Y(_02270_));
 AO21x1_ASAP7_75t_SL _24607_ (.A1(_01743_),
    .A2(_01698_),
    .B(_01660_),
    .Y(_02271_));
 OAI21x1_ASAP7_75t_R _24608_ (.A1(_01694_),
    .A2(_02270_),
    .B(_02271_),
    .Y(_02272_));
 NAND2x1_ASAP7_75t_R _24609_ (.A(_01208_),
    .B(_01923_),
    .Y(_02273_));
 NOR3x1_ASAP7_75t_R _24610_ (.A(_01848_),
    .B(_01829_),
    .C(_01736_),
    .Y(_02274_));
 AOI21x1_ASAP7_75t_R _24611_ (.A1(_02273_),
    .A2(_02274_),
    .B(_01687_),
    .Y(_02275_));
 OAI21x1_ASAP7_75t_R _24612_ (.A1(_01720_),
    .A2(_02272_),
    .B(_02275_),
    .Y(_02276_));
 AOI21x1_ASAP7_75t_R _24613_ (.A1(_02269_),
    .A2(_02276_),
    .B(_01801_),
    .Y(_02277_));
 NAND2x1_ASAP7_75t_SL _24614_ (.A(_02262_),
    .B(_02277_),
    .Y(_02278_));
 AO21x1_ASAP7_75t_R _24615_ (.A1(_02002_),
    .A2(_01946_),
    .B(_01687_),
    .Y(_02279_));
 AND3x1_ASAP7_75t_SL _24616_ (.A(_01704_),
    .B(_01660_),
    .C(_01770_),
    .Y(_02280_));
 NOR2x1_ASAP7_75t_R _24617_ (.A(_02279_),
    .B(_02280_),
    .Y(_02281_));
 NAND2x1_ASAP7_75t_R _24618_ (.A(_01635_),
    .B(_01660_),
    .Y(_02282_));
 AO21x1_ASAP7_75t_R _24619_ (.A1(_02109_),
    .A2(_02282_),
    .B(_01686_),
    .Y(_02283_));
 NAND2x1_ASAP7_75t_R _24620_ (.A(_01829_),
    .B(_02283_),
    .Y(_02284_));
 NOR2x1_ASAP7_75t_R _24621_ (.A(_01687_),
    .B(_01729_),
    .Y(_02285_));
 AOI21x1_ASAP7_75t_SL _24622_ (.A1(_02285_),
    .A2(_01925_),
    .B(_01829_),
    .Y(_02286_));
 AO21x1_ASAP7_75t_SL _24623_ (.A1(_01633_),
    .A2(_01703_),
    .B(_02151_),
    .Y(_02287_));
 AOI21x1_ASAP7_75t_R _24624_ (.A1(_01694_),
    .A2(_01819_),
    .B(_01686_),
    .Y(_02288_));
 NAND2x1_ASAP7_75t_L _24625_ (.A(_02287_),
    .B(_02288_),
    .Y(_02289_));
 AOI21x1_ASAP7_75t_SL _24626_ (.A1(_02289_),
    .A2(_02286_),
    .B(_01754_),
    .Y(_02290_));
 OAI21x1_ASAP7_75t_SL _24627_ (.A1(_02281_),
    .A2(_02284_),
    .B(_02290_),
    .Y(_02291_));
 AO21x1_ASAP7_75t_SL _24628_ (.A1(_01897_),
    .A2(_01808_),
    .B(_01660_),
    .Y(_02292_));
 AOI21x1_ASAP7_75t_SL _24629_ (.A1(_02292_),
    .A2(_02072_),
    .B(_01686_),
    .Y(_02293_));
 AO21x1_ASAP7_75t_R _24630_ (.A1(_01967_),
    .A2(_01897_),
    .B(_01694_),
    .Y(_02294_));
 AOI21x1_ASAP7_75t_R _24631_ (.A1(_02294_),
    .A2(_02006_),
    .B(_01687_),
    .Y(_02295_));
 OAI21x1_ASAP7_75t_SL _24632_ (.A1(_02293_),
    .A2(_02295_),
    .B(_01720_),
    .Y(_02296_));
 AOI21x1_ASAP7_75t_R _24633_ (.A1(_01660_),
    .A2(_01772_),
    .B(_01687_),
    .Y(_02297_));
 AOI21x1_ASAP7_75t_R _24634_ (.A1(_02297_),
    .A2(_02086_),
    .B(_01720_),
    .Y(_02298_));
 AO21x1_ASAP7_75t_R _24635_ (.A1(_01208_),
    .A2(_01638_),
    .B(_01611_),
    .Y(_02299_));
 AOI21x1_ASAP7_75t_R _24636_ (.A1(_01660_),
    .A2(_02299_),
    .B(_01686_),
    .Y(_02300_));
 OAI21x1_ASAP7_75t_R _24637_ (.A1(_01660_),
    .A2(_02270_),
    .B(_02300_),
    .Y(_02301_));
 AOI21x1_ASAP7_75t_R _24638_ (.A1(_02298_),
    .A2(_02301_),
    .B(_01753_),
    .Y(_02302_));
 AOI21x1_ASAP7_75t_SL _24639_ (.A1(_02302_),
    .A2(_02296_),
    .B(_01907_),
    .Y(_02303_));
 NAND2x1_ASAP7_75t_SL _24640_ (.A(_02303_),
    .B(_02291_),
    .Y(_02304_));
 NAND2x1_ASAP7_75t_SL _24641_ (.A(_02278_),
    .B(_02304_),
    .Y(_00095_));
 NOR2x1_ASAP7_75t_R _24642_ (.A(_00574_),
    .B(_00468_),
    .Y(_02305_));
 XOR2x2_ASAP7_75t_SL _24643_ (.A(_13463_),
    .B(_10706_),
    .Y(_02306_));
 XOR2x2_ASAP7_75t_SL _24644_ (.A(_00678_),
    .B(_00671_),
    .Y(_02307_));
 INVx1_ASAP7_75t_R _24645_ (.A(_00672_),
    .Y(_02308_));
 XOR2x2_ASAP7_75t_SL _24646_ (.A(_02307_),
    .B(_02308_),
    .Y(_02309_));
 INVx1_ASAP7_75t_SL _24647_ (.A(_02309_),
    .Y(_02310_));
 NAND2x1_ASAP7_75t_R _24648_ (.A(_02306_),
    .B(_02310_),
    .Y(_02311_));
 INVx1_ASAP7_75t_R _24649_ (.A(_02306_),
    .Y(_02312_));
 NAND2x1_ASAP7_75t_L _24650_ (.A(_02309_),
    .B(_02312_),
    .Y(_02313_));
 AOI21x1_ASAP7_75t_SL _24651_ (.A1(_02313_),
    .A2(_02311_),
    .B(_10675_),
    .Y(_02314_));
 OAI21x1_ASAP7_75t_SL _24652_ (.A1(_02305_),
    .A2(_02314_),
    .B(_00869_),
    .Y(_02315_));
 AND2x2_ASAP7_75t_R _24653_ (.A(_10675_),
    .B(_00468_),
    .Y(_02316_));
 XOR2x2_ASAP7_75t_SL _24654_ (.A(_02306_),
    .B(_02309_),
    .Y(_02317_));
 NOR2x1p5_ASAP7_75t_L _24655_ (.A(_10675_),
    .B(_02317_),
    .Y(_02318_));
 INVx1_ASAP7_75t_R _24656_ (.A(_00869_),
    .Y(_02319_));
 OAI21x1_ASAP7_75t_R _24657_ (.A1(_02316_),
    .A2(_02318_),
    .B(_02319_),
    .Y(_02320_));
 NAND2x2_ASAP7_75t_SL _24658_ (.A(_02320_),
    .B(_02315_),
    .Y(_01233_));
 NOR2x1_ASAP7_75t_L _24659_ (.A(_00574_),
    .B(_00469_),
    .Y(_02321_));
 XOR2x2_ASAP7_75t_SL _24660_ (.A(_00607_),
    .B(_00646_),
    .Y(_02322_));
 XOR2x2_ASAP7_75t_SL _24661_ (.A(_02322_),
    .B(_00575_),
    .Y(_02323_));
 NAND2x1_ASAP7_75t_R _24662_ (.A(_02307_),
    .B(_02323_),
    .Y(_02324_));
 NOR2x1_ASAP7_75t_L _24663_ (.A(_02307_),
    .B(_02323_),
    .Y(_02325_));
 INVx1_ASAP7_75t_R _24664_ (.A(_02325_),
    .Y(_02326_));
 AOI21x1_ASAP7_75t_SL _24665_ (.A1(_02324_),
    .A2(_02326_),
    .B(_10675_),
    .Y(_02327_));
 OAI21x1_ASAP7_75t_R _24666_ (.A1(_02321_),
    .A2(_02327_),
    .B(_00868_),
    .Y(_02328_));
 INVx1_ASAP7_75t_R _24667_ (.A(_02307_),
    .Y(_02329_));
 XNOR2x2_ASAP7_75t_R _24668_ (.A(_00575_),
    .B(_02322_),
    .Y(_02330_));
 NOR2x1_ASAP7_75t_SL _24669_ (.A(_02329_),
    .B(_02330_),
    .Y(_02331_));
 OAI21x1_ASAP7_75t_R _24670_ (.A1(_02325_),
    .A2(_02331_),
    .B(_00574_),
    .Y(_02332_));
 INVx1_ASAP7_75t_R _24671_ (.A(_00868_),
    .Y(_02333_));
 INVx1_ASAP7_75t_R _24672_ (.A(_02321_),
    .Y(_02334_));
 NAND3x1_ASAP7_75t_SL _24673_ (.A(_02332_),
    .B(_02333_),
    .C(_02334_),
    .Y(_02335_));
 NAND2x2_ASAP7_75t_SL _24674_ (.A(_02328_),
    .B(_02335_),
    .Y(_01236_));
 NAND2x1_ASAP7_75t_R _24675_ (.A(_00470_),
    .B(_10675_),
    .Y(_02336_));
 XOR2x2_ASAP7_75t_SL _24676_ (.A(_00577_),
    .B(_00609_),
    .Y(_02337_));
 INVx2_ASAP7_75t_SL _24677_ (.A(_02337_),
    .Y(_02338_));
 INVx1_ASAP7_75t_R _24678_ (.A(_00673_),
    .Y(_02339_));
 XOR2x1_ASAP7_75t_SL _24679_ (.A(_13464_),
    .Y(_02340_),
    .B(_02339_));
 NAND2x1_ASAP7_75t_SL _24680_ (.A(_02338_),
    .B(_02340_),
    .Y(_02341_));
 NOR2x1_ASAP7_75t_L _24681_ (.A(_02339_),
    .B(_13464_),
    .Y(_02342_));
 XNOR2x2_ASAP7_75t_L _24682_ (.A(_00640_),
    .B(_00672_),
    .Y(_02343_));
 NOR2x1_ASAP7_75t_R _24683_ (.A(_00673_),
    .B(_02343_),
    .Y(_02344_));
 OAI21x1_ASAP7_75t_SL _24684_ (.A1(_02342_),
    .A2(_02344_),
    .B(_02337_),
    .Y(_02345_));
 NAND3x1_ASAP7_75t_R _24685_ (.A(_02341_),
    .B(_00574_),
    .C(_02345_),
    .Y(_02346_));
 AOI21x1_ASAP7_75t_SL _24686_ (.A1(_02336_),
    .A2(_02346_),
    .B(_00839_),
    .Y(_02347_));
 NOR2x1_ASAP7_75t_R _24687_ (.A(_00574_),
    .B(_00470_),
    .Y(_02348_));
 INVx1_ASAP7_75t_R _24688_ (.A(_02348_),
    .Y(_02349_));
 AOI21x1_ASAP7_75t_SL _24689_ (.A1(_02345_),
    .A2(_02341_),
    .B(_10675_),
    .Y(_02350_));
 INVx1_ASAP7_75t_R _24690_ (.A(_02350_),
    .Y(_02351_));
 INVx1_ASAP7_75t_R _24691_ (.A(_00839_),
    .Y(_02352_));
 AOI21x1_ASAP7_75t_SL _24692_ (.A1(_02349_),
    .A2(_02351_),
    .B(_02352_),
    .Y(_02353_));
 NOR2x2_ASAP7_75t_SL _24693_ (.A(_02347_),
    .B(_02353_),
    .Y(_02354_));
 OAI21x1_ASAP7_75t_SL _24695_ (.A1(_02314_),
    .A2(_02305_),
    .B(_02319_),
    .Y(_02355_));
 OAI21x1_ASAP7_75t_SL _24696_ (.A1(_02318_),
    .A2(_02316_),
    .B(_00869_),
    .Y(_02356_));
 NAND2x1p5_ASAP7_75t_SL _24697_ (.A(_02356_),
    .B(_02355_),
    .Y(_02357_));
 AOI21x1_ASAP7_75t_SL _24699_ (.A1(_02336_),
    .A2(_02346_),
    .B(_02352_),
    .Y(_02358_));
 AOI21x1_ASAP7_75t_SL _24700_ (.A1(_02349_),
    .A2(_02351_),
    .B(_00839_),
    .Y(_02359_));
 NOR2x2_ASAP7_75t_SL _24701_ (.A(_02358_),
    .B(_02359_),
    .Y(_02360_));
 NAND2x1_ASAP7_75t_SL _24704_ (.A(_02360_),
    .B(_01236_),
    .Y(_02362_));
 OAI21x1_ASAP7_75t_SL _24705_ (.A1(_02358_),
    .A2(_02359_),
    .B(_01237_),
    .Y(_02363_));
 XNOR2x2_ASAP7_75t_L _24706_ (.A(_00674_),
    .B(_13519_),
    .Y(_02364_));
 XNOR2x2_ASAP7_75t_R _24707_ (.A(_00673_),
    .B(_00678_),
    .Y(_02365_));
 XOR2x2_ASAP7_75t_R _24708_ (.A(_00578_),
    .B(_00610_),
    .Y(_02366_));
 XOR2x2_ASAP7_75t_SL _24709_ (.A(_02365_),
    .B(_02366_),
    .Y(_02367_));
 AOI21x1_ASAP7_75t_R _24710_ (.A1(_02364_),
    .A2(_02367_),
    .B(_10675_),
    .Y(_02368_));
 OR2x2_ASAP7_75t_SL _24711_ (.A(_02367_),
    .B(_02364_),
    .Y(_02369_));
 AND2x2_ASAP7_75t_R _24712_ (.A(_10675_),
    .B(_00564_),
    .Y(_02370_));
 AOI21x1_ASAP7_75t_SL _24713_ (.A1(_02368_),
    .A2(_02369_),
    .B(_02370_),
    .Y(_02371_));
 XOR2x2_ASAP7_75t_SL _24714_ (.A(_02371_),
    .B(_00840_),
    .Y(_02372_));
 AO21x1_ASAP7_75t_SL _24717_ (.A1(_02362_),
    .A2(_02363_),
    .B(_02372_),
    .Y(_02375_));
 OAI21x1_ASAP7_75t_SL _24719_ (.A1(_02358_),
    .A2(_02359_),
    .B(_01231_),
    .Y(_02377_));
 NAND2x2_ASAP7_75t_SL _24720_ (.A(_02360_),
    .B(_02357_),
    .Y(_02378_));
 XNOR2x2_ASAP7_75t_SL _24721_ (.A(_00840_),
    .B(_02371_),
    .Y(_02379_));
 AOI21x1_ASAP7_75t_SL _24723_ (.A1(_02378_),
    .A2(_02377_),
    .B(_02379_),
    .Y(_02381_));
 INVx1_ASAP7_75t_SL _24724_ (.A(_02381_),
    .Y(_02382_));
 XOR2x2_ASAP7_75t_R _24725_ (.A(_00674_),
    .B(_00678_),
    .Y(_02383_));
 XOR2x2_ASAP7_75t_SL _24726_ (.A(_10828_),
    .B(_02383_),
    .Y(_02384_));
 XNOR2x2_ASAP7_75t_SL _24727_ (.A(_13551_),
    .B(_02384_),
    .Y(_02385_));
 NOR2x1_ASAP7_75t_R _24728_ (.A(_00574_),
    .B(_00563_),
    .Y(_02386_));
 AOI21x1_ASAP7_75t_R _24729_ (.A1(_00574_),
    .A2(_02385_),
    .B(_02386_),
    .Y(_02387_));
 XOR2x2_ASAP7_75t_SL _24730_ (.A(_02387_),
    .B(_00841_),
    .Y(_02388_));
 INVx2_ASAP7_75t_SL _24731_ (.A(_02388_),
    .Y(_02389_));
 AND3x1_ASAP7_75t_SL _24734_ (.A(_02375_),
    .B(_02382_),
    .C(_02389_),
    .Y(_02392_));
 INVx2_ASAP7_75t_SL _24738_ (.A(_01235_),
    .Y(_02396_));
 OA21x2_ASAP7_75t_R _24740_ (.A1(_02354_),
    .A2(_02396_),
    .B(_02379_),
    .Y(_02398_));
 NOR2x1_ASAP7_75t_SL _24741_ (.A(_02389_),
    .B(_02398_),
    .Y(_02399_));
 INVx1_ASAP7_75t_R _24742_ (.A(_01232_),
    .Y(_02400_));
 NAND2x1_ASAP7_75t_SL _24743_ (.A(_02400_),
    .B(_02360_),
    .Y(_02401_));
 NAND2x1_ASAP7_75t_SL _24744_ (.A(_01230_),
    .B(_02354_),
    .Y(_02402_));
 AO21x1_ASAP7_75t_SL _24746_ (.A1(_02401_),
    .A2(_02402_),
    .B(_02379_),
    .Y(_02404_));
 NOR2x1_ASAP7_75t_R _24747_ (.A(_00574_),
    .B(_00562_),
    .Y(_02405_));
 NAND2x1_ASAP7_75t_R _24748_ (.A(_00676_),
    .B(_10733_),
    .Y(_02406_));
 NAND2x1_ASAP7_75t_R _24749_ (.A(_13574_),
    .B(_10732_),
    .Y(_02407_));
 NAND3x1_ASAP7_75t_R _24750_ (.A(_02406_),
    .B(_02407_),
    .C(_10745_),
    .Y(_02408_));
 AOI21x1_ASAP7_75t_R _24751_ (.A1(_02407_),
    .A2(_02406_),
    .B(_10745_),
    .Y(_02409_));
 INVx1_ASAP7_75t_R _24752_ (.A(_02409_),
    .Y(_02410_));
 AOI21x1_ASAP7_75t_R _24753_ (.A1(_02408_),
    .A2(_02410_),
    .B(_10675_),
    .Y(_02411_));
 INVx1_ASAP7_75t_R _24754_ (.A(_00842_),
    .Y(_02412_));
 OAI21x1_ASAP7_75t_R _24755_ (.A1(_02405_),
    .A2(_02411_),
    .B(_02412_),
    .Y(_02413_));
 INVx1_ASAP7_75t_R _24756_ (.A(_10745_),
    .Y(_02414_));
 XOR2x2_ASAP7_75t_R _24757_ (.A(_10732_),
    .B(_00676_),
    .Y(_02415_));
 NOR2x1_ASAP7_75t_R _24758_ (.A(_02414_),
    .B(_02415_),
    .Y(_02416_));
 OAI21x1_ASAP7_75t_R _24759_ (.A1(_02409_),
    .A2(_02416_),
    .B(_00574_),
    .Y(_02417_));
 INVx1_ASAP7_75t_R _24760_ (.A(_02405_),
    .Y(_02418_));
 NAND3x1_ASAP7_75t_R _24761_ (.A(_02417_),
    .B(_00842_),
    .C(_02418_),
    .Y(_02419_));
 NAND2x1_ASAP7_75t_SL _24762_ (.A(_02413_),
    .B(_02419_),
    .Y(_02420_));
 AO21x1_ASAP7_75t_SL _24765_ (.A1(_02399_),
    .A2(_02404_),
    .B(_02420_),
    .Y(_02423_));
 OAI21x1_ASAP7_75t_R _24766_ (.A1(_02321_),
    .A2(_02327_),
    .B(_02333_),
    .Y(_02424_));
 NAND3x1_ASAP7_75t_L _24767_ (.A(_02332_),
    .B(_00868_),
    .C(_02334_),
    .Y(_02425_));
 NAND2x1_ASAP7_75t_SL _24768_ (.A(_02424_),
    .B(_02425_),
    .Y(_02426_));
 AOI21x1_ASAP7_75t_R _24771_ (.A1(_02354_),
    .A2(_02426_),
    .B(_02372_),
    .Y(_02428_));
 INVx2_ASAP7_75t_R _24772_ (.A(_01239_),
    .Y(_02429_));
 NAND2x1_ASAP7_75t_SL _24774_ (.A(_02429_),
    .B(_02360_),
    .Y(_02431_));
 OAI21x1_ASAP7_75t_SL _24776_ (.A1(_02358_),
    .A2(_02359_),
    .B(_02396_),
    .Y(_02433_));
 OAI21x1_ASAP7_75t_SL _24777_ (.A1(_02379_),
    .A2(_02433_),
    .B(_02389_),
    .Y(_02434_));
 AO21x1_ASAP7_75t_SL _24778_ (.A1(_02428_),
    .A2(_02431_),
    .B(_02434_),
    .Y(_02435_));
 INVx1_ASAP7_75t_R _24779_ (.A(_01238_),
    .Y(_02436_));
 OAI21x1_ASAP7_75t_R _24780_ (.A1(_02347_),
    .A2(_02353_),
    .B(_02436_),
    .Y(_02437_));
 AO21x2_ASAP7_75t_SL _24782_ (.A1(_02437_),
    .A2(_02433_),
    .B(_02379_),
    .Y(_02439_));
 OAI21x1_ASAP7_75t_SL _24783_ (.A1(_02347_),
    .A2(_02353_),
    .B(_01231_),
    .Y(_02440_));
 NAND2x1p5_ASAP7_75t_SL _24784_ (.A(_02440_),
    .B(_02379_),
    .Y(_02441_));
 AND2x2_ASAP7_75t_SL _24786_ (.A(_02441_),
    .B(_02388_),
    .Y(_02443_));
 INVx2_ASAP7_75t_SL _24787_ (.A(_02420_),
    .Y(_02444_));
 AOI21x1_ASAP7_75t_SL _24789_ (.A1(_02439_),
    .A2(_02443_),
    .B(_02444_),
    .Y(_02446_));
 XOR2x2_ASAP7_75t_R _24790_ (.A(_13608_),
    .B(_10879_),
    .Y(_02447_));
 XOR2x2_ASAP7_75t_SL _24791_ (.A(_02447_),
    .B(_10692_),
    .Y(_02448_));
 NOR2x1_ASAP7_75t_SL _24792_ (.A(_00574_),
    .B(_00560_),
    .Y(_02449_));
 AO21x1_ASAP7_75t_SL _24793_ (.A1(_02448_),
    .A2(_00574_),
    .B(_02449_),
    .Y(_02450_));
 XOR2x2_ASAP7_75t_SL _24794_ (.A(_02450_),
    .B(_00844_),
    .Y(_02451_));
 AOI21x1_ASAP7_75t_SL _24796_ (.A1(_02435_),
    .A2(_02446_),
    .B(_02451_),
    .Y(_02453_));
 OAI21x1_ASAP7_75t_SL _24797_ (.A1(_02392_),
    .A2(_02423_),
    .B(_02453_),
    .Y(_02454_));
 INVx2_ASAP7_75t_SL _24799_ (.A(_01234_),
    .Y(_02456_));
 NAND2x1_ASAP7_75t_SL _24800_ (.A(_02456_),
    .B(_02354_),
    .Y(_02457_));
 AND3x1_ASAP7_75t_SL _24801_ (.A(_02378_),
    .B(_02372_),
    .C(_02457_),
    .Y(_02458_));
 NAND2x2_ASAP7_75t_SL _24803_ (.A(_01240_),
    .B(_02360_),
    .Y(_02460_));
 AO21x1_ASAP7_75t_SL _24804_ (.A1(_02428_),
    .A2(_02460_),
    .B(_02389_),
    .Y(_02461_));
 NOR2x1_ASAP7_75t_SL _24805_ (.A(_01232_),
    .B(_02354_),
    .Y(_02462_));
 NOR2x1_ASAP7_75t_SL _24806_ (.A(_02360_),
    .B(_01233_),
    .Y(_02463_));
 OAI21x1_ASAP7_75t_SL _24807_ (.A1(_02462_),
    .A2(_02463_),
    .B(_02372_),
    .Y(_02464_));
 AOI21x1_ASAP7_75t_SL _24808_ (.A1(_02431_),
    .A2(_02428_),
    .B(_02388_),
    .Y(_02465_));
 AOI21x1_ASAP7_75t_SL _24809_ (.A1(_02464_),
    .A2(_02465_),
    .B(_02444_),
    .Y(_02466_));
 OAI21x1_ASAP7_75t_SL _24810_ (.A1(_02458_),
    .A2(_02461_),
    .B(_02466_),
    .Y(_02467_));
 NOR2x2_ASAP7_75t_SL _24811_ (.A(_02456_),
    .B(_02360_),
    .Y(_02468_));
 NOR2x1_ASAP7_75t_SL _24813_ (.A(_01235_),
    .B(_02354_),
    .Y(_02470_));
 OAI21x1_ASAP7_75t_SL _24815_ (.A1(_02468_),
    .A2(_02470_),
    .B(_02379_),
    .Y(_02472_));
 AOI21x1_ASAP7_75t_R _24817_ (.A1(_02354_),
    .A2(_02426_),
    .B(_02379_),
    .Y(_02474_));
 NOR2x1_ASAP7_75t_SL _24818_ (.A(_02388_),
    .B(_02474_),
    .Y(_02475_));
 AOI21x1_ASAP7_75t_SL _24819_ (.A1(_02472_),
    .A2(_02475_),
    .B(_02420_),
    .Y(_02476_));
 AOI21x1_ASAP7_75t_SL _24821_ (.A1(_01240_),
    .A2(_02354_),
    .B(_02372_),
    .Y(_02478_));
 NAND2x1_ASAP7_75t_SL _24822_ (.A(_02440_),
    .B(_02478_),
    .Y(_02479_));
 NAND2x1_ASAP7_75t_SL _24823_ (.A(_02360_),
    .B(_02426_),
    .Y(_02480_));
 OA21x2_ASAP7_75t_SL _24824_ (.A1(_02360_),
    .A2(_01234_),
    .B(_02372_),
    .Y(_02481_));
 AOI21x1_ASAP7_75t_SL _24826_ (.A1(_02480_),
    .A2(_02481_),
    .B(_02389_),
    .Y(_02483_));
 NAND2x1_ASAP7_75t_SL _24827_ (.A(_02479_),
    .B(_02483_),
    .Y(_02484_));
 INVx1_ASAP7_75t_SL _24828_ (.A(_02451_),
    .Y(_02485_));
 AOI21x1_ASAP7_75t_SL _24830_ (.A1(_02476_),
    .A2(_02484_),
    .B(_02485_),
    .Y(_02487_));
 XOR2x2_ASAP7_75t_SL _24831_ (.A(_00676_),
    .B(_00677_),
    .Y(_02488_));
 XOR2x2_ASAP7_75t_R _24832_ (.A(_02488_),
    .B(_00644_),
    .Y(_02489_));
 XOR2x2_ASAP7_75t_R _24833_ (.A(_02489_),
    .B(_10878_),
    .Y(_02490_));
 NOR2x1_ASAP7_75t_R _24834_ (.A(_00574_),
    .B(_00561_),
    .Y(_02491_));
 AO21x1_ASAP7_75t_SL _24835_ (.A1(_02490_),
    .A2(_00574_),
    .B(_02491_),
    .Y(_02492_));
 XOR2x2_ASAP7_75t_SL _24836_ (.A(_02492_),
    .B(_00843_),
    .Y(_02493_));
 AOI21x1_ASAP7_75t_SL _24838_ (.A1(_02467_),
    .A2(_02487_),
    .B(_02493_),
    .Y(_02495_));
 NAND2x1_ASAP7_75t_SL _24839_ (.A(_02454_),
    .B(_02495_),
    .Y(_02496_));
 OAI21x1_ASAP7_75t_SL _24840_ (.A1(_02347_),
    .A2(_02353_),
    .B(_01234_),
    .Y(_02497_));
 NOR2x1_ASAP7_75t_R _24841_ (.A(_02379_),
    .B(_02497_),
    .Y(_02498_));
 NOR2x1_ASAP7_75t_SL _24842_ (.A(_02498_),
    .B(_02434_),
    .Y(_02499_));
 INVx1_ASAP7_75t_SL _24843_ (.A(_02499_),
    .Y(_02500_));
 INVx1_ASAP7_75t_R _24844_ (.A(_01230_),
    .Y(_02501_));
 NAND2x1_ASAP7_75t_SL _24845_ (.A(_02501_),
    .B(_02360_),
    .Y(_02502_));
 AND3x1_ASAP7_75t_SL _24846_ (.A(_02354_),
    .B(_02400_),
    .C(_02372_),
    .Y(_02503_));
 AO21x1_ASAP7_75t_SL _24847_ (.A1(_02428_),
    .A2(_02502_),
    .B(_02503_),
    .Y(_02504_));
 NAND2x1_ASAP7_75t_R _24849_ (.A(_01245_),
    .B(_02379_),
    .Y(_02506_));
 INVx4_ASAP7_75t_R _24850_ (.A(_01231_),
    .Y(_02507_));
 AO21x1_ASAP7_75t_SL _24851_ (.A1(_02354_),
    .A2(_02507_),
    .B(_02379_),
    .Y(_02508_));
 NAND2x1_ASAP7_75t_SL _24852_ (.A(_02506_),
    .B(_02508_),
    .Y(_02509_));
 AOI21x1_ASAP7_75t_SL _24853_ (.A1(_02388_),
    .A2(_02509_),
    .B(_02444_),
    .Y(_02510_));
 OAI21x1_ASAP7_75t_SL _24854_ (.A1(_02500_),
    .A2(_02504_),
    .B(_02510_),
    .Y(_02511_));
 INVx1_ASAP7_75t_SL _24855_ (.A(_02497_),
    .Y(_02512_));
 NOR2x1_ASAP7_75t_SL _24856_ (.A(_01238_),
    .B(_02360_),
    .Y(_02513_));
 OAI21x1_ASAP7_75t_SL _24857_ (.A1(_02512_),
    .A2(_02513_),
    .B(_02379_),
    .Y(_02514_));
 NOR2x1_ASAP7_75t_R _24858_ (.A(_02379_),
    .B(_02401_),
    .Y(_02515_));
 INVx1_ASAP7_75t_SL _24859_ (.A(_02515_),
    .Y(_02516_));
 NAND3x1_ASAP7_75t_SL _24860_ (.A(_02514_),
    .B(_02516_),
    .C(_02389_),
    .Y(_02517_));
 OAI21x1_ASAP7_75t_R _24861_ (.A1(_02379_),
    .A2(_02497_),
    .B(_02388_),
    .Y(_02518_));
 INVx1_ASAP7_75t_SL _24862_ (.A(_02518_),
    .Y(_02519_));
 NOR2x1_ASAP7_75t_R _24863_ (.A(_02379_),
    .B(_02363_),
    .Y(_02520_));
 NOR2x1_ASAP7_75t_SL _24864_ (.A(_02372_),
    .B(_02401_),
    .Y(_02521_));
 NOR2x1_ASAP7_75t_SL _24865_ (.A(_02520_),
    .B(_02521_),
    .Y(_02522_));
 AOI21x1_ASAP7_75t_SL _24866_ (.A1(_02519_),
    .A2(_02522_),
    .B(_02420_),
    .Y(_02523_));
 AOI21x1_ASAP7_75t_SL _24867_ (.A1(_02517_),
    .A2(_02523_),
    .B(_02451_),
    .Y(_02524_));
 INVx1_ASAP7_75t_SL _24868_ (.A(_02493_),
    .Y(_02525_));
 AOI21x1_ASAP7_75t_SL _24870_ (.A1(_02511_),
    .A2(_02524_),
    .B(_02525_),
    .Y(_02527_));
 INVx1_ASAP7_75t_R _24871_ (.A(_01237_),
    .Y(_02528_));
 NOR2x1_ASAP7_75t_R _24872_ (.A(_02528_),
    .B(_02354_),
    .Y(_02529_));
 INVx1_ASAP7_75t_R _24873_ (.A(_02402_),
    .Y(_02530_));
 OAI21x1_ASAP7_75t_SL _24874_ (.A1(_02529_),
    .A2(_02530_),
    .B(_02379_),
    .Y(_02531_));
 NAND2x1_ASAP7_75t_SL _24875_ (.A(_02429_),
    .B(_02354_),
    .Y(_02532_));
 AND2x2_ASAP7_75t_L _24876_ (.A(_02440_),
    .B(_02372_),
    .Y(_02533_));
 NAND2x1_ASAP7_75t_SL _24877_ (.A(_02532_),
    .B(_02533_),
    .Y(_02534_));
 AOI21x1_ASAP7_75t_SL _24879_ (.A1(_02531_),
    .A2(_02534_),
    .B(_02388_),
    .Y(_02536_));
 NAND2x1_ASAP7_75t_SL _24880_ (.A(_02426_),
    .B(_02357_),
    .Y(_02537_));
 AOI21x1_ASAP7_75t_SL _24881_ (.A1(_02360_),
    .A2(_01236_),
    .B(_02379_),
    .Y(_02538_));
 NAND2x1_ASAP7_75t_SL _24882_ (.A(_02537_),
    .B(_02538_),
    .Y(_02539_));
 AO21x1_ASAP7_75t_SL _24884_ (.A1(_02537_),
    .A2(_02362_),
    .B(_02372_),
    .Y(_02541_));
 AOI21x1_ASAP7_75t_SL _24885_ (.A1(_02539_),
    .A2(_02541_),
    .B(_02389_),
    .Y(_02542_));
 OAI21x1_ASAP7_75t_SL _24887_ (.A1(_02536_),
    .A2(_02542_),
    .B(_02444_),
    .Y(_02544_));
 NAND2x2_ASAP7_75t_L _24888_ (.A(_02507_),
    .B(_02360_),
    .Y(_02545_));
 NAND2x1_ASAP7_75t_R _24889_ (.A(_02354_),
    .B(_01233_),
    .Y(_02546_));
 NAND2x1_ASAP7_75t_SL _24890_ (.A(_02545_),
    .B(_02546_),
    .Y(_02547_));
 AOI21x1_ASAP7_75t_SL _24891_ (.A1(_02379_),
    .A2(_02377_),
    .B(_02389_),
    .Y(_02548_));
 OAI21x1_ASAP7_75t_SL _24892_ (.A1(_02379_),
    .A2(_02547_),
    .B(_02548_),
    .Y(_02549_));
 OAI21x1_ASAP7_75t_R _24893_ (.A1(_02347_),
    .A2(_02353_),
    .B(_01230_),
    .Y(_02550_));
 AOI21x1_ASAP7_75t_SL _24894_ (.A1(_02363_),
    .A2(_02550_),
    .B(_02379_),
    .Y(_02551_));
 AOI21x1_ASAP7_75t_SL _24896_ (.A1(_02402_),
    .A2(_02545_),
    .B(_02372_),
    .Y(_02553_));
 OAI21x1_ASAP7_75t_SL _24897_ (.A1(_02551_),
    .A2(_02553_),
    .B(_02389_),
    .Y(_02554_));
 NAND2x1_ASAP7_75t_SL _24898_ (.A(_02549_),
    .B(_02554_),
    .Y(_02555_));
 AOI21x1_ASAP7_75t_SL _24899_ (.A1(_02420_),
    .A2(_02555_),
    .B(_02485_),
    .Y(_02556_));
 NAND2x1_ASAP7_75t_SL _24900_ (.A(_02544_),
    .B(_02556_),
    .Y(_02557_));
 NAND2x1_ASAP7_75t_SL _24901_ (.A(_02527_),
    .B(_02557_),
    .Y(_02558_));
 NAND2x1_ASAP7_75t_SL _24902_ (.A(_02496_),
    .B(_02558_),
    .Y(_00096_));
 OAI21x1_ASAP7_75t_R _24903_ (.A1(_02360_),
    .A2(_02426_),
    .B(_02372_),
    .Y(_02559_));
 INVx2_ASAP7_75t_R _24904_ (.A(_02550_),
    .Y(_02560_));
 INVx2_ASAP7_75t_SL _24905_ (.A(_02433_),
    .Y(_02561_));
 OAI22x1_ASAP7_75t_R _24906_ (.A1(_02559_),
    .A2(_02560_),
    .B1(_02441_),
    .B2(_02561_),
    .Y(_02562_));
 AND2x2_ASAP7_75t_R _24907_ (.A(_02562_),
    .B(_02388_),
    .Y(_02563_));
 NAND2x1p5_ASAP7_75t_SL _24908_ (.A(_02507_),
    .B(_02354_),
    .Y(_02564_));
 AND3x1_ASAP7_75t_L _24909_ (.A(_02480_),
    .B(_02564_),
    .C(_02372_),
    .Y(_02565_));
 NAND2x1_ASAP7_75t_R _24910_ (.A(_01236_),
    .B(_02357_),
    .Y(_02566_));
 AO21x1_ASAP7_75t_R _24911_ (.A1(_02428_),
    .A2(_02566_),
    .B(_02388_),
    .Y(_02567_));
 OAI21x1_ASAP7_75t_R _24912_ (.A1(_02565_),
    .A2(_02567_),
    .B(_02420_),
    .Y(_02568_));
 NAND2x1_ASAP7_75t_SL _24913_ (.A(_02378_),
    .B(_02478_),
    .Y(_02569_));
 NOR2x1p5_ASAP7_75t_L _24914_ (.A(_02429_),
    .B(_02354_),
    .Y(_02570_));
 NAND2x1_ASAP7_75t_R _24915_ (.A(_02372_),
    .B(_02570_),
    .Y(_02571_));
 NAND3x1_ASAP7_75t_SL _24916_ (.A(_02569_),
    .B(_02388_),
    .C(_02571_),
    .Y(_02572_));
 AOI21x1_ASAP7_75t_SL _24917_ (.A1(_02354_),
    .A2(_02429_),
    .B(_02372_),
    .Y(_02573_));
 NAND2x1_ASAP7_75t_L _24918_ (.A(_02545_),
    .B(_02573_),
    .Y(_02574_));
 NAND2x1_ASAP7_75t_SL _24919_ (.A(_02396_),
    .B(_02372_),
    .Y(_02575_));
 OA21x2_ASAP7_75t_R _24920_ (.A1(_02575_),
    .A2(_02354_),
    .B(_02389_),
    .Y(_02576_));
 AOI21x1_ASAP7_75t_R _24921_ (.A1(_02574_),
    .A2(_02576_),
    .B(_02420_),
    .Y(_02577_));
 AOI21x1_ASAP7_75t_R _24923_ (.A1(_02572_),
    .A2(_02577_),
    .B(_02493_),
    .Y(_02579_));
 OAI21x1_ASAP7_75t_R _24924_ (.A1(_02563_),
    .A2(_02568_),
    .B(_02579_),
    .Y(_02580_));
 NOR2x1_ASAP7_75t_SL _24925_ (.A(_02372_),
    .B(_02360_),
    .Y(_02581_));
 AOI21x1_ASAP7_75t_R _24926_ (.A1(_01234_),
    .A2(_02581_),
    .B(_02388_),
    .Y(_02582_));
 AOI21x1_ASAP7_75t_SL _24927_ (.A1(_02360_),
    .A2(_01233_),
    .B(_02379_),
    .Y(_02583_));
 NAND2x1_ASAP7_75t_SL _24928_ (.A(_02537_),
    .B(_02583_),
    .Y(_02584_));
 AOI21x1_ASAP7_75t_R _24929_ (.A1(_02582_),
    .A2(_02584_),
    .B(_02420_),
    .Y(_02585_));
 NOR2x1_ASAP7_75t_SL _24930_ (.A(_02360_),
    .B(_01236_),
    .Y(_02586_));
 NAND2x1_ASAP7_75t_SL _24931_ (.A(_02354_),
    .B(_01236_),
    .Y(_02587_));
 AOI21x1_ASAP7_75t_SL _24932_ (.A1(_01235_),
    .A2(_02360_),
    .B(_02379_),
    .Y(_02588_));
 AOI21x1_ASAP7_75t_R _24933_ (.A1(_02587_),
    .A2(_02588_),
    .B(_02389_),
    .Y(_02589_));
 OAI21x1_ASAP7_75t_R _24934_ (.A1(_02586_),
    .A2(_02441_),
    .B(_02589_),
    .Y(_02590_));
 AOI21x1_ASAP7_75t_R _24935_ (.A1(_02585_),
    .A2(_02590_),
    .B(_02525_),
    .Y(_02591_));
 INVx1_ASAP7_75t_SL _24936_ (.A(_02460_),
    .Y(_02592_));
 NAND2x1_ASAP7_75t_SL _24937_ (.A(_02379_),
    .B(_02377_),
    .Y(_02593_));
 OAI21x1_ASAP7_75t_R _24938_ (.A1(_02592_),
    .A2(_02593_),
    .B(_02499_),
    .Y(_02594_));
 INVx1_ASAP7_75t_SL _24939_ (.A(_02378_),
    .Y(_02595_));
 NAND2x1_ASAP7_75t_R _24940_ (.A(_02372_),
    .B(_02595_),
    .Y(_02596_));
 AND2x2_ASAP7_75t_R _24941_ (.A(_02379_),
    .B(_01249_),
    .Y(_02597_));
 AOI211x1_ASAP7_75t_R _24942_ (.A1(_02561_),
    .A2(_02372_),
    .B(_02389_),
    .C(_02597_),
    .Y(_02598_));
 AOI21x1_ASAP7_75t_R _24943_ (.A1(_02596_),
    .A2(_02598_),
    .B(_02444_),
    .Y(_02599_));
 NAND2x1_ASAP7_75t_R _24944_ (.A(_02594_),
    .B(_02599_),
    .Y(_02600_));
 AOI21x1_ASAP7_75t_R _24945_ (.A1(_02591_),
    .A2(_02600_),
    .B(_02451_),
    .Y(_02601_));
 NAND2x1_ASAP7_75t_R _24946_ (.A(_02580_),
    .B(_02601_),
    .Y(_02602_));
 AOI21x1_ASAP7_75t_SL _24947_ (.A1(_02456_),
    .A2(_02354_),
    .B(_02372_),
    .Y(_02603_));
 AOI21x1_ASAP7_75t_R _24949_ (.A1(_02402_),
    .A2(_02362_),
    .B(_02379_),
    .Y(_02605_));
 NAND2x1_ASAP7_75t_R _24950_ (.A(_02388_),
    .B(_02444_),
    .Y(_02606_));
 AOI211x1_ASAP7_75t_R _24951_ (.A1(_02431_),
    .A2(_02603_),
    .B(_02605_),
    .C(_02606_),
    .Y(_02607_));
 AO21x1_ASAP7_75t_R _24952_ (.A1(_02360_),
    .A2(_01235_),
    .B(_02372_),
    .Y(_02608_));
 OAI21x1_ASAP7_75t_R _24953_ (.A1(_02463_),
    .A2(_02608_),
    .B(_02388_),
    .Y(_02609_));
 AO21x1_ASAP7_75t_SL _24954_ (.A1(_02538_),
    .A2(_02546_),
    .B(_02444_),
    .Y(_02610_));
 NOR2x1_ASAP7_75t_R _24955_ (.A(_02609_),
    .B(_02610_),
    .Y(_02611_));
 INVx1_ASAP7_75t_R _24956_ (.A(_01247_),
    .Y(_02612_));
 NAND2x1_ASAP7_75t_R _24957_ (.A(_02379_),
    .B(_02420_),
    .Y(_02613_));
 OAI21x1_ASAP7_75t_R _24958_ (.A1(_02612_),
    .A2(_02613_),
    .B(_02389_),
    .Y(_02614_));
 INVx1_ASAP7_75t_R _24959_ (.A(_02363_),
    .Y(_02615_));
 OAI21x1_ASAP7_75t_R _24960_ (.A1(_02615_),
    .A2(_02570_),
    .B(_02372_),
    .Y(_02616_));
 INVx1_ASAP7_75t_R _24961_ (.A(_02616_),
    .Y(_02617_));
 OAI21x1_ASAP7_75t_R _24962_ (.A1(_02614_),
    .A2(_02617_),
    .B(_02493_),
    .Y(_02618_));
 NOR3x1_ASAP7_75t_R _24963_ (.A(_02607_),
    .B(_02611_),
    .C(_02618_),
    .Y(_02619_));
 AOI21x1_ASAP7_75t_R _24964_ (.A1(_01232_),
    .A2(_02354_),
    .B(_02379_),
    .Y(_02620_));
 INVx1_ASAP7_75t_R _24965_ (.A(_02620_),
    .Y(_02621_));
 AOI21x1_ASAP7_75t_R _24966_ (.A1(_02545_),
    .A2(_02573_),
    .B(_02389_),
    .Y(_02622_));
 OAI21x1_ASAP7_75t_R _24967_ (.A1(_02592_),
    .A2(_02621_),
    .B(_02622_),
    .Y(_02623_));
 NAND2x1_ASAP7_75t_R _24968_ (.A(_02431_),
    .B(_02474_),
    .Y(_02624_));
 AND2x2_ASAP7_75t_L _24969_ (.A(_02441_),
    .B(_02389_),
    .Y(_02625_));
 AOI21x1_ASAP7_75t_R _24970_ (.A1(_02624_),
    .A2(_02625_),
    .B(_02444_),
    .Y(_02626_));
 NAND2x1_ASAP7_75t_R _24971_ (.A(_02623_),
    .B(_02626_),
    .Y(_02627_));
 NOR2x2_ASAP7_75t_SL _24972_ (.A(_02360_),
    .B(_02426_),
    .Y(_02628_));
 AOI21x1_ASAP7_75t_SL _24973_ (.A1(_02372_),
    .A2(_02628_),
    .B(_02389_),
    .Y(_02629_));
 AOI21x1_ASAP7_75t_SL _24974_ (.A1(_02550_),
    .A2(_02564_),
    .B(_02372_),
    .Y(_02630_));
 NOR2x1_ASAP7_75t_L _24975_ (.A(_02515_),
    .B(_02630_),
    .Y(_02631_));
 NAND2x1_ASAP7_75t_L _24976_ (.A(_02629_),
    .B(_02631_),
    .Y(_02632_));
 NAND2x1_ASAP7_75t_R _24977_ (.A(_02501_),
    .B(_02354_),
    .Y(_02633_));
 AOI21x1_ASAP7_75t_R _24978_ (.A1(_02633_),
    .A2(_02538_),
    .B(_02388_),
    .Y(_02634_));
 NAND2x1_ASAP7_75t_SL _24979_ (.A(_02354_),
    .B(_02357_),
    .Y(_02635_));
 NAND2x1_ASAP7_75t_SL _24980_ (.A(_02635_),
    .B(_02398_),
    .Y(_02636_));
 AOI21x1_ASAP7_75t_R _24981_ (.A1(_02634_),
    .A2(_02636_),
    .B(_02420_),
    .Y(_02637_));
 NAND2x1_ASAP7_75t_R _24982_ (.A(_02632_),
    .B(_02637_),
    .Y(_02638_));
 AOI21x1_ASAP7_75t_R _24983_ (.A1(_02627_),
    .A2(_02638_),
    .B(_02493_),
    .Y(_02639_));
 OAI21x1_ASAP7_75t_SL _24984_ (.A1(_02619_),
    .A2(_02639_),
    .B(_02451_),
    .Y(_02640_));
 NAND2x1_ASAP7_75t_SL _24985_ (.A(_02602_),
    .B(_02640_),
    .Y(_00097_));
 OR2x2_ASAP7_75t_R _24987_ (.A(_02379_),
    .B(_01245_),
    .Y(_02642_));
 AO21x1_ASAP7_75t_SL _24988_ (.A1(_02497_),
    .A2(_02564_),
    .B(_02372_),
    .Y(_02643_));
 AOI21x1_ASAP7_75t_R _24989_ (.A1(_02642_),
    .A2(_02643_),
    .B(_02388_),
    .Y(_02644_));
 NOR2x1_ASAP7_75t_R _24990_ (.A(_02372_),
    .B(_02426_),
    .Y(_02645_));
 OAI21x1_ASAP7_75t_SL _24991_ (.A1(_02581_),
    .A2(_02645_),
    .B(_02635_),
    .Y(_02646_));
 AOI21x1_ASAP7_75t_R _24993_ (.A1(_02646_),
    .A2(_02382_),
    .B(_02389_),
    .Y(_02648_));
 NOR2x1_ASAP7_75t_L _24994_ (.A(_02644_),
    .B(_02648_),
    .Y(_02649_));
 NAND2x2_ASAP7_75t_SL _24995_ (.A(_02360_),
    .B(_01233_),
    .Y(_02650_));
 AOI21x1_ASAP7_75t_R _24996_ (.A1(_02426_),
    .A2(_02357_),
    .B(_02372_),
    .Y(_02651_));
 NOR2x1_ASAP7_75t_R _24997_ (.A(_02612_),
    .B(_02379_),
    .Y(_02652_));
 AOI21x1_ASAP7_75t_R _24998_ (.A1(_02650_),
    .A2(_02651_),
    .B(_02652_),
    .Y(_02653_));
 AOI21x1_ASAP7_75t_R _24999_ (.A1(_02389_),
    .A2(_02653_),
    .B(_02444_),
    .Y(_02654_));
 AND2x2_ASAP7_75t_SL _25000_ (.A(_02583_),
    .B(_02402_),
    .Y(_02655_));
 AO21x1_ASAP7_75t_SL _25001_ (.A1(_02507_),
    .A2(_02354_),
    .B(_02372_),
    .Y(_02656_));
 NOR2x1_ASAP7_75t_R _25002_ (.A(_02529_),
    .B(_02656_),
    .Y(_02657_));
 OAI21x1_ASAP7_75t_R _25004_ (.A1(_02655_),
    .A2(_02657_),
    .B(_02388_),
    .Y(_02659_));
 NAND2x1_ASAP7_75t_SL _25005_ (.A(_02654_),
    .B(_02659_),
    .Y(_02660_));
 OAI21x1_ASAP7_75t_R _25006_ (.A1(_02420_),
    .A2(_02649_),
    .B(_02660_),
    .Y(_02661_));
 NAND2x1_ASAP7_75t_SL _25007_ (.A(_02372_),
    .B(_02560_),
    .Y(_02662_));
 NOR2x1_ASAP7_75t_R _25008_ (.A(_01231_),
    .B(_02354_),
    .Y(_02663_));
 OAI21x1_ASAP7_75t_R _25009_ (.A1(_02561_),
    .A2(_02663_),
    .B(_02379_),
    .Y(_02664_));
 AOI21x1_ASAP7_75t_R _25010_ (.A1(_02662_),
    .A2(_02664_),
    .B(_02388_),
    .Y(_02665_));
 AND2x2_ASAP7_75t_R _25011_ (.A(_01232_),
    .B(_01235_),
    .Y(_02666_));
 NAND2x1_ASAP7_75t_SL _25012_ (.A(_02666_),
    .B(_02360_),
    .Y(_02667_));
 NAND2x1_ASAP7_75t_R _25013_ (.A(_02667_),
    .B(_02573_),
    .Y(_02668_));
 AOI21x1_ASAP7_75t_R _25014_ (.A1(_02668_),
    .A2(_02616_),
    .B(_02389_),
    .Y(_02669_));
 OAI21x1_ASAP7_75t_R _25015_ (.A1(_02665_),
    .A2(_02669_),
    .B(_02444_),
    .Y(_02670_));
 OA21x2_ASAP7_75t_R _25016_ (.A1(_01250_),
    .A2(_02379_),
    .B(_02388_),
    .Y(_02671_));
 NAND2x1_ASAP7_75t_R _25017_ (.A(_02650_),
    .B(_02603_),
    .Y(_02672_));
 AOI21x1_ASAP7_75t_R _25018_ (.A1(_02671_),
    .A2(_02672_),
    .B(_02444_),
    .Y(_02673_));
 AND2x2_ASAP7_75t_R _25019_ (.A(_02379_),
    .B(_01244_),
    .Y(_02674_));
 NOR2x1_ASAP7_75t_SL _25020_ (.A(_02674_),
    .B(_02481_),
    .Y(_02675_));
 NAND2x1_ASAP7_75t_R _25021_ (.A(_02389_),
    .B(_02675_),
    .Y(_02676_));
 AOI21x1_ASAP7_75t_R _25022_ (.A1(_02673_),
    .A2(_02676_),
    .B(_02525_),
    .Y(_02677_));
 AOI21x1_ASAP7_75t_SL _25023_ (.A1(_02670_),
    .A2(_02677_),
    .B(_02451_),
    .Y(_02678_));
 OAI21x1_ASAP7_75t_R _25024_ (.A1(_02493_),
    .A2(_02661_),
    .B(_02678_),
    .Y(_02679_));
 OAI21x1_ASAP7_75t_R _25026_ (.A1(_02663_),
    .A2(_02463_),
    .B(_02372_),
    .Y(_02681_));
 NOR2x1_ASAP7_75t_R _25027_ (.A(_01232_),
    .B(_02360_),
    .Y(_02682_));
 INVx1_ASAP7_75t_SL _25028_ (.A(_02362_),
    .Y(_02683_));
 OAI21x1_ASAP7_75t_R _25029_ (.A1(_02682_),
    .A2(_02683_),
    .B(_02379_),
    .Y(_02684_));
 NAND2x1_ASAP7_75t_SL _25030_ (.A(_02681_),
    .B(_02684_),
    .Y(_02685_));
 NAND2x1_ASAP7_75t_SL _25031_ (.A(_02460_),
    .B(_02573_),
    .Y(_02686_));
 AOI21x1_ASAP7_75t_R _25032_ (.A1(_02372_),
    .A2(_02457_),
    .B(_02388_),
    .Y(_02687_));
 AOI21x1_ASAP7_75t_R _25033_ (.A1(_02686_),
    .A2(_02687_),
    .B(_02420_),
    .Y(_02688_));
 OAI21x1_ASAP7_75t_SL _25034_ (.A1(_02389_),
    .A2(_02685_),
    .B(_02688_),
    .Y(_02689_));
 NAND2x1_ASAP7_75t_R _25035_ (.A(_02379_),
    .B(_02497_),
    .Y(_02690_));
 OAI21x1_ASAP7_75t_SL _25036_ (.A1(_02561_),
    .A2(_02690_),
    .B(_02389_),
    .Y(_02691_));
 NOR2x1_ASAP7_75t_R _25037_ (.A(_02381_),
    .B(_02691_),
    .Y(_02692_));
 NAND2x1_ASAP7_75t_R _25038_ (.A(_01240_),
    .B(_02354_),
    .Y(_02693_));
 NAND2x1_ASAP7_75t_R _25039_ (.A(_02693_),
    .B(_02588_),
    .Y(_02694_));
 AOI21x1_ASAP7_75t_R _25040_ (.A1(_02672_),
    .A2(_02694_),
    .B(_02389_),
    .Y(_02695_));
 OAI21x1_ASAP7_75t_R _25041_ (.A1(_02692_),
    .A2(_02695_),
    .B(_02420_),
    .Y(_02696_));
 AOI21x1_ASAP7_75t_R _25042_ (.A1(_02689_),
    .A2(_02696_),
    .B(_02525_),
    .Y(_02697_));
 AOI21x1_ASAP7_75t_R _25043_ (.A1(_01235_),
    .A2(_02354_),
    .B(_02372_),
    .Y(_02698_));
 NAND2x1_ASAP7_75t_R _25044_ (.A(_02378_),
    .B(_02698_),
    .Y(_02699_));
 AOI21x1_ASAP7_75t_R _25045_ (.A1(_02699_),
    .A2(_02439_),
    .B(_02388_),
    .Y(_02700_));
 NAND2x1_ASAP7_75t_R _25046_ (.A(_02480_),
    .B(_02698_),
    .Y(_02701_));
 INVx2_ASAP7_75t_R _25047_ (.A(_02437_),
    .Y(_02702_));
 NOR2x1_ASAP7_75t_SL _25048_ (.A(_01240_),
    .B(_02360_),
    .Y(_02703_));
 OAI21x1_ASAP7_75t_R _25050_ (.A1(_02702_),
    .A2(_02703_),
    .B(_02372_),
    .Y(_02705_));
 AOI21x1_ASAP7_75t_R _25051_ (.A1(_02701_),
    .A2(_02705_),
    .B(_02389_),
    .Y(_02706_));
 OAI21x1_ASAP7_75t_R _25052_ (.A1(_02700_),
    .A2(_02706_),
    .B(_02420_),
    .Y(_02707_));
 OAI21x1_ASAP7_75t_SL _25053_ (.A1(_02360_),
    .A2(_01233_),
    .B(_02379_),
    .Y(_02708_));
 NOR2x1_ASAP7_75t_R _25054_ (.A(_02702_),
    .B(_02708_),
    .Y(_02709_));
 OAI21x1_ASAP7_75t_R _25055_ (.A1(_02354_),
    .A2(_02426_),
    .B(_02372_),
    .Y(_02710_));
 OAI21x1_ASAP7_75t_R _25056_ (.A1(_02703_),
    .A2(_02710_),
    .B(_02388_),
    .Y(_02711_));
 NOR2x1_ASAP7_75t_R _25057_ (.A(_02709_),
    .B(_02711_),
    .Y(_02712_));
 AOI21x1_ASAP7_75t_R _25058_ (.A1(_01238_),
    .A2(_02354_),
    .B(_02379_),
    .Y(_02713_));
 NAND2x1_ASAP7_75t_SL _25059_ (.A(_02480_),
    .B(_02713_),
    .Y(_02714_));
 NAND3x1_ASAP7_75t_L _25060_ (.A(_02564_),
    .B(_02379_),
    .C(_02440_),
    .Y(_02715_));
 AOI21x1_ASAP7_75t_R _25061_ (.A1(_02714_),
    .A2(_02715_),
    .B(_02388_),
    .Y(_02716_));
 OAI21x1_ASAP7_75t_R _25062_ (.A1(_02712_),
    .A2(_02716_),
    .B(_02444_),
    .Y(_02717_));
 AOI21x1_ASAP7_75t_R _25063_ (.A1(_02707_),
    .A2(_02717_),
    .B(_02493_),
    .Y(_02718_));
 OAI21x1_ASAP7_75t_R _25064_ (.A1(_02697_),
    .A2(_02718_),
    .B(_02451_),
    .Y(_02719_));
 NAND2x1_ASAP7_75t_SL _25065_ (.A(_02679_),
    .B(_02719_),
    .Y(_00098_));
 NAND2x1_ASAP7_75t_SL _25066_ (.A(_02420_),
    .B(_02711_),
    .Y(_02720_));
 NOR2x1_ASAP7_75t_R _25067_ (.A(_02666_),
    .B(_02354_),
    .Y(_02721_));
 OAI21x1_ASAP7_75t_R _25068_ (.A1(_02513_),
    .A2(_02721_),
    .B(_02379_),
    .Y(_02722_));
 AOI21x1_ASAP7_75t_SL _25069_ (.A1(_02616_),
    .A2(_02722_),
    .B(_02388_),
    .Y(_02723_));
 OAI21x1_ASAP7_75t_SL _25070_ (.A1(_02720_),
    .A2(_02723_),
    .B(_02525_),
    .Y(_02724_));
 AOI21x1_ASAP7_75t_R _25071_ (.A1(_02502_),
    .A2(_02428_),
    .B(_02388_),
    .Y(_02725_));
 NAND2x1_ASAP7_75t_SL _25072_ (.A(_02584_),
    .B(_02725_),
    .Y(_02726_));
 OAI21x1_ASAP7_75t_SL _25073_ (.A1(_02702_),
    .A2(_02586_),
    .B(_02379_),
    .Y(_02727_));
 AOI21x1_ASAP7_75t_R _25074_ (.A1(_02693_),
    .A2(_02533_),
    .B(_02389_),
    .Y(_02728_));
 NAND2x1_ASAP7_75t_SL _25075_ (.A(_02727_),
    .B(_02728_),
    .Y(_02729_));
 AOI21x1_ASAP7_75t_SL _25076_ (.A1(_02726_),
    .A2(_02729_),
    .B(_02420_),
    .Y(_02730_));
 NOR2x1_ASAP7_75t_SL _25077_ (.A(_02724_),
    .B(_02730_),
    .Y(_02731_));
 INVx1_ASAP7_75t_R _25078_ (.A(_02478_),
    .Y(_02732_));
 INVx1_ASAP7_75t_SL _25079_ (.A(_02667_),
    .Y(_02733_));
 NAND2x1_ASAP7_75t_SL _25080_ (.A(_02440_),
    .B(_02474_),
    .Y(_02734_));
 OAI21x1_ASAP7_75t_SL _25081_ (.A1(_02732_),
    .A2(_02733_),
    .B(_02734_),
    .Y(_02735_));
 OA21x2_ASAP7_75t_SL _25082_ (.A1(_02437_),
    .A2(_02372_),
    .B(_02444_),
    .Y(_02736_));
 AOI21x1_ASAP7_75t_SL _25083_ (.A1(_02714_),
    .A2(_02736_),
    .B(_02388_),
    .Y(_02737_));
 OAI21x1_ASAP7_75t_SL _25084_ (.A1(_02444_),
    .A2(_02735_),
    .B(_02737_),
    .Y(_02738_));
 NAND2x1_ASAP7_75t_SL _25085_ (.A(_02528_),
    .B(_02354_),
    .Y(_02739_));
 AND3x1_ASAP7_75t_SL _25086_ (.A(_02583_),
    .B(_02739_),
    .C(_02420_),
    .Y(_02740_));
 OR3x1_ASAP7_75t_SL _25087_ (.A(_02440_),
    .B(_02379_),
    .C(_02420_),
    .Y(_02741_));
 NOR2x1_ASAP7_75t_R _25088_ (.A(_02377_),
    .B(_02613_),
    .Y(_02742_));
 NOR2x1_ASAP7_75t_SL _25089_ (.A(_02742_),
    .B(_02521_),
    .Y(_02743_));
 NAND2x1_ASAP7_75t_SL _25090_ (.A(_02741_),
    .B(_02743_),
    .Y(_02744_));
 OAI21x1_ASAP7_75t_SL _25091_ (.A1(_02740_),
    .A2(_02744_),
    .B(_02388_),
    .Y(_02745_));
 AOI21x1_ASAP7_75t_SL _25092_ (.A1(_02738_),
    .A2(_02745_),
    .B(_02525_),
    .Y(_02746_));
 OAI21x1_ASAP7_75t_SL _25093_ (.A1(_02731_),
    .A2(_02746_),
    .B(_02451_),
    .Y(_02747_));
 INVx2_ASAP7_75t_SL _25094_ (.A(_02440_),
    .Y(_02748_));
 NOR2x1_ASAP7_75t_R _25095_ (.A(_01236_),
    .B(_01233_),
    .Y(_02749_));
 OAI21x1_ASAP7_75t_SL _25096_ (.A1(_02628_),
    .A2(_02749_),
    .B(_02372_),
    .Y(_02750_));
 OAI21x1_ASAP7_75t_SL _25097_ (.A1(_02748_),
    .A2(_02708_),
    .B(_02750_),
    .Y(_02751_));
 AOI21x1_ASAP7_75t_R _25098_ (.A1(_02354_),
    .A2(_02357_),
    .B(_02379_),
    .Y(_02752_));
 NAND2x1_ASAP7_75t_SL _25099_ (.A(_02480_),
    .B(_02752_),
    .Y(_02753_));
 AOI21x1_ASAP7_75t_SL _25100_ (.A1(_02548_),
    .A2(_02753_),
    .B(_02444_),
    .Y(_02754_));
 OAI21x1_ASAP7_75t_SL _25101_ (.A1(_02388_),
    .A2(_02751_),
    .B(_02754_),
    .Y(_02755_));
 NOR2x1_ASAP7_75t_SL _25102_ (.A(_02560_),
    .B(_02593_),
    .Y(_02756_));
 NOR2x1_ASAP7_75t_SL _25103_ (.A(_02529_),
    .B(_02559_),
    .Y(_02757_));
 OAI21x1_ASAP7_75t_SL _25104_ (.A1(_02756_),
    .A2(_02757_),
    .B(_02388_),
    .Y(_02758_));
 NAND2x1_ASAP7_75t_SL _25105_ (.A(_02460_),
    .B(_02698_),
    .Y(_02759_));
 AOI21x1_ASAP7_75t_SL _25106_ (.A1(_02545_),
    .A2(_02752_),
    .B(_02388_),
    .Y(_02760_));
 AOI21x1_ASAP7_75t_SL _25107_ (.A1(_02759_),
    .A2(_02760_),
    .B(_02420_),
    .Y(_02761_));
 NAND2x1_ASAP7_75t_SL _25108_ (.A(_02758_),
    .B(_02761_),
    .Y(_02762_));
 AOI21x1_ASAP7_75t_SL _25109_ (.A1(_02755_),
    .A2(_02762_),
    .B(_02525_),
    .Y(_02763_));
 NAND2x1_ASAP7_75t_SL _25110_ (.A(_02545_),
    .B(_02713_),
    .Y(_02764_));
 AOI21x1_ASAP7_75t_SL _25111_ (.A1(_02569_),
    .A2(_02764_),
    .B(_02389_),
    .Y(_02765_));
 INVx1_ASAP7_75t_SL _25112_ (.A(_02603_),
    .Y(_02766_));
 AOI21x1_ASAP7_75t_SL _25113_ (.A1(_02766_),
    .A2(_02750_),
    .B(_02388_),
    .Y(_02767_));
 OAI21x1_ASAP7_75t_SL _25114_ (.A1(_02765_),
    .A2(_02767_),
    .B(_02420_),
    .Y(_02768_));
 AO21x1_ASAP7_75t_SL _25115_ (.A1(_02363_),
    .A2(_02440_),
    .B(_02379_),
    .Y(_02769_));
 NOR2x1_ASAP7_75t_R _25116_ (.A(_01236_),
    .B(_02357_),
    .Y(_02770_));
 OAI21x1_ASAP7_75t_SL _25117_ (.A1(_02628_),
    .A2(_02770_),
    .B(_02379_),
    .Y(_02771_));
 AOI21x1_ASAP7_75t_SL _25118_ (.A1(_02769_),
    .A2(_02771_),
    .B(_02389_),
    .Y(_02772_));
 OAI21x1_ASAP7_75t_SL _25119_ (.A1(_02468_),
    .A2(_02529_),
    .B(_02379_),
    .Y(_02773_));
 NOR2x1_ASAP7_75t_SL _25120_ (.A(_01231_),
    .B(_02360_),
    .Y(_02774_));
 OAI21x1_ASAP7_75t_SL _25121_ (.A1(_02774_),
    .A2(_02570_),
    .B(_02372_),
    .Y(_02775_));
 AOI21x1_ASAP7_75t_SL _25122_ (.A1(_02773_),
    .A2(_02775_),
    .B(_02388_),
    .Y(_02776_));
 OAI21x1_ASAP7_75t_SL _25123_ (.A1(_02772_),
    .A2(_02776_),
    .B(_02444_),
    .Y(_02777_));
 AOI21x1_ASAP7_75t_SL _25124_ (.A1(_02768_),
    .A2(_02777_),
    .B(_02493_),
    .Y(_02778_));
 OAI21x1_ASAP7_75t_SL _25125_ (.A1(_02763_),
    .A2(_02778_),
    .B(_02485_),
    .Y(_02779_));
 NAND2x1_ASAP7_75t_SL _25126_ (.A(_02747_),
    .B(_02779_),
    .Y(_00099_));
 NOR2x1_ASAP7_75t_R _25127_ (.A(_02360_),
    .B(_02357_),
    .Y(_02780_));
 OAI21x1_ASAP7_75t_R _25128_ (.A1(_02560_),
    .A2(_02780_),
    .B(_02379_),
    .Y(_02781_));
 AOI21x1_ASAP7_75t_R _25129_ (.A1(_02781_),
    .A2(_02499_),
    .B(_02444_),
    .Y(_02782_));
 AOI21x1_ASAP7_75t_SL _25130_ (.A1(_02456_),
    .A2(_02360_),
    .B(_02372_),
    .Y(_02783_));
 NAND2x1_ASAP7_75t_R _25131_ (.A(_02635_),
    .B(_02783_),
    .Y(_02784_));
 NAND3x1_ASAP7_75t_SL _25132_ (.A(_02694_),
    .B(_02784_),
    .C(_02388_),
    .Y(_02785_));
 NAND2x1_ASAP7_75t_SL _25133_ (.A(_02782_),
    .B(_02785_),
    .Y(_02786_));
 OAI21x1_ASAP7_75t_R _25134_ (.A1(_02702_),
    .A2(_02774_),
    .B(_02379_),
    .Y(_02787_));
 AOI21x1_ASAP7_75t_R _25135_ (.A1(_02439_),
    .A2(_02787_),
    .B(_02389_),
    .Y(_02788_));
 NOR2x1_ASAP7_75t_R _25136_ (.A(_01240_),
    .B(_02354_),
    .Y(_02789_));
 OAI21x1_ASAP7_75t_R _25137_ (.A1(_02774_),
    .A2(_02789_),
    .B(_02372_),
    .Y(_02790_));
 AOI21x1_ASAP7_75t_SL _25138_ (.A1(_02514_),
    .A2(_02790_),
    .B(_02388_),
    .Y(_02791_));
 OAI21x1_ASAP7_75t_R _25139_ (.A1(_02788_),
    .A2(_02791_),
    .B(_02444_),
    .Y(_02792_));
 NAND2x1_ASAP7_75t_R _25140_ (.A(_02786_),
    .B(_02792_),
    .Y(_02793_));
 OAI21x1_ASAP7_75t_R _25141_ (.A1(_02525_),
    .A2(_02793_),
    .B(_02485_),
    .Y(_02794_));
 NOR2x1_ASAP7_75t_SL _25142_ (.A(_02463_),
    .B(_02770_),
    .Y(_02795_));
 NAND2x1_ASAP7_75t_SL _25143_ (.A(_02372_),
    .B(_02795_),
    .Y(_02796_));
 AO21x1_ASAP7_75t_R _25144_ (.A1(_02378_),
    .A2(_02633_),
    .B(_02372_),
    .Y(_02797_));
 AO21x1_ASAP7_75t_R _25145_ (.A1(_02796_),
    .A2(_02797_),
    .B(_02389_),
    .Y(_02798_));
 INVx1_ASAP7_75t_SL _25146_ (.A(_02650_),
    .Y(_02799_));
 OAI21x1_ASAP7_75t_SL _25147_ (.A1(_01236_),
    .A2(_01233_),
    .B(_02379_),
    .Y(_02800_));
 OAI21x1_ASAP7_75t_R _25148_ (.A1(_02799_),
    .A2(_02800_),
    .B(_02389_),
    .Y(_02801_));
 NOR2x1_ASAP7_75t_R _25149_ (.A(_02780_),
    .B(_02710_),
    .Y(_02802_));
 OA21x2_ASAP7_75t_R _25150_ (.A1(_02801_),
    .A2(_02802_),
    .B(_02420_),
    .Y(_02803_));
 AO21x1_ASAP7_75t_R _25151_ (.A1(_02354_),
    .A2(_01238_),
    .B(_02372_),
    .Y(_02804_));
 AO21x1_ASAP7_75t_R _25152_ (.A1(_02804_),
    .A2(_02401_),
    .B(_02389_),
    .Y(_02805_));
 AOI21x1_ASAP7_75t_SL _25153_ (.A1(_02354_),
    .A2(_01233_),
    .B(_02372_),
    .Y(_02806_));
 AND2x2_ASAP7_75t_SL _25154_ (.A(_02806_),
    .B(_02480_),
    .Y(_02807_));
 OAI21x1_ASAP7_75t_R _25155_ (.A1(_02605_),
    .A2(_02807_),
    .B(_02389_),
    .Y(_02808_));
 AOI21x1_ASAP7_75t_R _25156_ (.A1(_02805_),
    .A2(_02808_),
    .B(_02420_),
    .Y(_02809_));
 AOI211x1_ASAP7_75t_R _25157_ (.A1(_02798_),
    .A2(_02803_),
    .B(_02809_),
    .C(_02493_),
    .Y(_02810_));
 INVx1_ASAP7_75t_R _25158_ (.A(_02404_),
    .Y(_02811_));
 INVx1_ASAP7_75t_R _25159_ (.A(_02541_),
    .Y(_02812_));
 OAI21x1_ASAP7_75t_R _25160_ (.A1(_02811_),
    .A2(_02812_),
    .B(_02389_),
    .Y(_02813_));
 NOR2x1_ASAP7_75t_R _25161_ (.A(_02683_),
    .B(_02804_),
    .Y(_02814_));
 INVx1_ASAP7_75t_R _25162_ (.A(_02796_),
    .Y(_02815_));
 OAI21x1_ASAP7_75t_R _25163_ (.A1(_02814_),
    .A2(_02815_),
    .B(_02388_),
    .Y(_02816_));
 AOI21x1_ASAP7_75t_R _25164_ (.A1(_02813_),
    .A2(_02816_),
    .B(_02525_),
    .Y(_02817_));
 AND3x1_ASAP7_75t_R _25165_ (.A(_02546_),
    .B(_02372_),
    .C(_02502_),
    .Y(_02818_));
 NOR2x1_ASAP7_75t_R _25166_ (.A(_02818_),
    .B(_02609_),
    .Y(_02819_));
 AO21x1_ASAP7_75t_R _25167_ (.A1(_02538_),
    .A2(_02693_),
    .B(_02581_),
    .Y(_02820_));
 OAI21x1_ASAP7_75t_R _25168_ (.A1(_02388_),
    .A2(_02820_),
    .B(_02525_),
    .Y(_02821_));
 OAI21x1_ASAP7_75t_R _25169_ (.A1(_02819_),
    .A2(_02821_),
    .B(_02420_),
    .Y(_02822_));
 OAI21x1_ASAP7_75t_R _25170_ (.A1(_02595_),
    .A2(_02804_),
    .B(_02519_),
    .Y(_02823_));
 OA21x2_ASAP7_75t_SL _25171_ (.A1(_02429_),
    .A2(_02379_),
    .B(_02389_),
    .Y(_02824_));
 AOI21x1_ASAP7_75t_R _25172_ (.A1(_02656_),
    .A2(_02824_),
    .B(_02525_),
    .Y(_02825_));
 AOI21x1_ASAP7_75t_R _25173_ (.A1(_02823_),
    .A2(_02825_),
    .B(_02420_),
    .Y(_02826_));
 INVx1_ASAP7_75t_SL _25174_ (.A(_02465_),
    .Y(_02827_));
 AND2x2_ASAP7_75t_R _25175_ (.A(_02588_),
    .B(_02564_),
    .Y(_02828_));
 NOR2x1_ASAP7_75t_SL _25176_ (.A(_02389_),
    .B(_02573_),
    .Y(_02829_));
 AOI21x1_ASAP7_75t_R _25177_ (.A1(_02621_),
    .A2(_02829_),
    .B(_02493_),
    .Y(_02830_));
 OAI21x1_ASAP7_75t_R _25178_ (.A1(_02827_),
    .A2(_02828_),
    .B(_02830_),
    .Y(_02831_));
 AOI21x1_ASAP7_75t_R _25179_ (.A1(_02826_),
    .A2(_02831_),
    .B(_02485_),
    .Y(_02832_));
 OAI21x1_ASAP7_75t_SL _25180_ (.A1(_02817_),
    .A2(_02822_),
    .B(_02832_),
    .Y(_02833_));
 OAI21x1_ASAP7_75t_SL _25181_ (.A1(_02794_),
    .A2(_02810_),
    .B(_02833_),
    .Y(_00100_));
 INVx1_ASAP7_75t_SL _25182_ (.A(_02739_),
    .Y(_02834_));
 OAI21x1_ASAP7_75t_SL _25183_ (.A1(_02748_),
    .A2(_02703_),
    .B(_02372_),
    .Y(_02835_));
 OAI21x1_ASAP7_75t_SL _25184_ (.A1(_02834_),
    .A2(_02441_),
    .B(_02835_),
    .Y(_02836_));
 NOR2x1_ASAP7_75t_R _25185_ (.A(_02528_),
    .B(_02372_),
    .Y(_02837_));
 AOI21x1_ASAP7_75t_SL _25186_ (.A1(_02372_),
    .A2(_02431_),
    .B(_02837_),
    .Y(_02838_));
 AOI21x1_ASAP7_75t_SL _25187_ (.A1(_02389_),
    .A2(_02838_),
    .B(_02444_),
    .Y(_02839_));
 OAI21x1_ASAP7_75t_SL _25188_ (.A1(_02389_),
    .A2(_02836_),
    .B(_02839_),
    .Y(_02840_));
 AO21x1_ASAP7_75t_SL _25189_ (.A1(_02561_),
    .A2(_02372_),
    .B(_02389_),
    .Y(_02841_));
 AOI21x1_ASAP7_75t_SL _25190_ (.A1(_02379_),
    .A2(_02667_),
    .B(_02388_),
    .Y(_02842_));
 OAI21x1_ASAP7_75t_SL _25191_ (.A1(_02468_),
    .A2(_02570_),
    .B(_02372_),
    .Y(_02843_));
 AOI21x1_ASAP7_75t_SL _25192_ (.A1(_02842_),
    .A2(_02843_),
    .B(_02420_),
    .Y(_02844_));
 OAI21x1_ASAP7_75t_SL _25193_ (.A1(_02478_),
    .A2(_02841_),
    .B(_02844_),
    .Y(_02845_));
 AOI21x1_ASAP7_75t_SL _25194_ (.A1(_02840_),
    .A2(_02845_),
    .B(_02525_),
    .Y(_02846_));
 OA21x2_ASAP7_75t_SL _25195_ (.A1(_02683_),
    .A2(_02561_),
    .B(_02372_),
    .Y(_02847_));
 OA21x2_ASAP7_75t_SL _25196_ (.A1(_02363_),
    .A2(_02372_),
    .B(_02388_),
    .Y(_02848_));
 OAI21x1_ASAP7_75t_SL _25197_ (.A1(_02570_),
    .A2(_02703_),
    .B(_02372_),
    .Y(_02849_));
 AOI21x1_ASAP7_75t_SL _25198_ (.A1(_02848_),
    .A2(_02849_),
    .B(_02444_),
    .Y(_02850_));
 OAI21x1_ASAP7_75t_SL _25199_ (.A1(_02827_),
    .A2(_02847_),
    .B(_02850_),
    .Y(_02851_));
 NAND2x1_ASAP7_75t_SL _25200_ (.A(_02378_),
    .B(_02713_),
    .Y(_02852_));
 NAND2x1_ASAP7_75t_SL _25201_ (.A(_02440_),
    .B(_02603_),
    .Y(_02853_));
 AOI21x1_ASAP7_75t_SL _25202_ (.A1(_02852_),
    .A2(_02853_),
    .B(_02389_),
    .Y(_02854_));
 AOI21x1_ASAP7_75t_SL _25203_ (.A1(_02537_),
    .A2(_02538_),
    .B(_02645_),
    .Y(_02855_));
 NOR2x1_ASAP7_75t_SL _25204_ (.A(_02388_),
    .B(_02855_),
    .Y(_02856_));
 OAI21x1_ASAP7_75t_SL _25205_ (.A1(_02854_),
    .A2(_02856_),
    .B(_02444_),
    .Y(_02857_));
 AOI21x1_ASAP7_75t_SL _25206_ (.A1(_02851_),
    .A2(_02857_),
    .B(_02493_),
    .Y(_02858_));
 OAI21x1_ASAP7_75t_SL _25207_ (.A1(_02846_),
    .A2(_02858_),
    .B(_02451_),
    .Y(_02859_));
 OAI21x1_ASAP7_75t_SL _25208_ (.A1(_02379_),
    .A2(_02703_),
    .B(_02389_),
    .Y(_02860_));
 NOR2x1_ASAP7_75t_SL _25209_ (.A(_02530_),
    .B(_02441_),
    .Y(_02861_));
 NOR2x1_ASAP7_75t_SL _25210_ (.A(_02860_),
    .B(_02861_),
    .Y(_02862_));
 NAND2x1_ASAP7_75t_SL _25211_ (.A(_02379_),
    .B(_02774_),
    .Y(_02863_));
 NAND2x1_ASAP7_75t_SL _25212_ (.A(_02650_),
    .B(_02620_),
    .Y(_02864_));
 AOI21x1_ASAP7_75t_SL _25213_ (.A1(_02863_),
    .A2(_02864_),
    .B(_02389_),
    .Y(_02865_));
 OAI21x1_ASAP7_75t_SL _25214_ (.A1(_02862_),
    .A2(_02865_),
    .B(_02420_),
    .Y(_02866_));
 AO21x1_ASAP7_75t_SL _25215_ (.A1(_02357_),
    .A2(_02379_),
    .B(_02388_),
    .Y(_02867_));
 AOI21x1_ASAP7_75t_SL _25216_ (.A1(_02372_),
    .A2(_02795_),
    .B(_02867_),
    .Y(_02868_));
 OAI21x1_ASAP7_75t_SL _25217_ (.A1(_02615_),
    .A2(_02570_),
    .B(_02379_),
    .Y(_02869_));
 NOR2x1_ASAP7_75t_R _25218_ (.A(_02426_),
    .B(_02357_),
    .Y(_02870_));
 OAI21x1_ASAP7_75t_SL _25219_ (.A1(_02586_),
    .A2(_02870_),
    .B(_02372_),
    .Y(_02871_));
 AOI21x1_ASAP7_75t_SL _25220_ (.A1(_02869_),
    .A2(_02871_),
    .B(_02389_),
    .Y(_02872_));
 OAI21x1_ASAP7_75t_SL _25221_ (.A1(_02868_),
    .A2(_02872_),
    .B(_02444_),
    .Y(_02873_));
 AOI21x1_ASAP7_75t_SL _25222_ (.A1(_02866_),
    .A2(_02873_),
    .B(_02525_),
    .Y(_02874_));
 OR3x1_ASAP7_75t_SL _25223_ (.A(_02588_),
    .B(_02389_),
    .C(_02468_),
    .Y(_02875_));
 NOR2x1_ASAP7_75t_SL _25224_ (.A(_02388_),
    .B(_02533_),
    .Y(_02876_));
 AOI21x1_ASAP7_75t_SL _25225_ (.A1(_02727_),
    .A2(_02876_),
    .B(_02444_),
    .Y(_02877_));
 NAND2x1_ASAP7_75t_SL _25226_ (.A(_02875_),
    .B(_02877_),
    .Y(_02878_));
 INVx1_ASAP7_75t_R _25227_ (.A(_02666_),
    .Y(_02879_));
 NAND2x1_ASAP7_75t_SL _25228_ (.A(_02879_),
    .B(_02698_),
    .Y(_02880_));
 OAI21x1_ASAP7_75t_SL _25229_ (.A1(_02512_),
    .A2(_02513_),
    .B(_02372_),
    .Y(_02881_));
 AOI21x1_ASAP7_75t_SL _25230_ (.A1(_02880_),
    .A2(_02881_),
    .B(_02389_),
    .Y(_02882_));
 OAI21x1_ASAP7_75t_SL _25231_ (.A1(_02703_),
    .A2(_02470_),
    .B(_02379_),
    .Y(_02883_));
 AOI21x1_ASAP7_75t_SL _25232_ (.A1(_02883_),
    .A2(_02464_),
    .B(_02388_),
    .Y(_02884_));
 OAI21x1_ASAP7_75t_SL _25233_ (.A1(_02882_),
    .A2(_02884_),
    .B(_02444_),
    .Y(_02885_));
 AOI21x1_ASAP7_75t_SL _25234_ (.A1(_02878_),
    .A2(_02885_),
    .B(_02493_),
    .Y(_02886_));
 OAI21x1_ASAP7_75t_SL _25235_ (.A1(_02874_),
    .A2(_02886_),
    .B(_02485_),
    .Y(_02887_));
 NAND2x1_ASAP7_75t_SL _25236_ (.A(_02859_),
    .B(_02887_),
    .Y(_00101_));
 NOR2x1_ASAP7_75t_R _25237_ (.A(_02389_),
    .B(_02520_),
    .Y(_02888_));
 OAI21x1_ASAP7_75t_SL _25238_ (.A1(_02512_),
    .A2(_02463_),
    .B(_02379_),
    .Y(_02889_));
 AOI21x1_ASAP7_75t_SL _25239_ (.A1(_02888_),
    .A2(_02889_),
    .B(_02525_),
    .Y(_02890_));
 AOI21x1_ASAP7_75t_SL _25240_ (.A1(_02587_),
    .A2(_02783_),
    .B(_02388_),
    .Y(_02891_));
 OAI21x1_ASAP7_75t_SL _25241_ (.A1(_02508_),
    .A2(_02733_),
    .B(_02891_),
    .Y(_02892_));
 AOI21x1_ASAP7_75t_SL _25242_ (.A1(_02890_),
    .A2(_02892_),
    .B(_02451_),
    .Y(_02893_));
 AOI21x1_ASAP7_75t_SL _25243_ (.A1(_02460_),
    .A2(_02713_),
    .B(_02388_),
    .Y(_02894_));
 OAI21x1_ASAP7_75t_SL _25244_ (.A1(_02358_),
    .A2(_02359_),
    .B(_01239_),
    .Y(_02895_));
 AO21x1_ASAP7_75t_SL _25245_ (.A1(_02401_),
    .A2(_02895_),
    .B(_02372_),
    .Y(_02896_));
 AOI21x1_ASAP7_75t_SL _25246_ (.A1(_02894_),
    .A2(_02896_),
    .B(_02493_),
    .Y(_02897_));
 OA21x2_ASAP7_75t_SL _25247_ (.A1(_02437_),
    .A2(_02372_),
    .B(_02388_),
    .Y(_02898_));
 AOI22x1_ASAP7_75t_SL _25248_ (.A1(_02581_),
    .A2(_02879_),
    .B1(_02538_),
    .B2(_02564_),
    .Y(_02899_));
 NAND2x1_ASAP7_75t_SL _25249_ (.A(_02898_),
    .B(_02899_),
    .Y(_02900_));
 NAND2x1_ASAP7_75t_SL _25250_ (.A(_02897_),
    .B(_02900_),
    .Y(_02901_));
 AOI21x1_ASAP7_75t_SL _25251_ (.A1(_02893_),
    .A2(_02901_),
    .B(_02444_),
    .Y(_02902_));
 OAI21x1_ASAP7_75t_SL _25252_ (.A1(_02513_),
    .A2(_02799_),
    .B(_02379_),
    .Y(_02903_));
 OAI21x1_ASAP7_75t_SL _25253_ (.A1(_02379_),
    .A2(_02834_),
    .B(_02903_),
    .Y(_02904_));
 NAND2x1_ASAP7_75t_SL _25254_ (.A(_02493_),
    .B(_02691_),
    .Y(_02905_));
 AOI21x1_ASAP7_75t_SL _25255_ (.A1(_02388_),
    .A2(_02904_),
    .B(_02905_),
    .Y(_02906_));
 NAND2x1_ASAP7_75t_SL _25256_ (.A(_02372_),
    .B(_02663_),
    .Y(_02907_));
 NAND3x1_ASAP7_75t_SL _25257_ (.A(_02727_),
    .B(_02389_),
    .C(_02907_),
    .Y(_02908_));
 INVx1_ASAP7_75t_SL _25258_ (.A(_02597_),
    .Y(_02909_));
 NAND2x1_ASAP7_75t_SL _25259_ (.A(_02909_),
    .B(_02483_),
    .Y(_02910_));
 AOI21x1_ASAP7_75t_SL _25260_ (.A1(_02908_),
    .A2(_02910_),
    .B(_02493_),
    .Y(_02911_));
 OAI21x1_ASAP7_75t_SL _25261_ (.A1(_02906_),
    .A2(_02911_),
    .B(_02451_),
    .Y(_02912_));
 NAND2x1_ASAP7_75t_SL _25262_ (.A(_02902_),
    .B(_02912_),
    .Y(_02913_));
 NAND2x1_ASAP7_75t_SL _25263_ (.A(_02545_),
    .B(_02620_),
    .Y(_02914_));
 NAND2x1_ASAP7_75t_SL _25264_ (.A(_02378_),
    .B(_02603_),
    .Y(_02915_));
 AOI21x1_ASAP7_75t_SL _25265_ (.A1(_02914_),
    .A2(_02915_),
    .B(_02388_),
    .Y(_02916_));
 AO21x1_ASAP7_75t_SL _25266_ (.A1(_02748_),
    .A2(_02372_),
    .B(_02389_),
    .Y(_02917_));
 OAI21x1_ASAP7_75t_SL _25267_ (.A1(_02917_),
    .A2(_02675_),
    .B(_02493_),
    .Y(_02918_));
 NOR2x1_ASAP7_75t_SL _25268_ (.A(_02916_),
    .B(_02918_),
    .Y(_02919_));
 OAI21x1_ASAP7_75t_SL _25269_ (.A1(_02870_),
    .A2(_02595_),
    .B(_02379_),
    .Y(_02920_));
 AO21x1_ASAP7_75t_R _25270_ (.A1(_01248_),
    .A2(_01242_),
    .B(_02379_),
    .Y(_02921_));
 AND2x2_ASAP7_75t_SL _25271_ (.A(_02921_),
    .B(_02389_),
    .Y(_02922_));
 NAND2x1_ASAP7_75t_SL _25272_ (.A(_02920_),
    .B(_02922_),
    .Y(_02923_));
 NAND2x1_ASAP7_75t_SL _25273_ (.A(_02400_),
    .B(_02581_),
    .Y(_02924_));
 NAND3x1_ASAP7_75t_SL _25274_ (.A(_02898_),
    .B(_02662_),
    .C(_02924_),
    .Y(_02925_));
 AOI21x1_ASAP7_75t_SL _25275_ (.A1(_02923_),
    .A2(_02925_),
    .B(_02493_),
    .Y(_02926_));
 OAI21x1_ASAP7_75t_SL _25276_ (.A1(_02919_),
    .A2(_02926_),
    .B(_02485_),
    .Y(_02927_));
 AO21x1_ASAP7_75t_SL _25277_ (.A1(_01243_),
    .A2(_02379_),
    .B(_02388_),
    .Y(_02928_));
 AO21x1_ASAP7_75t_SL _25278_ (.A1(_02378_),
    .A2(_02713_),
    .B(_02928_),
    .Y(_02929_));
 OAI21x1_ASAP7_75t_SL _25279_ (.A1(_02748_),
    .A2(_02703_),
    .B(_02379_),
    .Y(_02930_));
 AOI21x1_ASAP7_75t_SL _25280_ (.A1(_02930_),
    .A2(_02629_),
    .B(_02525_),
    .Y(_02931_));
 AOI21x1_ASAP7_75t_SL _25281_ (.A1(_02929_),
    .A2(_02931_),
    .B(_02485_),
    .Y(_02932_));
 AO21x1_ASAP7_75t_SL _25282_ (.A1(_02360_),
    .A2(_01240_),
    .B(_02379_),
    .Y(_02933_));
 AOI211x1_ASAP7_75t_SL _25283_ (.A1(_02933_),
    .A2(_02800_),
    .B(_02389_),
    .C(_02628_),
    .Y(_02934_));
 OAI21x1_ASAP7_75t_SL _25284_ (.A1(_02468_),
    .A2(_02595_),
    .B(_02372_),
    .Y(_02935_));
 AO21x1_ASAP7_75t_SL _25285_ (.A1(_02537_),
    .A2(_02587_),
    .B(_02372_),
    .Y(_02936_));
 AOI21x1_ASAP7_75t_SL _25286_ (.A1(_02935_),
    .A2(_02936_),
    .B(_02388_),
    .Y(_02937_));
 OAI21x1_ASAP7_75t_SL _25287_ (.A1(_02934_),
    .A2(_02937_),
    .B(_02525_),
    .Y(_02938_));
 AOI21x1_ASAP7_75t_SL _25288_ (.A1(_02932_),
    .A2(_02938_),
    .B(_02420_),
    .Y(_02939_));
 NAND2x1_ASAP7_75t_SL _25289_ (.A(_02927_),
    .B(_02939_),
    .Y(_02940_));
 NAND2x1_ASAP7_75t_SL _25290_ (.A(_02913_),
    .B(_02940_),
    .Y(_00102_));
 NOR2x1_ASAP7_75t_SL _25291_ (.A(_02379_),
    .B(_01236_),
    .Y(_02941_));
 OAI21x1_ASAP7_75t_SL _25292_ (.A1(_02941_),
    .A2(_02807_),
    .B(_02388_),
    .Y(_02942_));
 AO21x1_ASAP7_75t_SL _25293_ (.A1(_02650_),
    .A2(_02895_),
    .B(_02379_),
    .Y(_02943_));
 INVx1_ASAP7_75t_SL _25294_ (.A(_02801_),
    .Y(_02944_));
 AOI21x1_ASAP7_75t_SL _25295_ (.A1(_02943_),
    .A2(_02944_),
    .B(_02525_),
    .Y(_02945_));
 NAND2x1_ASAP7_75t_SL _25296_ (.A(_02942_),
    .B(_02945_),
    .Y(_02946_));
 AOI21x1_ASAP7_75t_SL _25297_ (.A1(_02502_),
    .A2(_02573_),
    .B(_02389_),
    .Y(_02947_));
 AO21x1_ASAP7_75t_SL _25298_ (.A1(_02587_),
    .A2(_02497_),
    .B(_02379_),
    .Y(_02948_));
 NAND2x1_ASAP7_75t_SL _25299_ (.A(_02947_),
    .B(_02948_),
    .Y(_02949_));
 AND2x2_ASAP7_75t_SL _25300_ (.A(_02933_),
    .B(_02389_),
    .Y(_02950_));
 AOI21x1_ASAP7_75t_SL _25301_ (.A1(_02903_),
    .A2(_02950_),
    .B(_02493_),
    .Y(_02951_));
 AOI21x1_ASAP7_75t_SL _25302_ (.A1(_02949_),
    .A2(_02951_),
    .B(_02485_),
    .Y(_02952_));
 NAND2x1_ASAP7_75t_SL _25303_ (.A(_02946_),
    .B(_02952_),
    .Y(_02953_));
 AO21x1_ASAP7_75t_SL _25304_ (.A1(_01239_),
    .A2(_02379_),
    .B(_02388_),
    .Y(_02954_));
 OA21x2_ASAP7_75t_SL _25305_ (.A1(_02503_),
    .A2(_02954_),
    .B(_02493_),
    .Y(_02955_));
 AOI21x1_ASAP7_75t_SL _25306_ (.A1(_02372_),
    .A2(_02463_),
    .B(_02518_),
    .Y(_02956_));
 NAND2x1_ASAP7_75t_SL _25307_ (.A(_02636_),
    .B(_02956_),
    .Y(_02957_));
 AOI21x1_ASAP7_75t_SL _25308_ (.A1(_02955_),
    .A2(_02957_),
    .B(_02451_),
    .Y(_02958_));
 AND2x2_ASAP7_75t_SL _25309_ (.A(_02583_),
    .B(_02532_),
    .Y(_02959_));
 NAND2x1_ASAP7_75t_SL _25310_ (.A(_02388_),
    .B(_02722_),
    .Y(_02960_));
 AOI21x1_ASAP7_75t_R _25311_ (.A1(_02363_),
    .A2(_02440_),
    .B(_02372_),
    .Y(_02961_));
 AOI21x1_ASAP7_75t_SL _25312_ (.A1(_02895_),
    .A2(_02550_),
    .B(_02379_),
    .Y(_02962_));
 NOR2x1_ASAP7_75t_SL _25313_ (.A(_02961_),
    .B(_02962_),
    .Y(_02963_));
 AOI21x1_ASAP7_75t_SL _25314_ (.A1(_02389_),
    .A2(_02963_),
    .B(_02493_),
    .Y(_02964_));
 OAI21x1_ASAP7_75t_SL _25315_ (.A1(_02959_),
    .A2(_02960_),
    .B(_02964_),
    .Y(_02965_));
 AOI21x1_ASAP7_75t_SL _25316_ (.A1(_02958_),
    .A2(_02965_),
    .B(_02420_),
    .Y(_02966_));
 NAND2x1_ASAP7_75t_SL _25317_ (.A(_02953_),
    .B(_02966_),
    .Y(_02967_));
 NOR2x1_ASAP7_75t_SL _25318_ (.A(_01248_),
    .B(_02372_),
    .Y(_02968_));
 AOI21x1_ASAP7_75t_SL _25319_ (.A1(_02377_),
    .A2(_02437_),
    .B(_02379_),
    .Y(_02969_));
 OAI21x1_ASAP7_75t_SL _25320_ (.A1(_02968_),
    .A2(_02969_),
    .B(_02389_),
    .Y(_02970_));
 NAND2x1_ASAP7_75t_SL _25321_ (.A(_02493_),
    .B(_02970_),
    .Y(_02971_));
 NOR2x1_ASAP7_75t_SL _25322_ (.A(_02774_),
    .B(_02441_),
    .Y(_02972_));
 AOI211x1_ASAP7_75t_SL _25323_ (.A1(_02583_),
    .A2(_02587_),
    .B(_02972_),
    .C(_02389_),
    .Y(_02973_));
 NOR2x1_ASAP7_75t_SL _25324_ (.A(_02971_),
    .B(_02973_),
    .Y(_02974_));
 NAND2x1_ASAP7_75t_SL _25325_ (.A(_02389_),
    .B(_02502_),
    .Y(_02975_));
 NOR2x1_ASAP7_75t_SL _25326_ (.A(_02620_),
    .B(_02806_),
    .Y(_02976_));
 OAI21x1_ASAP7_75t_SL _25327_ (.A1(_02975_),
    .A2(_02976_),
    .B(_02525_),
    .Y(_02977_));
 AOI21x1_ASAP7_75t_SL _25328_ (.A1(_02575_),
    .A2(_02920_),
    .B(_02389_),
    .Y(_02978_));
 OAI21x1_ASAP7_75t_SL _25329_ (.A1(_02977_),
    .A2(_02978_),
    .B(_02485_),
    .Y(_02979_));
 NOR2x1_ASAP7_75t_SL _25330_ (.A(_02974_),
    .B(_02979_),
    .Y(_02980_));
 NOR2x1_ASAP7_75t_SL _25331_ (.A(_02372_),
    .B(_02570_),
    .Y(_02981_));
 NOR3x1_ASAP7_75t_SL _25332_ (.A(_02981_),
    .B(_02388_),
    .C(_02533_),
    .Y(_02982_));
 AOI21x1_ASAP7_75t_SL _25333_ (.A1(_02440_),
    .A2(_02895_),
    .B(_02379_),
    .Y(_02983_));
 OA21x2_ASAP7_75t_SL _25334_ (.A1(_02983_),
    .A2(_02783_),
    .B(_02388_),
    .Y(_02984_));
 OAI21x1_ASAP7_75t_SL _25335_ (.A1(_02982_),
    .A2(_02984_),
    .B(_02493_),
    .Y(_02985_));
 OAI21x1_ASAP7_75t_SL _25336_ (.A1(_02592_),
    .A2(_02593_),
    .B(_02734_),
    .Y(_02986_));
 AOI21x1_ASAP7_75t_SL _25337_ (.A1(_02646_),
    .A2(_02894_),
    .B(_02493_),
    .Y(_02987_));
 OAI21x1_ASAP7_75t_SL _25338_ (.A1(_02389_),
    .A2(_02986_),
    .B(_02987_),
    .Y(_02988_));
 AOI21x1_ASAP7_75t_SL _25339_ (.A1(_02985_),
    .A2(_02988_),
    .B(_02485_),
    .Y(_02989_));
 OAI21x1_ASAP7_75t_SL _25340_ (.A1(_02980_),
    .A2(_02989_),
    .B(_02420_),
    .Y(_02990_));
 NAND2x1_ASAP7_75t_SL _25341_ (.A(_02967_),
    .B(_02990_),
    .Y(_00103_));
 NOR2x1p5_ASAP7_75t_L _25342_ (.A(_00574_),
    .B(_00471_),
    .Y(_02991_));
 XOR2x2_ASAP7_75t_SL _25343_ (.A(_00686_),
    .B(_00679_),
    .Y(_02992_));
 XOR2x2_ASAP7_75t_SL _25344_ (.A(_11392_),
    .B(_02992_),
    .Y(_02993_));
 XOR2x2_ASAP7_75t_SL _25345_ (.A(_14180_),
    .B(_11434_),
    .Y(_02994_));
 NAND2x1p5_ASAP7_75t_SL _25346_ (.A(_02994_),
    .B(_02993_),
    .Y(_02995_));
 XOR2x2_ASAP7_75t_SL _25347_ (.A(_00680_),
    .B(_02992_),
    .Y(_02996_));
 XOR2x2_ASAP7_75t_SL _25348_ (.A(_14180_),
    .B(_11426_),
    .Y(_02997_));
 NAND2x1p5_ASAP7_75t_L _25349_ (.A(_02996_),
    .B(_02997_),
    .Y(_02998_));
 AOI21x1_ASAP7_75t_SL _25350_ (.A1(_02998_),
    .A2(_02995_),
    .B(_10675_),
    .Y(_02999_));
 OAI21x1_ASAP7_75t_R _25351_ (.A1(_02991_),
    .A2(_02999_),
    .B(_00901_),
    .Y(_03000_));
 AND2x2_ASAP7_75t_R _25352_ (.A(_10675_),
    .B(_00471_),
    .Y(_03001_));
 NAND2x1p5_ASAP7_75t_SL _25353_ (.A(_02994_),
    .B(_02996_),
    .Y(_03002_));
 NAND2x1p5_ASAP7_75t_SL _25354_ (.A(_02997_),
    .B(_02993_),
    .Y(_03003_));
 AOI21x1_ASAP7_75t_SL _25355_ (.A1(_03003_),
    .A2(_03002_),
    .B(_10675_),
    .Y(_03004_));
 OAI21x1_ASAP7_75t_R _25356_ (.A1(_03001_),
    .A2(_03004_),
    .B(_08729_),
    .Y(_03005_));
 NAND2x2_ASAP7_75t_SL _25357_ (.A(_03005_),
    .B(_03000_),
    .Y(_01256_));
 NOR2x1p5_ASAP7_75t_L _25358_ (.A(_00574_),
    .B(_00472_),
    .Y(_03006_));
 XOR2x2_ASAP7_75t_SL _25359_ (.A(_00615_),
    .B(_00583_),
    .Y(_03007_));
 INVx1_ASAP7_75t_SL _25360_ (.A(_03007_),
    .Y(_03008_));
 NAND2x1p5_ASAP7_75t_L _25361_ (.A(_00654_),
    .B(_03008_),
    .Y(_03009_));
 INVx1_ASAP7_75t_R _25362_ (.A(_00654_),
    .Y(_03010_));
 NAND2x1_ASAP7_75t_L _25363_ (.A(_03010_),
    .B(_03007_),
    .Y(_03011_));
 INVx2_ASAP7_75t_L _25364_ (.A(_02992_),
    .Y(_03012_));
 NAND3x1_ASAP7_75t_R _25365_ (.A(_03009_),
    .B(_03011_),
    .C(_03012_),
    .Y(_03013_));
 AOI21x1_ASAP7_75t_SL _25366_ (.A1(_03011_),
    .A2(_03009_),
    .B(_03012_),
    .Y(_03014_));
 INVx1_ASAP7_75t_SL _25367_ (.A(_03014_),
    .Y(_03015_));
 AOI21x1_ASAP7_75t_SL _25368_ (.A1(_03013_),
    .A2(_03015_),
    .B(_10675_),
    .Y(_03016_));
 OAI21x1_ASAP7_75t_R _25369_ (.A1(_03006_),
    .A2(_03016_),
    .B(_00900_),
    .Y(_03017_));
 XOR2x2_ASAP7_75t_SL _25370_ (.A(_00654_),
    .B(_03007_),
    .Y(_03018_));
 NOR2x1_ASAP7_75t_L _25371_ (.A(_02992_),
    .B(_03018_),
    .Y(_03019_));
 OAI21x1_ASAP7_75t_SL _25372_ (.A1(_03019_),
    .A2(_03014_),
    .B(_00574_),
    .Y(_03020_));
 INVx1_ASAP7_75t_R _25373_ (.A(_00900_),
    .Y(_03021_));
 INVx2_ASAP7_75t_R _25374_ (.A(_03006_),
    .Y(_03022_));
 NAND3x1_ASAP7_75t_R _25375_ (.A(_03020_),
    .B(_03021_),
    .C(_03022_),
    .Y(_03023_));
 NAND2x2_ASAP7_75t_SL _25376_ (.A(_03017_),
    .B(_03023_),
    .Y(_01259_));
 NAND2x1_ASAP7_75t_R _25377_ (.A(_00473_),
    .B(_10675_),
    .Y(_03024_));
 XOR2x2_ASAP7_75t_SL _25378_ (.A(_00585_),
    .B(_00617_),
    .Y(_03025_));
 INVx2_ASAP7_75t_L _25379_ (.A(_03025_),
    .Y(_03026_));
 INVx1_ASAP7_75t_R _25380_ (.A(_00681_),
    .Y(_03027_));
 XOR2x2_ASAP7_75t_SL _25381_ (.A(_14181_),
    .B(_03027_),
    .Y(_03028_));
 NAND2x1_ASAP7_75t_SL _25382_ (.A(_03026_),
    .B(_03028_),
    .Y(_03029_));
 NOR2x1_ASAP7_75t_R _25383_ (.A(_03027_),
    .B(_14181_),
    .Y(_03030_));
 XNOR2x2_ASAP7_75t_L _25384_ (.A(_00648_),
    .B(_00680_),
    .Y(_03031_));
 NOR2x1_ASAP7_75t_R _25385_ (.A(_00681_),
    .B(_03031_),
    .Y(_03032_));
 OAI21x1_ASAP7_75t_SL _25386_ (.A1(_03030_),
    .A2(_03032_),
    .B(_03025_),
    .Y(_03033_));
 NAND3x1_ASAP7_75t_SL _25387_ (.A(_03029_),
    .B(_00574_),
    .C(_03033_),
    .Y(_03034_));
 AOI21x1_ASAP7_75t_SL _25388_ (.A1(_03024_),
    .A2(_03034_),
    .B(_00871_),
    .Y(_03035_));
 NOR2x1_ASAP7_75t_R _25389_ (.A(_00574_),
    .B(_00473_),
    .Y(_03036_));
 AOI21x1_ASAP7_75t_SL _25390_ (.A1(_03033_),
    .A2(_03029_),
    .B(_10675_),
    .Y(_03037_));
 OAI21x1_ASAP7_75t_SL _25391_ (.A1(_03036_),
    .A2(_03037_),
    .B(_00871_),
    .Y(_03038_));
 INVx2_ASAP7_75t_SL _25392_ (.A(_03038_),
    .Y(_03039_));
 NOR2x2_ASAP7_75t_SL _25393_ (.A(_03035_),
    .B(_03039_),
    .Y(_03040_));
 OAI21x1_ASAP7_75t_SL _25395_ (.A1(_02999_),
    .A2(_02991_),
    .B(_08729_),
    .Y(_03041_));
 OAI21x1_ASAP7_75t_SL _25396_ (.A1(_03004_),
    .A2(_03001_),
    .B(_00901_),
    .Y(_03042_));
 NAND2x1p5_ASAP7_75t_SL _25397_ (.A(_03042_),
    .B(_03041_),
    .Y(_03043_));
 INVx1_ASAP7_75t_R _25399_ (.A(_00871_),
    .Y(_03044_));
 AOI21x1_ASAP7_75t_SL _25400_ (.A1(_03024_),
    .A2(_03034_),
    .B(_03044_),
    .Y(_03045_));
 OAI21x1_ASAP7_75t_SL _25401_ (.A1(_03036_),
    .A2(_03037_),
    .B(_03044_),
    .Y(_03046_));
 INVx2_ASAP7_75t_SL _25402_ (.A(_03046_),
    .Y(_03047_));
 NOR2x1_ASAP7_75t_SL _25403_ (.A(_03045_),
    .B(_03047_),
    .Y(_03048_));
 OAI21x1_ASAP7_75t_SL _25406_ (.A1(_03016_),
    .A2(_03006_),
    .B(_03021_),
    .Y(_03050_));
 NAND3x1_ASAP7_75t_SL _25407_ (.A(_03022_),
    .B(_00900_),
    .C(_03020_),
    .Y(_03051_));
 NAND2x1p5_ASAP7_75t_SL _25408_ (.A(_03051_),
    .B(_03050_),
    .Y(_03052_));
 XNOR2x2_ASAP7_75t_SL _25411_ (.A(_00682_),
    .B(_14239_),
    .Y(_03054_));
 XNOR2x2_ASAP7_75t_L _25412_ (.A(_00681_),
    .B(_00686_),
    .Y(_03055_));
 XOR2x2_ASAP7_75t_R _25413_ (.A(_00586_),
    .B(_00618_),
    .Y(_03056_));
 XOR2x2_ASAP7_75t_L _25414_ (.A(_03055_),
    .B(_03056_),
    .Y(_03057_));
 AOI21x1_ASAP7_75t_R _25415_ (.A1(_03054_),
    .A2(_03057_),
    .B(_10675_),
    .Y(_03058_));
 OR2x2_ASAP7_75t_SL _25416_ (.A(_03057_),
    .B(_03054_),
    .Y(_03059_));
 AND2x2_ASAP7_75t_R _25417_ (.A(_10675_),
    .B(_00505_),
    .Y(_03060_));
 AOI21x1_ASAP7_75t_SL _25418_ (.A1(_03058_),
    .A2(_03059_),
    .B(_03060_),
    .Y(_03061_));
 XOR2x2_ASAP7_75t_SL _25419_ (.A(_03061_),
    .B(_00872_),
    .Y(_03062_));
 AOI21x1_ASAP7_75t_SL _25421_ (.A1(_03052_),
    .A2(_03040_),
    .B(_03062_),
    .Y(_03064_));
 INVx1_ASAP7_75t_SL _25422_ (.A(_01263_),
    .Y(_03065_));
 NOR2x1_ASAP7_75t_L _25423_ (.A(_03065_),
    .B(_03040_),
    .Y(_03066_));
 INVx1_ASAP7_75t_SL _25424_ (.A(_03066_),
    .Y(_03067_));
 INVx2_ASAP7_75t_R _25425_ (.A(_01257_),
    .Y(_03068_));
 NOR2x1_ASAP7_75t_L _25427_ (.A(_03068_),
    .B(_03048_),
    .Y(_03070_));
 NOR2x1_ASAP7_75t_SL _25428_ (.A(_03043_),
    .B(_03040_),
    .Y(_03071_));
 OA21x2_ASAP7_75t_R _25431_ (.A1(_03070_),
    .A2(_03071_),
    .B(_03062_),
    .Y(_03074_));
 XOR2x2_ASAP7_75t_R _25432_ (.A(_00682_),
    .B(_00686_),
    .Y(_03075_));
 XOR2x2_ASAP7_75t_SL _25433_ (.A(_11545_),
    .B(_03075_),
    .Y(_03076_));
 XNOR2x2_ASAP7_75t_SL _25434_ (.A(_14269_),
    .B(_03076_),
    .Y(_03077_));
 NOR2x1_ASAP7_75t_R _25435_ (.A(_00574_),
    .B(_00504_),
    .Y(_03078_));
 AOI21x1_ASAP7_75t_R _25436_ (.A1(_00574_),
    .A2(_03077_),
    .B(_03078_),
    .Y(_03079_));
 XNOR2x2_ASAP7_75t_SL _25437_ (.A(_00873_),
    .B(_03079_),
    .Y(_03080_));
 AOI211x1_ASAP7_75t_R _25440_ (.A1(_03064_),
    .A2(_03067_),
    .B(_03074_),
    .C(_03080_),
    .Y(_03083_));
 INVx1_ASAP7_75t_SL _25441_ (.A(_03080_),
    .Y(_03084_));
 INVx2_ASAP7_75t_R _25444_ (.A(_01262_),
    .Y(_03087_));
 NAND2x1_ASAP7_75t_R _25445_ (.A(_03087_),
    .B(_03048_),
    .Y(_03088_));
 NAND2x1_ASAP7_75t_SL _25446_ (.A(_03088_),
    .B(_03064_),
    .Y(_03089_));
 NAND2x2_ASAP7_75t_SL _25447_ (.A(_03043_),
    .B(_03040_),
    .Y(_03090_));
 INVx1_ASAP7_75t_SL _25448_ (.A(_01255_),
    .Y(_03091_));
 OAI21x1_ASAP7_75t_R _25449_ (.A1(_03035_),
    .A2(_03039_),
    .B(_03091_),
    .Y(_03092_));
 XNOR2x2_ASAP7_75t_SL _25450_ (.A(_00872_),
    .B(_03061_),
    .Y(_03093_));
 AO21x1_ASAP7_75t_SL _25453_ (.A1(_03090_),
    .A2(_03092_),
    .B(_03093_),
    .Y(_03096_));
 NAND2x1_ASAP7_75t_SL _25454_ (.A(_03089_),
    .B(_03096_),
    .Y(_03097_));
 XOR2x2_ASAP7_75t_SL _25455_ (.A(_00684_),
    .B(_00685_),
    .Y(_03098_));
 XOR2x2_ASAP7_75t_R _25456_ (.A(_03098_),
    .B(_00652_),
    .Y(_03099_));
 XOR2x2_ASAP7_75t_R _25457_ (.A(_03099_),
    .B(_11588_),
    .Y(_03100_));
 NOR2x1_ASAP7_75t_R _25458_ (.A(_00574_),
    .B(_00502_),
    .Y(_03101_));
 AO21x1_ASAP7_75t_R _25459_ (.A1(_03100_),
    .A2(_00574_),
    .B(_03101_),
    .Y(_03102_));
 XOR2x2_ASAP7_75t_SL _25460_ (.A(_03102_),
    .B(_00875_),
    .Y(_03103_));
 INVx2_ASAP7_75t_SL _25461_ (.A(_03103_),
    .Y(_03104_));
 OAI21x1_ASAP7_75t_R _25463_ (.A1(_03084_),
    .A2(_03097_),
    .B(_03104_),
    .Y(_03106_));
 NOR2x1_ASAP7_75t_L _25464_ (.A(_03083_),
    .B(_03106_),
    .Y(_03107_));
 AOI21x1_ASAP7_75t_SL _25469_ (.A1(_03040_),
    .A2(_01254_),
    .B(_03062_),
    .Y(_03112_));
 OAI21x1_ASAP7_75t_SL _25470_ (.A1(_03035_),
    .A2(_03039_),
    .B(_01254_),
    .Y(_03113_));
 AOI21x1_ASAP7_75t_R _25474_ (.A1(_03113_),
    .A2(_03090_),
    .B(_03093_),
    .Y(_03117_));
 OAI21x1_ASAP7_75t_R _25477_ (.A1(_03112_),
    .A2(_03117_),
    .B(_03084_),
    .Y(_03120_));
 NAND2x1_ASAP7_75t_R _25478_ (.A(_03103_),
    .B(_03120_),
    .Y(_03121_));
 INVx1_ASAP7_75t_R _25479_ (.A(_01253_),
    .Y(_03122_));
 NAND2x1_ASAP7_75t_R _25480_ (.A(_03122_),
    .B(_03040_),
    .Y(_03123_));
 NAND2x1p5_ASAP7_75t_SL _25481_ (.A(_03113_),
    .B(_03093_),
    .Y(_03124_));
 INVx2_ASAP7_75t_SL _25482_ (.A(_03124_),
    .Y(_03125_));
 OAI21x1_ASAP7_75t_R _25484_ (.A1(_03035_),
    .A2(_03039_),
    .B(_01253_),
    .Y(_03127_));
 NOR2x1_ASAP7_75t_L _25485_ (.A(_03093_),
    .B(_03127_),
    .Y(_03128_));
 NOR2x1_ASAP7_75t_SL _25486_ (.A(_03084_),
    .B(_03128_),
    .Y(_03129_));
 INVx1_ASAP7_75t_R _25487_ (.A(_03129_),
    .Y(_03130_));
 OAI21x1_ASAP7_75t_SL _25488_ (.A1(_03045_),
    .A2(_03047_),
    .B(_01260_),
    .Y(_03131_));
 NOR2x1_ASAP7_75t_R _25489_ (.A(_03093_),
    .B(_03131_),
    .Y(_03132_));
 AOI211x1_ASAP7_75t_R _25490_ (.A1(_03123_),
    .A2(_03125_),
    .B(_03130_),
    .C(_03132_),
    .Y(_03133_));
 NOR2x1_ASAP7_75t_R _25491_ (.A(_00574_),
    .B(_00503_),
    .Y(_03134_));
 XOR2x2_ASAP7_75t_R _25492_ (.A(_11503_),
    .B(_00684_),
    .Y(_03135_));
 XOR2x2_ASAP7_75t_SL _25493_ (.A(_03135_),
    .B(_11482_),
    .Y(_03136_));
 NOR2x1_ASAP7_75t_R _25494_ (.A(_10675_),
    .B(_03136_),
    .Y(_03137_));
 INVx1_ASAP7_75t_R _25495_ (.A(_00874_),
    .Y(_03138_));
 OAI21x1_ASAP7_75t_R _25496_ (.A1(_03134_),
    .A2(_03137_),
    .B(_03138_),
    .Y(_03139_));
 XNOR2x2_ASAP7_75t_R _25497_ (.A(_11482_),
    .B(_03135_),
    .Y(_03140_));
 NAND2x1_ASAP7_75t_R _25498_ (.A(_00574_),
    .B(_03140_),
    .Y(_03141_));
 INVx1_ASAP7_75t_R _25499_ (.A(_03134_),
    .Y(_03142_));
 NAND3x1_ASAP7_75t_SL _25500_ (.A(_03141_),
    .B(_00874_),
    .C(_03142_),
    .Y(_03143_));
 NAND2x2_ASAP7_75t_SL _25501_ (.A(_03139_),
    .B(_03143_),
    .Y(_03144_));
 OAI21x1_ASAP7_75t_R _25503_ (.A1(_03121_),
    .A2(_03133_),
    .B(_03144_),
    .Y(_03146_));
 NOR2x1_ASAP7_75t_L _25504_ (.A(_03107_),
    .B(_03146_),
    .Y(_03147_));
 INVx4_ASAP7_75t_SL _25505_ (.A(_01254_),
    .Y(_03148_));
 NAND2x2_ASAP7_75t_L _25506_ (.A(_03148_),
    .B(_03048_),
    .Y(_03149_));
 OAI21x1_ASAP7_75t_R _25507_ (.A1(_03045_),
    .A2(_03047_),
    .B(_01262_),
    .Y(_03150_));
 AO21x1_ASAP7_75t_R _25509_ (.A1(_03149_),
    .A2(_03150_),
    .B(_03093_),
    .Y(_03152_));
 NOR2x1_ASAP7_75t_R _25511_ (.A(_03122_),
    .B(_03048_),
    .Y(_03154_));
 INVx1_ASAP7_75t_R _25512_ (.A(_01260_),
    .Y(_03155_));
 NOR2x1_ASAP7_75t_SL _25513_ (.A(_03155_),
    .B(_03040_),
    .Y(_03156_));
 OAI21x1_ASAP7_75t_R _25514_ (.A1(_03154_),
    .A2(_03156_),
    .B(_03093_),
    .Y(_03157_));
 AND3x1_ASAP7_75t_R _25515_ (.A(_03152_),
    .B(_03080_),
    .C(_03157_),
    .Y(_03158_));
 NOR2x1_ASAP7_75t_R _25516_ (.A(_01256_),
    .B(_01259_),
    .Y(_03159_));
 OAI21x1_ASAP7_75t_R _25517_ (.A1(_03052_),
    .A2(_03040_),
    .B(_03062_),
    .Y(_03160_));
 NOR2x1_ASAP7_75t_R _25518_ (.A(_03159_),
    .B(_03160_),
    .Y(_03161_));
 NAND2x1_ASAP7_75t_R _25519_ (.A(_01259_),
    .B(_03048_),
    .Y(_03162_));
 NAND2x2_ASAP7_75t_SL _25520_ (.A(_03043_),
    .B(_03052_),
    .Y(_03163_));
 AO21x1_ASAP7_75t_R _25522_ (.A1(_03162_),
    .A2(_03163_),
    .B(_03062_),
    .Y(_03165_));
 NAND2x1_ASAP7_75t_R _25523_ (.A(_03084_),
    .B(_03165_),
    .Y(_03166_));
 OAI21x1_ASAP7_75t_R _25525_ (.A1(_03161_),
    .A2(_03166_),
    .B(_03103_),
    .Y(_03168_));
 NOR2x1_ASAP7_75t_R _25526_ (.A(_03158_),
    .B(_03168_),
    .Y(_03169_));
 NAND2x1_ASAP7_75t_L _25527_ (.A(_03052_),
    .B(_03048_),
    .Y(_03170_));
 AOI21x1_ASAP7_75t_SL _25528_ (.A1(_03068_),
    .A2(_03040_),
    .B(_03093_),
    .Y(_03171_));
 NAND2x1_ASAP7_75t_R _25529_ (.A(_03170_),
    .B(_03171_),
    .Y(_03172_));
 AOI21x1_ASAP7_75t_SL _25530_ (.A1(_01263_),
    .A2(_03040_),
    .B(_03062_),
    .Y(_03173_));
 NAND2x1_ASAP7_75t_R _25531_ (.A(_03113_),
    .B(_03173_),
    .Y(_03174_));
 AOI21x1_ASAP7_75t_R _25532_ (.A1(_03172_),
    .A2(_03174_),
    .B(_03080_),
    .Y(_03175_));
 AOI21x1_ASAP7_75t_SL _25533_ (.A1(_03052_),
    .A2(_03040_),
    .B(_03093_),
    .Y(_03176_));
 INVx1_ASAP7_75t_R _25534_ (.A(_03176_),
    .Y(_03177_));
 NOR2x1_ASAP7_75t_SL _25536_ (.A(_01258_),
    .B(_03040_),
    .Y(_03179_));
 OAI21x1_ASAP7_75t_R _25538_ (.A1(_03070_),
    .A2(_03179_),
    .B(_03093_),
    .Y(_03181_));
 AOI21x1_ASAP7_75t_R _25539_ (.A1(_03177_),
    .A2(_03181_),
    .B(_03084_),
    .Y(_03182_));
 NOR2x1_ASAP7_75t_R _25540_ (.A(_03175_),
    .B(_03182_),
    .Y(_03183_));
 INVx2_ASAP7_75t_SL _25541_ (.A(_03144_),
    .Y(_03184_));
 OAI21x1_ASAP7_75t_R _25543_ (.A1(_03103_),
    .A2(_03183_),
    .B(_03184_),
    .Y(_03186_));
 XOR2x2_ASAP7_75t_R _25544_ (.A(_14325_),
    .B(_11589_),
    .Y(_03187_));
 XOR2x2_ASAP7_75t_R _25545_ (.A(_03187_),
    .B(_11409_),
    .Y(_03188_));
 NOR2x1_ASAP7_75t_R _25546_ (.A(_00574_),
    .B(_00501_),
    .Y(_03189_));
 AO21x1_ASAP7_75t_R _25547_ (.A1(_03188_),
    .A2(_00574_),
    .B(_03189_),
    .Y(_03190_));
 XOR2x2_ASAP7_75t_R _25548_ (.A(_03190_),
    .B(_00876_),
    .Y(_03191_));
 OAI21x1_ASAP7_75t_R _25550_ (.A1(_03169_),
    .A2(_03186_),
    .B(_03191_),
    .Y(_03193_));
 AO21x1_ASAP7_75t_R _25551_ (.A1(_03048_),
    .A2(_01258_),
    .B(_03062_),
    .Y(_03194_));
 INVx1_ASAP7_75t_R _25552_ (.A(_03092_),
    .Y(_03195_));
 OAI21x1_ASAP7_75t_R _25554_ (.A1(_03195_),
    .A2(_03154_),
    .B(_03062_),
    .Y(_03197_));
 AOI21x1_ASAP7_75t_R _25555_ (.A1(_03194_),
    .A2(_03197_),
    .B(_03080_),
    .Y(_03198_));
 NAND2x1p5_ASAP7_75t_SL _25556_ (.A(_03148_),
    .B(_03040_),
    .Y(_03199_));
 AOI21x1_ASAP7_75t_SL _25557_ (.A1(_01256_),
    .A2(_03048_),
    .B(_03093_),
    .Y(_03200_));
 NAND2x1p5_ASAP7_75t_SL _25558_ (.A(_03200_),
    .B(_03199_),
    .Y(_03201_));
 INVx1_ASAP7_75t_R _25559_ (.A(_03131_),
    .Y(_03202_));
 NOR2x1_ASAP7_75t_R _25560_ (.A(_03052_),
    .B(_03040_),
    .Y(_03203_));
 OAI21x1_ASAP7_75t_R _25561_ (.A1(_03202_),
    .A2(_03203_),
    .B(_03093_),
    .Y(_03204_));
 AOI21x1_ASAP7_75t_R _25562_ (.A1(_03201_),
    .A2(_03204_),
    .B(_03084_),
    .Y(_03205_));
 OAI21x1_ASAP7_75t_R _25563_ (.A1(_03198_),
    .A2(_03205_),
    .B(_03104_),
    .Y(_03206_));
 NAND2x1_ASAP7_75t_R _25564_ (.A(_03062_),
    .B(_03195_),
    .Y(_03207_));
 NAND2x1_ASAP7_75t_R _25565_ (.A(_01261_),
    .B(_03040_),
    .Y(_03208_));
 AOI21x1_ASAP7_75t_R _25566_ (.A1(_03068_),
    .A2(_03048_),
    .B(_03062_),
    .Y(_03209_));
 AOI21x1_ASAP7_75t_R _25567_ (.A1(_03208_),
    .A2(_03209_),
    .B(_03084_),
    .Y(_03210_));
 NAND2x1_ASAP7_75t_SL _25568_ (.A(_03207_),
    .B(_03210_),
    .Y(_03211_));
 OAI21x1_ASAP7_75t_R _25569_ (.A1(_03035_),
    .A2(_03039_),
    .B(_01257_),
    .Y(_03212_));
 OA21x2_ASAP7_75t_R _25570_ (.A1(_03212_),
    .A2(_03093_),
    .B(_03084_),
    .Y(_03213_));
 NOR2x1_ASAP7_75t_R _25571_ (.A(_03062_),
    .B(_03092_),
    .Y(_03214_));
 NOR2x1_ASAP7_75t_R _25572_ (.A(_03132_),
    .B(_03214_),
    .Y(_03215_));
 AOI21x1_ASAP7_75t_R _25573_ (.A1(_03213_),
    .A2(_03215_),
    .B(_03104_),
    .Y(_03216_));
 AOI21x1_ASAP7_75t_R _25574_ (.A1(_03211_),
    .A2(_03216_),
    .B(_03144_),
    .Y(_03217_));
 AOI21x1_ASAP7_75t_R _25575_ (.A1(_03206_),
    .A2(_03217_),
    .B(_03191_),
    .Y(_03218_));
 OAI21x1_ASAP7_75t_R _25576_ (.A1(_03045_),
    .A2(_03047_),
    .B(_03091_),
    .Y(_03219_));
 INVx1_ASAP7_75t_R _25577_ (.A(_03219_),
    .Y(_03220_));
 NAND2x1_ASAP7_75t_R _25578_ (.A(_03062_),
    .B(_03220_),
    .Y(_03221_));
 NOR2x1_ASAP7_75t_R _25579_ (.A(_01253_),
    .B(_03040_),
    .Y(_03222_));
 INVx1_ASAP7_75t_R _25580_ (.A(_03222_),
    .Y(_03223_));
 NAND2x1_ASAP7_75t_SL _25581_ (.A(_03223_),
    .B(_03064_),
    .Y(_03224_));
 NAND2x1_ASAP7_75t_R _25582_ (.A(_03221_),
    .B(_03224_),
    .Y(_03225_));
 INVx1_ASAP7_75t_R _25583_ (.A(_01258_),
    .Y(_03226_));
 NAND2x1_ASAP7_75t_R _25584_ (.A(_03226_),
    .B(_03062_),
    .Y(_03227_));
 OA21x2_ASAP7_75t_SL _25585_ (.A1(_03227_),
    .A2(_03048_),
    .B(_03080_),
    .Y(_03228_));
 OAI21x1_ASAP7_75t_SL _25586_ (.A1(_03093_),
    .A2(_03212_),
    .B(_03228_),
    .Y(_03229_));
 AND2x2_ASAP7_75t_R _25587_ (.A(_03093_),
    .B(_01268_),
    .Y(_03230_));
 AO21x1_ASAP7_75t_R _25588_ (.A1(_03062_),
    .A2(_03199_),
    .B(_03230_),
    .Y(_03231_));
 AOI21x1_ASAP7_75t_R _25589_ (.A1(_03084_),
    .A2(_03231_),
    .B(_03104_),
    .Y(_03232_));
 OAI21x1_ASAP7_75t_R _25590_ (.A1(_03225_),
    .A2(_03229_),
    .B(_03232_),
    .Y(_03233_));
 NAND2x1_ASAP7_75t_R _25591_ (.A(_03089_),
    .B(_03228_),
    .Y(_03234_));
 OA21x2_ASAP7_75t_R _25592_ (.A1(_03227_),
    .A2(_03048_),
    .B(_03084_),
    .Y(_03235_));
 INVx1_ASAP7_75t_R _25593_ (.A(_03035_),
    .Y(_03236_));
 AOI21x1_ASAP7_75t_SL _25594_ (.A1(_03038_),
    .A2(_03236_),
    .B(_01261_),
    .Y(_03237_));
 INVx1_ASAP7_75t_R _25595_ (.A(_03237_),
    .Y(_03238_));
 OA21x2_ASAP7_75t_SL _25596_ (.A1(_03093_),
    .A2(_03238_),
    .B(_03124_),
    .Y(_03239_));
 AOI21x1_ASAP7_75t_R _25597_ (.A1(_03235_),
    .A2(_03239_),
    .B(_03103_),
    .Y(_03240_));
 AOI21x1_ASAP7_75t_R _25598_ (.A1(_03234_),
    .A2(_03240_),
    .B(_03184_),
    .Y(_03241_));
 NAND2x1_ASAP7_75t_R _25599_ (.A(_03233_),
    .B(_03241_),
    .Y(_03242_));
 NAND2x1_ASAP7_75t_SL _25600_ (.A(_03218_),
    .B(_03242_),
    .Y(_03243_));
 OAI21x1_ASAP7_75t_SL _25601_ (.A1(_03147_),
    .A2(_03193_),
    .B(_03243_),
    .Y(_00104_));
 INVx2_ASAP7_75t_SL _25602_ (.A(_03191_),
    .Y(_03244_));
 INVx2_ASAP7_75t_SL _25603_ (.A(_03090_),
    .Y(_03245_));
 NOR2x1_ASAP7_75t_R _25604_ (.A(_03245_),
    .B(_03194_),
    .Y(_03246_));
 INVx1_ASAP7_75t_SL _25605_ (.A(_03160_),
    .Y(_03247_));
 AO21x1_ASAP7_75t_R _25607_ (.A1(_03247_),
    .A2(_03123_),
    .B(_03084_),
    .Y(_03249_));
 NOR2x1_ASAP7_75t_R _25608_ (.A(_03246_),
    .B(_03249_),
    .Y(_03250_));
 OAI21x1_ASAP7_75t_SL _25609_ (.A1(_03045_),
    .A2(_03047_),
    .B(_01254_),
    .Y(_03251_));
 NAND2x1p5_ASAP7_75t_SL _25610_ (.A(_03251_),
    .B(_03093_),
    .Y(_03252_));
 NOR2x1_ASAP7_75t_R _25611_ (.A(_03222_),
    .B(_03252_),
    .Y(_03253_));
 NOR2x1_ASAP7_75t_SL _25612_ (.A(_03052_),
    .B(_03048_),
    .Y(_03254_));
 NAND2x1_ASAP7_75t_R _25613_ (.A(_03062_),
    .B(_03254_),
    .Y(_03255_));
 OA21x2_ASAP7_75t_R _25614_ (.A1(_03092_),
    .A2(_03093_),
    .B(_03084_),
    .Y(_03256_));
 NAND2x1_ASAP7_75t_R _25615_ (.A(_03255_),
    .B(_03256_),
    .Y(_03257_));
 OAI21x1_ASAP7_75t_R _25616_ (.A1(_03253_),
    .A2(_03257_),
    .B(_03184_),
    .Y(_03258_));
 OA21x2_ASAP7_75t_R _25617_ (.A1(_03048_),
    .A2(_03091_),
    .B(_03062_),
    .Y(_03259_));
 AND2x2_ASAP7_75t_R _25618_ (.A(_03259_),
    .B(_03067_),
    .Y(_03260_));
 AOI21x1_ASAP7_75t_SL _25619_ (.A1(_03087_),
    .A2(_03040_),
    .B(_03062_),
    .Y(_03261_));
 AO21x1_ASAP7_75t_R _25620_ (.A1(_03261_),
    .A2(_03149_),
    .B(_03080_),
    .Y(_03262_));
 AOI21x1_ASAP7_75t_R _25621_ (.A1(_03093_),
    .A2(_03113_),
    .B(_03084_),
    .Y(_03263_));
 NAND2x1_ASAP7_75t_R _25622_ (.A(_03088_),
    .B(_03176_),
    .Y(_03264_));
 AOI21x1_ASAP7_75t_R _25624_ (.A1(_03263_),
    .A2(_03264_),
    .B(_03184_),
    .Y(_03266_));
 OAI21x1_ASAP7_75t_R _25625_ (.A1(_03260_),
    .A2(_03262_),
    .B(_03266_),
    .Y(_03267_));
 OAI21x1_ASAP7_75t_R _25626_ (.A1(_03250_),
    .A2(_03258_),
    .B(_03267_),
    .Y(_03268_));
 AOI21x1_ASAP7_75t_SL _25627_ (.A1(_03068_),
    .A2(_03040_),
    .B(_03062_),
    .Y(_03269_));
 AND2x2_ASAP7_75t_R _25628_ (.A(_03269_),
    .B(_03088_),
    .Y(_03270_));
 INVx1_ASAP7_75t_R _25629_ (.A(_03170_),
    .Y(_03271_));
 AO21x1_ASAP7_75t_R _25630_ (.A1(_03040_),
    .A2(_03122_),
    .B(_03093_),
    .Y(_03272_));
 NOR2x1_ASAP7_75t_R _25631_ (.A(_03080_),
    .B(_03144_),
    .Y(_03273_));
 OAI21x1_ASAP7_75t_R _25632_ (.A1(_03271_),
    .A2(_03272_),
    .B(_03273_),
    .Y(_03274_));
 NOR2x1_ASAP7_75t_R _25633_ (.A(_03270_),
    .B(_03274_),
    .Y(_03275_));
 NOR2x1_ASAP7_75t_SL _25634_ (.A(_03043_),
    .B(_03048_),
    .Y(_03276_));
 OAI21x1_ASAP7_75t_R _25635_ (.A1(_03276_),
    .A2(_03160_),
    .B(_03144_),
    .Y(_03277_));
 OAI21x1_ASAP7_75t_R _25636_ (.A1(_03245_),
    .A2(_03194_),
    .B(_03084_),
    .Y(_03278_));
 NOR2x1_ASAP7_75t_R _25637_ (.A(_03277_),
    .B(_03278_),
    .Y(_03279_));
 NAND2x1_ASAP7_75t_R _25638_ (.A(_01262_),
    .B(_03048_),
    .Y(_03280_));
 AOI21x1_ASAP7_75t_R _25639_ (.A1(_03131_),
    .A2(_03280_),
    .B(_03093_),
    .Y(_03281_));
 INVx1_ASAP7_75t_R _25640_ (.A(_01270_),
    .Y(_03282_));
 NAND2x1_ASAP7_75t_R _25641_ (.A(_03093_),
    .B(_03144_),
    .Y(_03283_));
 OAI21x1_ASAP7_75t_R _25642_ (.A1(_03282_),
    .A2(_03283_),
    .B(_03080_),
    .Y(_03284_));
 OAI21x1_ASAP7_75t_R _25643_ (.A1(_03281_),
    .A2(_03284_),
    .B(_03103_),
    .Y(_03285_));
 NOR3x1_ASAP7_75t_SL _25644_ (.A(_03275_),
    .B(_03279_),
    .C(_03285_),
    .Y(_03286_));
 AOI21x1_ASAP7_75t_SL _25645_ (.A1(_03104_),
    .A2(_03268_),
    .B(_03286_),
    .Y(_03287_));
 NAND2x1_ASAP7_75t_SL _25646_ (.A(_03163_),
    .B(_03200_),
    .Y(_03288_));
 AOI21x1_ASAP7_75t_R _25647_ (.A1(_03093_),
    .A2(_03070_),
    .B(_03084_),
    .Y(_03289_));
 AOI21x1_ASAP7_75t_SL _25649_ (.A1(_03288_),
    .A2(_03289_),
    .B(_03144_),
    .Y(_03291_));
 AOI21x1_ASAP7_75t_R _25651_ (.A1(_03113_),
    .A2(_03064_),
    .B(_03080_),
    .Y(_03293_));
 OAI21x1_ASAP7_75t_R _25652_ (.A1(_03052_),
    .A2(_03048_),
    .B(_03062_),
    .Y(_03294_));
 AO21x1_ASAP7_75t_R _25653_ (.A1(_01258_),
    .A2(_03048_),
    .B(_03294_),
    .Y(_03295_));
 NAND2x1_ASAP7_75t_R _25654_ (.A(_03293_),
    .B(_03295_),
    .Y(_03296_));
 AOI21x1_ASAP7_75t_R _25655_ (.A1(_03291_),
    .A2(_03296_),
    .B(_03104_),
    .Y(_03297_));
 NOR2x1p5_ASAP7_75t_SL _25656_ (.A(_03066_),
    .B(_03252_),
    .Y(_03298_));
 NAND2x1_ASAP7_75t_SL _25657_ (.A(_03043_),
    .B(_03048_),
    .Y(_03299_));
 NAND2x1_ASAP7_75t_R _25659_ (.A(_01272_),
    .B(_03093_),
    .Y(_03301_));
 OA21x2_ASAP7_75t_R _25660_ (.A1(_03299_),
    .A2(_03093_),
    .B(_03301_),
    .Y(_03302_));
 AOI21x1_ASAP7_75t_R _25661_ (.A1(_03235_),
    .A2(_03302_),
    .B(_03184_),
    .Y(_03303_));
 OAI21x1_ASAP7_75t_R _25662_ (.A1(_03229_),
    .A2(_03298_),
    .B(_03303_),
    .Y(_03304_));
 NAND2x1_ASAP7_75t_SL _25663_ (.A(_03297_),
    .B(_03304_),
    .Y(_03305_));
 NOR2x1_ASAP7_75t_R _25664_ (.A(_01258_),
    .B(_03048_),
    .Y(_03306_));
 NOR2x1_ASAP7_75t_R _25665_ (.A(_03306_),
    .B(_03124_),
    .Y(_03307_));
 INVx1_ASAP7_75t_R _25666_ (.A(_03127_),
    .Y(_03308_));
 NOR2x1_ASAP7_75t_R _25667_ (.A(_03308_),
    .B(_03294_),
    .Y(_03309_));
 OAI21x1_ASAP7_75t_R _25668_ (.A1(_03307_),
    .A2(_03309_),
    .B(_03084_),
    .Y(_03310_));
 NAND2x1_ASAP7_75t_R _25669_ (.A(_03043_),
    .B(_01259_),
    .Y(_03311_));
 AOI21x1_ASAP7_75t_R _25670_ (.A1(_03311_),
    .A2(_03064_),
    .B(_03084_),
    .Y(_03312_));
 AO21x1_ASAP7_75t_R _25671_ (.A1(_03162_),
    .A2(_03251_),
    .B(_03093_),
    .Y(_03313_));
 AOI21x1_ASAP7_75t_R _25672_ (.A1(_03312_),
    .A2(_03313_),
    .B(_03184_),
    .Y(_03314_));
 NAND2x1_ASAP7_75t_SL _25673_ (.A(_03310_),
    .B(_03314_),
    .Y(_03315_));
 NAND2x1_ASAP7_75t_R _25674_ (.A(_03149_),
    .B(_03261_),
    .Y(_03316_));
 AOI21x1_ASAP7_75t_R _25675_ (.A1(_03062_),
    .A2(_03179_),
    .B(_03084_),
    .Y(_03317_));
 AOI21x1_ASAP7_75t_R _25676_ (.A1(_03316_),
    .A2(_03317_),
    .B(_03144_),
    .Y(_03318_));
 AOI21x1_ASAP7_75t_R _25677_ (.A1(_03299_),
    .A2(_03173_),
    .B(_03080_),
    .Y(_03319_));
 OAI21x1_ASAP7_75t_R _25678_ (.A1(_03093_),
    .A2(_03280_),
    .B(_03319_),
    .Y(_03320_));
 AOI21x1_ASAP7_75t_R _25679_ (.A1(_03318_),
    .A2(_03320_),
    .B(_03103_),
    .Y(_03321_));
 AOI21x1_ASAP7_75t_R _25680_ (.A1(_03315_),
    .A2(_03321_),
    .B(_03191_),
    .Y(_03322_));
 NAND2x1_ASAP7_75t_SL _25681_ (.A(_03305_),
    .B(_03322_),
    .Y(_03323_));
 OAI21x1_ASAP7_75t_SL _25682_ (.A1(_03244_),
    .A2(_03287_),
    .B(_03323_),
    .Y(_00105_));
 INVx1_ASAP7_75t_R _25683_ (.A(_03045_),
    .Y(_03324_));
 AOI21x1_ASAP7_75t_SL _25684_ (.A1(_03046_),
    .A2(_03324_),
    .B(_01263_),
    .Y(_03325_));
 OAI21x1_ASAP7_75t_R _25685_ (.A1(_03237_),
    .A2(_03325_),
    .B(_03062_),
    .Y(_03326_));
 AOI21x1_ASAP7_75t_R _25686_ (.A1(_01258_),
    .A2(_03040_),
    .B(_03062_),
    .Y(_03327_));
 NAND2x1_ASAP7_75t_R _25687_ (.A(_03170_),
    .B(_03327_),
    .Y(_03328_));
 AOI21x1_ASAP7_75t_R _25688_ (.A1(_03326_),
    .A2(_03328_),
    .B(_03080_),
    .Y(_03329_));
 NAND2x1_ASAP7_75t_R _25689_ (.A(_03299_),
    .B(_03327_),
    .Y(_03330_));
 OAI21x1_ASAP7_75t_R _25690_ (.A1(_03237_),
    .A2(_03306_),
    .B(_03062_),
    .Y(_03331_));
 AOI21x1_ASAP7_75t_R _25692_ (.A1(_03330_),
    .A2(_03331_),
    .B(_03084_),
    .Y(_03333_));
 OAI21x1_ASAP7_75t_R _25693_ (.A1(_03329_),
    .A2(_03333_),
    .B(_03144_),
    .Y(_03334_));
 OAI21x1_ASAP7_75t_R _25694_ (.A1(_03325_),
    .A2(_03160_),
    .B(_03084_),
    .Y(_03335_));
 AO21x1_ASAP7_75t_SL _25695_ (.A1(_03040_),
    .A2(_03043_),
    .B(_03062_),
    .Y(_03336_));
 NOR2x1_ASAP7_75t_SL _25696_ (.A(_03237_),
    .B(_03336_),
    .Y(_03337_));
 NOR2x1_ASAP7_75t_SL _25697_ (.A(_03335_),
    .B(_03337_),
    .Y(_03338_));
 AOI21x1_ASAP7_75t_SL _25698_ (.A1(_01261_),
    .A2(_03040_),
    .B(_03093_),
    .Y(_03339_));
 NAND2x1_ASAP7_75t_R _25699_ (.A(_03170_),
    .B(_03339_),
    .Y(_03340_));
 NAND2x1p5_ASAP7_75t_SL _25700_ (.A(_03125_),
    .B(_03199_),
    .Y(_03341_));
 AOI21x1_ASAP7_75t_SL _25701_ (.A1(_03340_),
    .A2(_03341_),
    .B(_03084_),
    .Y(_03342_));
 OAI21x1_ASAP7_75t_SL _25702_ (.A1(_03342_),
    .A2(_03338_),
    .B(_03184_),
    .Y(_03343_));
 AOI21x1_ASAP7_75t_SL _25703_ (.A1(_03343_),
    .A2(_03334_),
    .B(_03103_),
    .Y(_03344_));
 OAI21x1_ASAP7_75t_R _25704_ (.A1(_03325_),
    .A2(_03179_),
    .B(_03062_),
    .Y(_03345_));
 INVx1_ASAP7_75t_SL _25705_ (.A(_03071_),
    .Y(_03346_));
 NAND2x1_ASAP7_75t_SL _25706_ (.A(_03269_),
    .B(_03346_),
    .Y(_03347_));
 AOI21x1_ASAP7_75t_R _25707_ (.A1(_03345_),
    .A2(_03347_),
    .B(_03080_),
    .Y(_03348_));
 INVx1_ASAP7_75t_SL _25708_ (.A(_03201_),
    .Y(_03349_));
 NAND2x1_ASAP7_75t_R _25709_ (.A(_03093_),
    .B(_03212_),
    .Y(_03350_));
 OAI21x1_ASAP7_75t_R _25710_ (.A1(_03306_),
    .A2(_03350_),
    .B(_03080_),
    .Y(_03351_));
 OAI21x1_ASAP7_75t_R _25711_ (.A1(_03349_),
    .A2(_03351_),
    .B(_03144_),
    .Y(_03352_));
 NOR2x1_ASAP7_75t_SL _25712_ (.A(_03348_),
    .B(_03352_),
    .Y(_03353_));
 INVx1_ASAP7_75t_R _25713_ (.A(_03171_),
    .Y(_03354_));
 NAND2x1_ASAP7_75t_R _25714_ (.A(_03261_),
    .B(_03067_),
    .Y(_03355_));
 AOI21x1_ASAP7_75t_R _25715_ (.A1(_03354_),
    .A2(_03355_),
    .B(_03084_),
    .Y(_03356_));
 AOI21x1_ASAP7_75t_R _25716_ (.A1(_03043_),
    .A2(_03040_),
    .B(_03093_),
    .Y(_03357_));
 AND2x2_ASAP7_75t_SL _25717_ (.A(_03357_),
    .B(_03149_),
    .Y(_03358_));
 OAI21x1_ASAP7_75t_R _25718_ (.A1(_03052_),
    .A2(_03040_),
    .B(_03093_),
    .Y(_03359_));
 OAI21x1_ASAP7_75t_R _25719_ (.A1(_03220_),
    .A2(_03359_),
    .B(_03084_),
    .Y(_03360_));
 OAI21x1_ASAP7_75t_R _25720_ (.A1(_03358_),
    .A2(_03360_),
    .B(_03184_),
    .Y(_03361_));
 OAI21x1_ASAP7_75t_R _25721_ (.A1(_03356_),
    .A2(_03361_),
    .B(_03103_),
    .Y(_03362_));
 OAI21x1_ASAP7_75t_R _25722_ (.A1(_03362_),
    .A2(_03353_),
    .B(_03191_),
    .Y(_03363_));
 NOR2x1_ASAP7_75t_SL _25723_ (.A(_03363_),
    .B(_03344_),
    .Y(_03364_));
 AND2x2_ASAP7_75t_R _25724_ (.A(_01258_),
    .B(_01255_),
    .Y(_03365_));
 NAND2x1p5_ASAP7_75t_L _25725_ (.A(_03365_),
    .B(_03048_),
    .Y(_03366_));
 AOI211x1_ASAP7_75t_R _25726_ (.A1(_03261_),
    .A2(_03366_),
    .B(_03281_),
    .C(_03080_),
    .Y(_03367_));
 AO21x1_ASAP7_75t_SL _25727_ (.A1(_01258_),
    .A2(_03040_),
    .B(_03124_),
    .Y(_03368_));
 AO21x1_ASAP7_75t_R _25728_ (.A1(_03368_),
    .A2(_03129_),
    .B(_03144_),
    .Y(_03369_));
 AND2x2_ASAP7_75t_R _25729_ (.A(_03093_),
    .B(_01267_),
    .Y(_03370_));
 NOR2x1_ASAP7_75t_R _25730_ (.A(_03370_),
    .B(_03171_),
    .Y(_03371_));
 NAND2x1_ASAP7_75t_R _25731_ (.A(_03080_),
    .B(_03371_),
    .Y(_03372_));
 OA21x2_ASAP7_75t_R _25732_ (.A1(_01273_),
    .A2(_03093_),
    .B(_03084_),
    .Y(_03373_));
 AOI21x1_ASAP7_75t_R _25733_ (.A1(_03373_),
    .A2(_03347_),
    .B(_03184_),
    .Y(_03374_));
 AOI21x1_ASAP7_75t_R _25734_ (.A1(_03372_),
    .A2(_03374_),
    .B(_03104_),
    .Y(_03375_));
 OAI21x1_ASAP7_75t_SL _25735_ (.A1(_03369_),
    .A2(_03367_),
    .B(_03375_),
    .Y(_03376_));
 NAND2x1_ASAP7_75t_L _25736_ (.A(_03068_),
    .B(_03048_),
    .Y(_03377_));
 NOR2x1_ASAP7_75t_R _25737_ (.A(_01268_),
    .B(_03093_),
    .Y(_03378_));
 AOI21x1_ASAP7_75t_R _25738_ (.A1(_03377_),
    .A2(_03112_),
    .B(_03378_),
    .Y(_03379_));
 AOI21x1_ASAP7_75t_R _25739_ (.A1(_03080_),
    .A2(_03379_),
    .B(_03144_),
    .Y(_03380_));
 NOR2x1_ASAP7_75t_R _25740_ (.A(_03062_),
    .B(_03052_),
    .Y(_03381_));
 NOR2x1_ASAP7_75t_R _25741_ (.A(_03062_),
    .B(_03048_),
    .Y(_03382_));
 OAI21x1_ASAP7_75t_R _25742_ (.A1(_03381_),
    .A2(_03382_),
    .B(_03090_),
    .Y(_03383_));
 NAND3x1_ASAP7_75t_R _25743_ (.A(_03383_),
    .B(_03201_),
    .C(_03084_),
    .Y(_03384_));
 AOI21x1_ASAP7_75t_R _25744_ (.A1(_03380_),
    .A2(_03384_),
    .B(_03103_),
    .Y(_03385_));
 NAND2x1_ASAP7_75t_R _25745_ (.A(_01253_),
    .B(_03040_),
    .Y(_03386_));
 AND2x2_ASAP7_75t_R _25746_ (.A(_03200_),
    .B(_03386_),
    .Y(_03387_));
 AO21x1_ASAP7_75t_R _25747_ (.A1(_03040_),
    .A2(_03148_),
    .B(_03062_),
    .Y(_03388_));
 NOR2x1_ASAP7_75t_R _25748_ (.A(_03156_),
    .B(_03388_),
    .Y(_03389_));
 OAI21x1_ASAP7_75t_SL _25749_ (.A1(_03387_),
    .A2(_03389_),
    .B(_03084_),
    .Y(_03390_));
 NAND2x1_ASAP7_75t_R _25750_ (.A(_01270_),
    .B(_03062_),
    .Y(_03391_));
 NOR2x1_ASAP7_75t_SL _25751_ (.A(_03062_),
    .B(_03071_),
    .Y(_03392_));
 AOI21x1_ASAP7_75t_SL _25752_ (.A1(_03163_),
    .A2(_03392_),
    .B(_03084_),
    .Y(_03393_));
 AOI21x1_ASAP7_75t_R _25753_ (.A1(_03391_),
    .A2(_03393_),
    .B(_03184_),
    .Y(_03394_));
 NAND2x1_ASAP7_75t_L _25754_ (.A(_03390_),
    .B(_03394_),
    .Y(_03395_));
 NAND2x1_ASAP7_75t_R _25755_ (.A(_03385_),
    .B(_03395_),
    .Y(_03396_));
 AOI21x1_ASAP7_75t_SL _25756_ (.A1(_03376_),
    .A2(_03396_),
    .B(_03191_),
    .Y(_03397_));
 NOR2x1_ASAP7_75t_SL _25757_ (.A(_03397_),
    .B(_03364_),
    .Y(_00106_));
 NOR2x1_ASAP7_75t_L _25758_ (.A(_03308_),
    .B(_03252_),
    .Y(_03398_));
 NOR2x1_ASAP7_75t_R _25759_ (.A(_03156_),
    .B(_03294_),
    .Y(_03399_));
 OAI21x1_ASAP7_75t_R _25760_ (.A1(_03398_),
    .A2(_03399_),
    .B(_03084_),
    .Y(_03400_));
 NAND2x1_ASAP7_75t_R _25761_ (.A(_03327_),
    .B(_03067_),
    .Y(_03401_));
 AOI21x1_ASAP7_75t_R _25762_ (.A1(_03149_),
    .A2(_03357_),
    .B(_03084_),
    .Y(_03402_));
 AOI21x1_ASAP7_75t_R _25763_ (.A1(_03401_),
    .A2(_03402_),
    .B(_03144_),
    .Y(_03403_));
 NAND2x1_ASAP7_75t_R _25764_ (.A(_03400_),
    .B(_03403_),
    .Y(_03404_));
 INVx2_ASAP7_75t_R _25765_ (.A(_03113_),
    .Y(_03405_));
 OAI21x1_ASAP7_75t_SL _25766_ (.A1(_03159_),
    .A2(_03254_),
    .B(_03062_),
    .Y(_03406_));
 OAI21x1_ASAP7_75t_R _25767_ (.A1(_03405_),
    .A2(_03336_),
    .B(_03406_),
    .Y(_03407_));
 NAND2x1_ASAP7_75t_R _25768_ (.A(_03170_),
    .B(_03357_),
    .Y(_03408_));
 NOR2x1_ASAP7_75t_R _25769_ (.A(_03080_),
    .B(_03112_),
    .Y(_03409_));
 AOI21x1_ASAP7_75t_R _25770_ (.A1(_03408_),
    .A2(_03409_),
    .B(_03184_),
    .Y(_03410_));
 OAI21x1_ASAP7_75t_R _25771_ (.A1(_03084_),
    .A2(_03407_),
    .B(_03410_),
    .Y(_03411_));
 AOI21x1_ASAP7_75t_R _25772_ (.A1(_03404_),
    .A2(_03411_),
    .B(_03104_),
    .Y(_03412_));
 INVx1_ASAP7_75t_R _25773_ (.A(_03269_),
    .Y(_03413_));
 NAND3x1_ASAP7_75t_SL _25774_ (.A(_03406_),
    .B(_03080_),
    .C(_03413_),
    .Y(_03414_));
 NAND2x1_ASAP7_75t_R _25775_ (.A(_03149_),
    .B(_03339_),
    .Y(_03415_));
 AOI21x1_ASAP7_75t_SL _25776_ (.A1(_03415_),
    .A2(_03319_),
    .B(_03184_),
    .Y(_03416_));
 NAND2x1_ASAP7_75t_R _25777_ (.A(_03414_),
    .B(_03416_),
    .Y(_03417_));
 AO21x1_ASAP7_75t_SL _25778_ (.A1(_03113_),
    .A2(_03131_),
    .B(_03093_),
    .Y(_03418_));
 NOR2x1_ASAP7_75t_R _25779_ (.A(_03043_),
    .B(_01259_),
    .Y(_03419_));
 OAI21x1_ASAP7_75t_R _25780_ (.A1(_03419_),
    .A2(_03254_),
    .B(_03093_),
    .Y(_03420_));
 AOI21x1_ASAP7_75t_SL _25781_ (.A1(_03420_),
    .A2(_03418_),
    .B(_03080_),
    .Y(_03421_));
 NOR2x1_ASAP7_75t_R _25782_ (.A(_03087_),
    .B(_03040_),
    .Y(_03422_));
 NOR2x1_ASAP7_75t_R _25783_ (.A(_01254_),
    .B(_03048_),
    .Y(_03423_));
 OAI21x1_ASAP7_75t_R _25784_ (.A1(_03422_),
    .A2(_03423_),
    .B(_03062_),
    .Y(_03424_));
 OAI21x1_ASAP7_75t_R _25785_ (.A1(_03070_),
    .A2(_03156_),
    .B(_03093_),
    .Y(_03425_));
 AOI21x1_ASAP7_75t_R _25786_ (.A1(_03424_),
    .A2(_03425_),
    .B(_03084_),
    .Y(_03426_));
 OAI21x1_ASAP7_75t_SL _25787_ (.A1(_03426_),
    .A2(_03421_),
    .B(_03184_),
    .Y(_03427_));
 AOI21x1_ASAP7_75t_SL _25788_ (.A1(_03427_),
    .A2(_03417_),
    .B(_03103_),
    .Y(_03428_));
 OAI21x1_ASAP7_75t_SL _25789_ (.A1(_03428_),
    .A2(_03412_),
    .B(_03244_),
    .Y(_03429_));
 NOR2x1_ASAP7_75t_SL _25790_ (.A(_03113_),
    .B(_03093_),
    .Y(_03430_));
 OA21x2_ASAP7_75t_R _25791_ (.A1(_03430_),
    .A2(_03214_),
    .B(_03084_),
    .Y(_03431_));
 NAND2x1_ASAP7_75t_R _25792_ (.A(_03093_),
    .B(_03237_),
    .Y(_03432_));
 AOI21x1_ASAP7_75t_R _25793_ (.A1(_03432_),
    .A2(_03340_),
    .B(_03084_),
    .Y(_03433_));
 OAI21x1_ASAP7_75t_SL _25794_ (.A1(_03431_),
    .A2(_03433_),
    .B(_03184_),
    .Y(_03434_));
 NAND2x1_ASAP7_75t_R _25795_ (.A(_03366_),
    .B(_03173_),
    .Y(_03435_));
 NAND2x1p5_ASAP7_75t_SL _25796_ (.A(_03176_),
    .B(_03113_),
    .Y(_03436_));
 AOI21x1_ASAP7_75t_SL _25797_ (.A1(_03436_),
    .A2(_03435_),
    .B(_03084_),
    .Y(_03437_));
 AO21x1_ASAP7_75t_R _25798_ (.A1(_03092_),
    .A2(_03251_),
    .B(_03062_),
    .Y(_03438_));
 NOR2x1_ASAP7_75t_R _25799_ (.A(_01256_),
    .B(_03040_),
    .Y(_03439_));
 OAI21x1_ASAP7_75t_R _25800_ (.A1(_03202_),
    .A2(_03439_),
    .B(_03062_),
    .Y(_03440_));
 AOI21x1_ASAP7_75t_R _25801_ (.A1(_03438_),
    .A2(_03440_),
    .B(_03080_),
    .Y(_03441_));
 OAI21x1_ASAP7_75t_SL _25802_ (.A1(_03441_),
    .A2(_03437_),
    .B(_03144_),
    .Y(_03442_));
 AOI21x1_ASAP7_75t_SL _25803_ (.A1(_03442_),
    .A2(_03434_),
    .B(_03104_),
    .Y(_03443_));
 INVx1_ASAP7_75t_R _25804_ (.A(_03335_),
    .Y(_03444_));
 AOI21x1_ASAP7_75t_SL _25805_ (.A1(_01261_),
    .A2(_03040_),
    .B(_03062_),
    .Y(_03445_));
 NAND2x1_ASAP7_75t_SL _25806_ (.A(_03366_),
    .B(_03445_),
    .Y(_03446_));
 OAI21x1_ASAP7_75t_R _25807_ (.A1(_03202_),
    .A2(_03422_),
    .B(_03062_),
    .Y(_03447_));
 AOI21x1_ASAP7_75t_R _25808_ (.A1(_03446_),
    .A2(_03447_),
    .B(_03084_),
    .Y(_03448_));
 OAI21x1_ASAP7_75t_R _25809_ (.A1(_03444_),
    .A2(_03448_),
    .B(_03144_),
    .Y(_03449_));
 AOI21x1_ASAP7_75t_R _25810_ (.A1(_03288_),
    .A2(_03224_),
    .B(_03084_),
    .Y(_03450_));
 NOR2x1_ASAP7_75t_R _25811_ (.A(_01254_),
    .B(_03040_),
    .Y(_03451_));
 OAI21x1_ASAP7_75t_R _25812_ (.A1(_03325_),
    .A2(_03451_),
    .B(_03062_),
    .Y(_03452_));
 NOR2x1_ASAP7_75t_R _25813_ (.A(_01259_),
    .B(_03048_),
    .Y(_03453_));
 OAI21x1_ASAP7_75t_R _25814_ (.A1(_03237_),
    .A2(_03453_),
    .B(_03093_),
    .Y(_03454_));
 AOI21x1_ASAP7_75t_R _25815_ (.A1(_03452_),
    .A2(_03454_),
    .B(_03080_),
    .Y(_03455_));
 OAI21x1_ASAP7_75t_R _25816_ (.A1(_03450_),
    .A2(_03455_),
    .B(_03184_),
    .Y(_03456_));
 AOI21x1_ASAP7_75t_R _25817_ (.A1(_03449_),
    .A2(_03456_),
    .B(_03103_),
    .Y(_03457_));
 OAI21x1_ASAP7_75t_R _25818_ (.A1(_03457_),
    .A2(_03443_),
    .B(_03191_),
    .Y(_03458_));
 NAND2x1_ASAP7_75t_SL _25819_ (.A(_03458_),
    .B(_03429_),
    .Y(_00107_));
 NAND2x1_ASAP7_75t_R _25820_ (.A(_01256_),
    .B(_01259_),
    .Y(_03459_));
 AOI21x1_ASAP7_75t_R _25821_ (.A1(_03459_),
    .A2(_03299_),
    .B(_03093_),
    .Y(_03460_));
 AND2x2_ASAP7_75t_R _25822_ (.A(_03445_),
    .B(_03162_),
    .Y(_03461_));
 OAI21x1_ASAP7_75t_R _25823_ (.A1(_03460_),
    .A2(_03461_),
    .B(_03084_),
    .Y(_03462_));
 AO21x1_ASAP7_75t_R _25824_ (.A1(_03165_),
    .A2(_03197_),
    .B(_03084_),
    .Y(_03463_));
 AOI21x1_ASAP7_75t_R _25825_ (.A1(_03462_),
    .A2(_03463_),
    .B(_03104_),
    .Y(_03464_));
 OA21x2_ASAP7_75t_R _25826_ (.A1(_03245_),
    .A2(_03308_),
    .B(_03062_),
    .Y(_03465_));
 NOR2x1_ASAP7_75t_R _25827_ (.A(_03278_),
    .B(_03465_),
    .Y(_03466_));
 NAND2x1_ASAP7_75t_R _25828_ (.A(_03065_),
    .B(_03040_),
    .Y(_03467_));
 AO21x1_ASAP7_75t_R _25829_ (.A1(_03170_),
    .A2(_03467_),
    .B(_03093_),
    .Y(_03468_));
 NOR2x1_ASAP7_75t_R _25830_ (.A(_03084_),
    .B(_03382_),
    .Y(_03469_));
 AO21x1_ASAP7_75t_R _25831_ (.A1(_03468_),
    .A2(_03469_),
    .B(_03103_),
    .Y(_03470_));
 OAI21x1_ASAP7_75t_R _25832_ (.A1(_03466_),
    .A2(_03470_),
    .B(_03191_),
    .Y(_03471_));
 OAI21x1_ASAP7_75t_R _25833_ (.A1(_03464_),
    .A2(_03471_),
    .B(_03144_),
    .Y(_03472_));
 NAND2x1_ASAP7_75t_R _25834_ (.A(_03090_),
    .B(_03209_),
    .Y(_03473_));
 AND3x1_ASAP7_75t_SL _25835_ (.A(_03345_),
    .B(_03473_),
    .C(_03084_),
    .Y(_03474_));
 NOR2x1_ASAP7_75t_R _25836_ (.A(_03222_),
    .B(_03336_),
    .Y(_03475_));
 OAI21x1_ASAP7_75t_R _25837_ (.A1(_03475_),
    .A2(_03229_),
    .B(_03103_),
    .Y(_03476_));
 NOR2x1_ASAP7_75t_R _25838_ (.A(_03474_),
    .B(_03476_),
    .Y(_03477_));
 OA21x2_ASAP7_75t_R _25839_ (.A1(_03276_),
    .A2(_03160_),
    .B(_03393_),
    .Y(_03478_));
 AOI21x1_ASAP7_75t_R _25840_ (.A1(_03386_),
    .A2(_03392_),
    .B(_03460_),
    .Y(_03479_));
 OAI21x1_ASAP7_75t_R _25841_ (.A1(_03080_),
    .A2(_03479_),
    .B(_03104_),
    .Y(_03480_));
 OAI21x1_ASAP7_75t_R _25842_ (.A1(_03478_),
    .A2(_03480_),
    .B(_03244_),
    .Y(_03481_));
 NOR2x1_ASAP7_75t_R _25843_ (.A(_03477_),
    .B(_03481_),
    .Y(_03482_));
 OA21x2_ASAP7_75t_R _25844_ (.A1(_03087_),
    .A2(_03093_),
    .B(_03080_),
    .Y(_03483_));
 AOI21x1_ASAP7_75t_R _25845_ (.A1(_03388_),
    .A2(_03483_),
    .B(_03104_),
    .Y(_03484_));
 NAND2x1_ASAP7_75t_SL _25846_ (.A(_03299_),
    .B(_03445_),
    .Y(_03485_));
 NAND2x1_ASAP7_75t_R _25847_ (.A(_03485_),
    .B(_03213_),
    .Y(_03486_));
 AOI21x1_ASAP7_75t_R _25848_ (.A1(_03484_),
    .A2(_03486_),
    .B(_03244_),
    .Y(_03487_));
 AO21x1_ASAP7_75t_R _25849_ (.A1(_03048_),
    .A2(_01258_),
    .B(_03093_),
    .Y(_03488_));
 NOR2x1_ASAP7_75t_R _25850_ (.A(_03423_),
    .B(_03488_),
    .Y(_03489_));
 AO21x1_ASAP7_75t_L _25851_ (.A1(_03064_),
    .A2(_03088_),
    .B(_03084_),
    .Y(_03490_));
 INVx1_ASAP7_75t_R _25852_ (.A(_03259_),
    .Y(_03491_));
 NOR2x1_ASAP7_75t_R _25853_ (.A(_03080_),
    .B(_03261_),
    .Y(_03492_));
 AOI21x1_ASAP7_75t_R _25854_ (.A1(_03491_),
    .A2(_03492_),
    .B(_03103_),
    .Y(_03493_));
 OAI21x1_ASAP7_75t_R _25855_ (.A1(_03489_),
    .A2(_03490_),
    .B(_03493_),
    .Y(_03494_));
 AOI21x1_ASAP7_75t_R _25856_ (.A1(_03487_),
    .A2(_03494_),
    .B(_03144_),
    .Y(_03495_));
 AO21x1_ASAP7_75t_R _25857_ (.A1(_03040_),
    .A2(_01256_),
    .B(_03062_),
    .Y(_03496_));
 AOI21x1_ASAP7_75t_R _25858_ (.A1(_03272_),
    .A2(_03496_),
    .B(_03271_),
    .Y(_03497_));
 OAI21x1_ASAP7_75t_R _25859_ (.A1(_03195_),
    .A2(_03445_),
    .B(_03084_),
    .Y(_03498_));
 NAND2x1_ASAP7_75t_R _25860_ (.A(_03104_),
    .B(_03498_),
    .Y(_03499_));
 AOI21x1_ASAP7_75t_R _25861_ (.A1(_03080_),
    .A2(_03497_),
    .B(_03499_),
    .Y(_03500_));
 AOI21x1_ASAP7_75t_R _25862_ (.A1(_01263_),
    .A2(_03048_),
    .B(_03093_),
    .Y(_03501_));
 NAND2x1_ASAP7_75t_R _25863_ (.A(_03251_),
    .B(_03501_),
    .Y(_03502_));
 NAND2x1_ASAP7_75t_R _25864_ (.A(_03502_),
    .B(_03210_),
    .Y(_03503_));
 AOI21x1_ASAP7_75t_R _25865_ (.A1(_03093_),
    .A2(_03237_),
    .B(_03080_),
    .Y(_03504_));
 NAND2x1_ASAP7_75t_R _25866_ (.A(_03093_),
    .B(_03423_),
    .Y(_03505_));
 NAND3x1_ASAP7_75t_R _25867_ (.A(_03331_),
    .B(_03504_),
    .C(_03505_),
    .Y(_03506_));
 AOI21x1_ASAP7_75t_R _25868_ (.A1(_03503_),
    .A2(_03506_),
    .B(_03104_),
    .Y(_03507_));
 OAI21x1_ASAP7_75t_R _25869_ (.A1(_03500_),
    .A2(_03507_),
    .B(_03244_),
    .Y(_03508_));
 NAND2x1_ASAP7_75t_SL _25870_ (.A(_03495_),
    .B(_03508_),
    .Y(_03509_));
 OAI21x1_ASAP7_75t_SL _25871_ (.A1(_03472_),
    .A2(_03482_),
    .B(_03509_),
    .Y(_00108_));
 AOI21x1_ASAP7_75t_R _25872_ (.A1(_03093_),
    .A2(_03366_),
    .B(_03084_),
    .Y(_03510_));
 NAND2x1_ASAP7_75t_R _25873_ (.A(_03088_),
    .B(_03171_),
    .Y(_03511_));
 NAND2x1_ASAP7_75t_R _25874_ (.A(_03510_),
    .B(_03511_),
    .Y(_03512_));
 INVx1_ASAP7_75t_R _25875_ (.A(_03173_),
    .Y(_03513_));
 NAND2x1_ASAP7_75t_R _25876_ (.A(_03513_),
    .B(_03235_),
    .Y(_03514_));
 AOI21x1_ASAP7_75t_R _25877_ (.A1(_03512_),
    .A2(_03514_),
    .B(_03144_),
    .Y(_03515_));
 NOR2x1_ASAP7_75t_R _25878_ (.A(_03155_),
    .B(_03062_),
    .Y(_03516_));
 AOI21x1_ASAP7_75t_R _25879_ (.A1(_03062_),
    .A2(_03088_),
    .B(_03516_),
    .Y(_03517_));
 OAI21x1_ASAP7_75t_R _25880_ (.A1(_03084_),
    .A2(_03517_),
    .B(_03144_),
    .Y(_03518_));
 OAI21x1_ASAP7_75t_R _25881_ (.A1(_03325_),
    .A2(_03405_),
    .B(_03062_),
    .Y(_03519_));
 AO21x1_ASAP7_75t_R _25882_ (.A1(_03149_),
    .A2(_03131_),
    .B(_03062_),
    .Y(_03520_));
 AOI21x1_ASAP7_75t_R _25883_ (.A1(_03519_),
    .A2(_03520_),
    .B(_03080_),
    .Y(_03521_));
 OAI21x1_ASAP7_75t_R _25884_ (.A1(_03518_),
    .A2(_03521_),
    .B(_03103_),
    .Y(_03522_));
 OAI21x1_ASAP7_75t_R _25885_ (.A1(_03515_),
    .A2(_03522_),
    .B(_03191_),
    .Y(_03523_));
 NAND2x1_ASAP7_75t_R _25886_ (.A(_03299_),
    .B(_03339_),
    .Y(_03524_));
 NAND2x1_ASAP7_75t_R _25887_ (.A(_03113_),
    .B(_03269_),
    .Y(_03525_));
 AOI21x1_ASAP7_75t_R _25888_ (.A1(_03524_),
    .A2(_03525_),
    .B(_03080_),
    .Y(_03526_));
 AOI21x1_ASAP7_75t_R _25889_ (.A1(_03163_),
    .A2(_03247_),
    .B(_03381_),
    .Y(_03527_));
 NOR2x1_ASAP7_75t_SL _25890_ (.A(_03084_),
    .B(_03527_),
    .Y(_03528_));
 OAI21x1_ASAP7_75t_R _25891_ (.A1(_03526_),
    .A2(_03528_),
    .B(_03184_),
    .Y(_03529_));
 OA21x2_ASAP7_75t_R _25892_ (.A1(_03203_),
    .A2(_03306_),
    .B(_03062_),
    .Y(_03530_));
 OA21x2_ASAP7_75t_R _25893_ (.A1(_03131_),
    .A2(_03062_),
    .B(_03084_),
    .Y(_03531_));
 AO21x1_ASAP7_75t_R _25894_ (.A1(_03280_),
    .A2(_03467_),
    .B(_03093_),
    .Y(_03532_));
 AOI21x1_ASAP7_75t_R _25895_ (.A1(_03531_),
    .A2(_03532_),
    .B(_03184_),
    .Y(_03533_));
 OAI21x1_ASAP7_75t_SL _25896_ (.A1(_03490_),
    .A2(_03530_),
    .B(_03533_),
    .Y(_03534_));
 AOI21x1_ASAP7_75t_R _25897_ (.A1(_03529_),
    .A2(_03534_),
    .B(_03103_),
    .Y(_03535_));
 NOR2x1_ASAP7_75t_SL _25898_ (.A(_03523_),
    .B(_03535_),
    .Y(_03536_));
 INVx1_ASAP7_75t_R _25899_ (.A(_03454_),
    .Y(_03537_));
 AO21x1_ASAP7_75t_R _25900_ (.A1(_03113_),
    .A2(_03062_),
    .B(_03084_),
    .Y(_03538_));
 NOR2x1_ASAP7_75t_R _25901_ (.A(_03080_),
    .B(_03070_),
    .Y(_03539_));
 AOI21x1_ASAP7_75t_R _25902_ (.A1(_03488_),
    .A2(_03539_),
    .B(_03184_),
    .Y(_03540_));
 OAI21x1_ASAP7_75t_R _25903_ (.A1(_03537_),
    .A2(_03538_),
    .B(_03540_),
    .Y(_03541_));
 NAND2x1_ASAP7_75t_R _25904_ (.A(_03377_),
    .B(_03339_),
    .Y(_03542_));
 INVx1_ASAP7_75t_R _25905_ (.A(_03365_),
    .Y(_03543_));
 NAND2x1_ASAP7_75t_R _25906_ (.A(_03543_),
    .B(_03327_),
    .Y(_03544_));
 AOI21x1_ASAP7_75t_R _25907_ (.A1(_03542_),
    .A2(_03544_),
    .B(_03080_),
    .Y(_03545_));
 OAI21x1_ASAP7_75t_R _25908_ (.A1(_03325_),
    .A2(_03179_),
    .B(_03093_),
    .Y(_03546_));
 AOI21x1_ASAP7_75t_R _25909_ (.A1(_03546_),
    .A2(_03096_),
    .B(_03084_),
    .Y(_03547_));
 OAI21x1_ASAP7_75t_R _25910_ (.A1(_03545_),
    .A2(_03547_),
    .B(_03184_),
    .Y(_03548_));
 AOI21x1_ASAP7_75t_R _25911_ (.A1(_03541_),
    .A2(_03548_),
    .B(_03103_),
    .Y(_03549_));
 NOR2x1_ASAP7_75t_L _25912_ (.A(_03154_),
    .B(_03124_),
    .Y(_03550_));
 AO21x1_ASAP7_75t_R _25913_ (.A1(_03467_),
    .A2(_03062_),
    .B(_03084_),
    .Y(_03551_));
 OAI21x1_ASAP7_75t_R _25914_ (.A1(_03550_),
    .A2(_03551_),
    .B(_03144_),
    .Y(_03552_));
 AO21x1_ASAP7_75t_R _25915_ (.A1(_03299_),
    .A2(_03219_),
    .B(_03093_),
    .Y(_03553_));
 AOI21x1_ASAP7_75t_R _25916_ (.A1(_03505_),
    .A2(_03553_),
    .B(_03080_),
    .Y(_03554_));
 NOR2x1_ASAP7_75t_R _25917_ (.A(_03552_),
    .B(_03554_),
    .Y(_03555_));
 AO21x1_ASAP7_75t_R _25918_ (.A1(_03043_),
    .A2(_03093_),
    .B(_03084_),
    .Y(_03556_));
 OAI21x1_ASAP7_75t_R _25919_ (.A1(_03556_),
    .A2(_03460_),
    .B(_03184_),
    .Y(_03557_));
 AND3x1_ASAP7_75t_R _25920_ (.A(_03280_),
    .B(_03093_),
    .C(_03131_),
    .Y(_03558_));
 AO21x1_ASAP7_75t_R _25921_ (.A1(_03176_),
    .A2(_03459_),
    .B(_03080_),
    .Y(_03559_));
 NOR2x1_ASAP7_75t_R _25922_ (.A(_03558_),
    .B(_03559_),
    .Y(_03560_));
 OAI21x1_ASAP7_75t_SL _25923_ (.A1(_03557_),
    .A2(_03560_),
    .B(_03103_),
    .Y(_03561_));
 OAI21x1_ASAP7_75t_R _25924_ (.A1(_03555_),
    .A2(_03561_),
    .B(_03244_),
    .Y(_03562_));
 NOR2x1_ASAP7_75t_SL _25925_ (.A(_03549_),
    .B(_03562_),
    .Y(_03563_));
 NOR2x1_ASAP7_75t_SL _25926_ (.A(_03536_),
    .B(_03563_),
    .Y(_00109_));
 AOI21x1_ASAP7_75t_R _25927_ (.A1(_03301_),
    .A2(_03172_),
    .B(_03080_),
    .Y(_03564_));
 NAND2x1_ASAP7_75t_R _25928_ (.A(_03062_),
    .B(_03451_),
    .Y(_03565_));
 AOI21x1_ASAP7_75t_R _25929_ (.A1(_03565_),
    .A2(_03454_),
    .B(_03084_),
    .Y(_03566_));
 OAI21x1_ASAP7_75t_R _25930_ (.A1(_03564_),
    .A2(_03566_),
    .B(_03144_),
    .Y(_03567_));
 OAI21x1_ASAP7_75t_SL _25931_ (.A1(_03419_),
    .A2(_03203_),
    .B(_03093_),
    .Y(_03568_));
 INVx1_ASAP7_75t_R _25932_ (.A(_03254_),
    .Y(_03569_));
 NAND2x1_ASAP7_75t_R _25933_ (.A(_03501_),
    .B(_03569_),
    .Y(_03570_));
 AOI21x1_ASAP7_75t_R _25934_ (.A1(_03568_),
    .A2(_03570_),
    .B(_03080_),
    .Y(_03571_));
 OAI21x1_ASAP7_75t_R _25935_ (.A1(_03159_),
    .A2(_03254_),
    .B(_03093_),
    .Y(_03572_));
 OAI21x1_ASAP7_75t_R _25936_ (.A1(_03439_),
    .A2(_03070_),
    .B(_03062_),
    .Y(_03573_));
 AOI21x1_ASAP7_75t_R _25937_ (.A1(_03572_),
    .A2(_03573_),
    .B(_03084_),
    .Y(_03574_));
 OAI21x1_ASAP7_75t_R _25938_ (.A1(_03571_),
    .A2(_03574_),
    .B(_03184_),
    .Y(_03575_));
 NAND2x1_ASAP7_75t_SL _25939_ (.A(_03567_),
    .B(_03575_),
    .Y(_03576_));
 NOR2x1_ASAP7_75t_R _25940_ (.A(_03062_),
    .B(_03219_),
    .Y(_03577_));
 NOR2x1_ASAP7_75t_R _25941_ (.A(_03128_),
    .B(_03577_),
    .Y(_03578_));
 AOI21x1_ASAP7_75t_R _25942_ (.A1(_03504_),
    .A2(_03578_),
    .B(_03144_),
    .Y(_03579_));
 AO21x1_ASAP7_75t_SL _25943_ (.A1(_03299_),
    .A2(_03459_),
    .B(_03062_),
    .Y(_03580_));
 AO21x1_ASAP7_75t_R _25944_ (.A1(_01265_),
    .A2(_01271_),
    .B(_03093_),
    .Y(_03581_));
 AND2x2_ASAP7_75t_R _25945_ (.A(_03581_),
    .B(_03080_),
    .Y(_03582_));
 NAND2x1_ASAP7_75t_R _25946_ (.A(_03580_),
    .B(_03582_),
    .Y(_03583_));
 AOI21x1_ASAP7_75t_R _25947_ (.A1(_03579_),
    .A2(_03583_),
    .B(_03191_),
    .Y(_03584_));
 NAND2x1_ASAP7_75t_R _25948_ (.A(_03199_),
    .B(_03247_),
    .Y(_03585_));
 NAND2x1_ASAP7_75t_R _25949_ (.A(_03543_),
    .B(_03382_),
    .Y(_03586_));
 AND2x2_ASAP7_75t_R _25950_ (.A(_03504_),
    .B(_03586_),
    .Y(_03587_));
 NAND2x1_ASAP7_75t_R _25951_ (.A(_03585_),
    .B(_03587_),
    .Y(_03588_));
 NAND2x1_ASAP7_75t_R _25952_ (.A(_03339_),
    .B(_03067_),
    .Y(_03589_));
 OAI21x1_ASAP7_75t_R _25953_ (.A1(_03062_),
    .A2(_03092_),
    .B(_03080_),
    .Y(_03590_));
 AND3x1_ASAP7_75t_R _25954_ (.A(_03040_),
    .B(_01262_),
    .C(_03093_),
    .Y(_03591_));
 NOR2x1_ASAP7_75t_R _25955_ (.A(_03590_),
    .B(_03591_),
    .Y(_03592_));
 AOI21x1_ASAP7_75t_R _25956_ (.A1(_03589_),
    .A2(_03592_),
    .B(_03184_),
    .Y(_03593_));
 NAND2x1_ASAP7_75t_SL _25957_ (.A(_03588_),
    .B(_03593_),
    .Y(_03594_));
 NAND2x1_ASAP7_75t_SL _25958_ (.A(_03584_),
    .B(_03594_),
    .Y(_03595_));
 OAI21x1_ASAP7_75t_R _25959_ (.A1(_03244_),
    .A2(_03576_),
    .B(_03595_),
    .Y(_03596_));
 OAI21x1_ASAP7_75t_R _25960_ (.A1(_03093_),
    .A2(_03113_),
    .B(_03084_),
    .Y(_03597_));
 OAI21x1_ASAP7_75t_R _25961_ (.A1(_03597_),
    .A2(_03371_),
    .B(_03184_),
    .Y(_03598_));
 NAND2x1_ASAP7_75t_R _25962_ (.A(_03299_),
    .B(_03269_),
    .Y(_03599_));
 AO21x1_ASAP7_75t_R _25963_ (.A1(_03113_),
    .A2(_03219_),
    .B(_03093_),
    .Y(_03600_));
 AOI21x1_ASAP7_75t_R _25964_ (.A1(_03599_),
    .A2(_03600_),
    .B(_03084_),
    .Y(_03601_));
 OAI21x1_ASAP7_75t_R _25965_ (.A1(_03598_),
    .A2(_03601_),
    .B(_03244_),
    .Y(_03602_));
 INVx1_ASAP7_75t_R _25966_ (.A(_03377_),
    .Y(_03603_));
 NOR2x1_ASAP7_75t_R _25967_ (.A(_03080_),
    .B(_03132_),
    .Y(_03604_));
 OAI21x1_ASAP7_75t_R _25968_ (.A1(_03603_),
    .A2(_03496_),
    .B(_03604_),
    .Y(_03605_));
 OA21x2_ASAP7_75t_R _25969_ (.A1(_03040_),
    .A2(_03365_),
    .B(_03251_),
    .Y(_03606_));
 AOI21x1_ASAP7_75t_R _25970_ (.A1(_03209_),
    .A2(_03569_),
    .B(_03084_),
    .Y(_03607_));
 OAI21x1_ASAP7_75t_R _25971_ (.A1(_03093_),
    .A2(_03606_),
    .B(_03607_),
    .Y(_03608_));
 AOI21x1_ASAP7_75t_R _25972_ (.A1(_03605_),
    .A2(_03608_),
    .B(_03184_),
    .Y(_03609_));
 NOR2x1_ASAP7_75t_SL _25973_ (.A(_03602_),
    .B(_03609_),
    .Y(_03610_));
 NAND2x1_ASAP7_75t_R _25974_ (.A(_01266_),
    .B(_03093_),
    .Y(_03611_));
 AOI21x1_ASAP7_75t_R _25975_ (.A1(_03611_),
    .A2(_03524_),
    .B(_03084_),
    .Y(_03612_));
 NAND2x1_ASAP7_75t_R _25976_ (.A(_03084_),
    .B(_03294_),
    .Y(_03613_));
 NOR3x1_ASAP7_75t_R _25977_ (.A(_03405_),
    .B(_03325_),
    .C(_03062_),
    .Y(_03614_));
 OAI21x1_ASAP7_75t_R _25978_ (.A1(_03613_),
    .A2(_03614_),
    .B(_03184_),
    .Y(_03615_));
 NOR2x1_ASAP7_75t_R _25979_ (.A(_03612_),
    .B(_03615_),
    .Y(_03616_));
 NAND2x1_ASAP7_75t_R _25980_ (.A(_03144_),
    .B(_03351_),
    .Y(_03617_));
 AO21x1_ASAP7_75t_R _25981_ (.A1(_03040_),
    .A2(_03155_),
    .B(_03093_),
    .Y(_03618_));
 AOI21x1_ASAP7_75t_R _25982_ (.A1(_03618_),
    .A2(_03485_),
    .B(_03080_),
    .Y(_03619_));
 OAI21x1_ASAP7_75t_R _25983_ (.A1(_03617_),
    .A2(_03619_),
    .B(_03191_),
    .Y(_03620_));
 OAI21x1_ASAP7_75t_R _25984_ (.A1(_03616_),
    .A2(_03620_),
    .B(_03103_),
    .Y(_03621_));
 NOR2x1_ASAP7_75t_SL _25985_ (.A(_03610_),
    .B(_03621_),
    .Y(_03622_));
 AOI21x1_ASAP7_75t_SL _25986_ (.A1(_03104_),
    .A2(_03596_),
    .B(_03622_),
    .Y(_00110_));
 AO21x1_ASAP7_75t_R _25987_ (.A1(_03346_),
    .A2(_03150_),
    .B(_03093_),
    .Y(_03623_));
 NAND2x1_ASAP7_75t_SL _25988_ (.A(_03623_),
    .B(_03393_),
    .Y(_03624_));
 NAND2x1_ASAP7_75t_R _25989_ (.A(_03062_),
    .B(_03052_),
    .Y(_03625_));
 OAI21x1_ASAP7_75t_R _25990_ (.A1(_03271_),
    .A2(_03496_),
    .B(_03625_),
    .Y(_03626_));
 AOI21x1_ASAP7_75t_R _25991_ (.A1(_03084_),
    .A2(_03626_),
    .B(_03104_),
    .Y(_03627_));
 NAND2x1_ASAP7_75t_R _25992_ (.A(_03624_),
    .B(_03627_),
    .Y(_03628_));
 NOR2x1_ASAP7_75t_R _25993_ (.A(_03084_),
    .B(_03501_),
    .Y(_03629_));
 AOI21x1_ASAP7_75t_R _25994_ (.A1(_03485_),
    .A2(_03629_),
    .B(_03103_),
    .Y(_03630_));
 AOI22x1_ASAP7_75t_R _25995_ (.A1(_03223_),
    .A2(_03261_),
    .B1(_03176_),
    .B2(_03377_),
    .Y(_03631_));
 NAND2x1_ASAP7_75t_R _25996_ (.A(_03084_),
    .B(_03631_),
    .Y(_03632_));
 AOI21x1_ASAP7_75t_R _25997_ (.A1(_03630_),
    .A2(_03632_),
    .B(_03144_),
    .Y(_03633_));
 NAND2x1_ASAP7_75t_SL _25998_ (.A(_03628_),
    .B(_03633_),
    .Y(_03634_));
 AO21x1_ASAP7_75t_SL _25999_ (.A1(_03150_),
    .A2(_03113_),
    .B(_03093_),
    .Y(_03635_));
 NOR2x1_ASAP7_75t_R _26000_ (.A(_03080_),
    .B(_03209_),
    .Y(_03636_));
 NAND2x1_ASAP7_75t_R _26001_ (.A(_03635_),
    .B(_03636_),
    .Y(_03637_));
 NAND2x1_ASAP7_75t_R _26002_ (.A(_03093_),
    .B(_03422_),
    .Y(_03638_));
 NOR2x1_ASAP7_75t_L _26003_ (.A(_03084_),
    .B(_03430_),
    .Y(_03639_));
 AOI21x1_ASAP7_75t_R _26004_ (.A1(_03638_),
    .A2(_03639_),
    .B(_03104_),
    .Y(_03640_));
 AOI21x1_ASAP7_75t_SL _26005_ (.A1(_03640_),
    .A2(_03637_),
    .B(_03184_),
    .Y(_03641_));
 NAND3x1_ASAP7_75t_R _26006_ (.A(_03589_),
    .B(_03383_),
    .C(_03080_),
    .Y(_03642_));
 NOR2x1_ASAP7_75t_L _26007_ (.A(_03080_),
    .B(_03298_),
    .Y(_03643_));
 AOI21x1_ASAP7_75t_SL _26008_ (.A1(_03643_),
    .A2(_03436_),
    .B(_03103_),
    .Y(_03644_));
 NAND2x1_ASAP7_75t_SL _26009_ (.A(_03642_),
    .B(_03644_),
    .Y(_03645_));
 AOI21x1_ASAP7_75t_SL _26010_ (.A1(_03645_),
    .A2(_03641_),
    .B(_03244_),
    .Y(_03646_));
 NAND2x1_ASAP7_75t_SL _26011_ (.A(_03634_),
    .B(_03646_),
    .Y(_03647_));
 AOI21x1_ASAP7_75t_R _26012_ (.A1(_03227_),
    .A2(_03580_),
    .B(_03080_),
    .Y(_03648_));
 AO21x1_ASAP7_75t_R _26013_ (.A1(_03048_),
    .A2(_03122_),
    .B(_03084_),
    .Y(_03649_));
 NOR2x1_ASAP7_75t_R _26014_ (.A(_03062_),
    .B(_03276_),
    .Y(_03650_));
 NOR2x1_ASAP7_75t_R _26015_ (.A(_03259_),
    .B(_03650_),
    .Y(_03651_));
 OAI21x1_ASAP7_75t_SL _26016_ (.A1(_03649_),
    .A2(_03651_),
    .B(_03104_),
    .Y(_03652_));
 NOR2x1_ASAP7_75t_R _26017_ (.A(_03648_),
    .B(_03652_),
    .Y(_03653_));
 AO21x1_ASAP7_75t_R _26018_ (.A1(_01271_),
    .A2(_03093_),
    .B(_03084_),
    .Y(_03654_));
 NAND2x1_ASAP7_75t_L _26019_ (.A(_03062_),
    .B(_03251_),
    .Y(_03655_));
 NOR2x1_ASAP7_75t_R _26020_ (.A(_03237_),
    .B(_03655_),
    .Y(_03656_));
 OAI21x1_ASAP7_75t_R _26021_ (.A1(_03654_),
    .A2(_03656_),
    .B(_03103_),
    .Y(_03657_));
 OAI21x1_ASAP7_75t_SL _26022_ (.A1(_03124_),
    .A2(_03423_),
    .B(_03084_),
    .Y(_03658_));
 AOI21x1_ASAP7_75t_SL _26023_ (.A1(_03569_),
    .A2(_03200_),
    .B(_03658_),
    .Y(_03659_));
 OAI21x1_ASAP7_75t_SL _26024_ (.A1(_03659_),
    .A2(_03657_),
    .B(_03144_),
    .Y(_03660_));
 NOR2x1_ASAP7_75t_SL _26025_ (.A(_03653_),
    .B(_03660_),
    .Y(_03661_));
 OAI21x1_ASAP7_75t_R _26026_ (.A1(_03093_),
    .A2(_03090_),
    .B(_03213_),
    .Y(_03662_));
 OA21x2_ASAP7_75t_R _26027_ (.A1(_03087_),
    .A2(_03062_),
    .B(_03080_),
    .Y(_03663_));
 AOI21x1_ASAP7_75t_R _26028_ (.A1(_03221_),
    .A2(_03663_),
    .B(_03104_),
    .Y(_03664_));
 OAI21x1_ASAP7_75t_R _26029_ (.A1(_03246_),
    .A2(_03662_),
    .B(_03664_),
    .Y(_03665_));
 AOI21x1_ASAP7_75t_SL _26030_ (.A1(_03131_),
    .A2(_03113_),
    .B(_03062_),
    .Y(_03666_));
 AOI21x1_ASAP7_75t_R _26031_ (.A1(_03127_),
    .A2(_03150_),
    .B(_03093_),
    .Y(_03667_));
 NOR2x1_ASAP7_75t_L _26032_ (.A(_03667_),
    .B(_03666_),
    .Y(_03668_));
 AOI21x1_ASAP7_75t_R _26033_ (.A1(_03080_),
    .A2(_03668_),
    .B(_03103_),
    .Y(_03669_));
 OAI21x1_ASAP7_75t_R _26034_ (.A1(_01262_),
    .A2(_03048_),
    .B(_03200_),
    .Y(_03670_));
 NAND3x1_ASAP7_75t_R _26035_ (.A(_03670_),
    .B(_03446_),
    .C(_03084_),
    .Y(_03671_));
 NAND2x1_ASAP7_75t_L _26036_ (.A(_03669_),
    .B(_03671_),
    .Y(_03672_));
 AOI21x1_ASAP7_75t_R _26037_ (.A1(_03665_),
    .A2(_03672_),
    .B(_03144_),
    .Y(_03673_));
 OAI21x1_ASAP7_75t_SL _26038_ (.A1(_03673_),
    .A2(_03661_),
    .B(_03244_),
    .Y(_03674_));
 NAND2x1_ASAP7_75t_SL _26039_ (.A(_03647_),
    .B(_03674_),
    .Y(_00111_));
 NOR2x1p5_ASAP7_75t_L _26040_ (.A(_00574_),
    .B(_00474_),
    .Y(_03675_));
 XOR2x2_ASAP7_75t_SL _26041_ (.A(_14895_),
    .B(_12116_),
    .Y(_03676_));
 XOR2x2_ASAP7_75t_SL _26042_ (.A(_00694_),
    .B(_00687_),
    .Y(_03677_));
 XOR2x2_ASAP7_75t_SL _26043_ (.A(_12082_),
    .B(_03677_),
    .Y(_03678_));
 INVx2_ASAP7_75t_R _26044_ (.A(_03678_),
    .Y(_03679_));
 NAND2x1_ASAP7_75t_L _26045_ (.A(_03676_),
    .B(_03679_),
    .Y(_03680_));
 INVx2_ASAP7_75t_R _26046_ (.A(_03676_),
    .Y(_03681_));
 NAND2x1_ASAP7_75t_SL _26047_ (.A(_03681_),
    .B(_03678_),
    .Y(_03682_));
 AOI21x1_ASAP7_75t_SL _26048_ (.A1(_03682_),
    .A2(_03680_),
    .B(_10675_),
    .Y(_03683_));
 OAI21x1_ASAP7_75t_R _26049_ (.A1(_03675_),
    .A2(_03683_),
    .B(_00933_),
    .Y(_03684_));
 AND2x2_ASAP7_75t_R _26050_ (.A(_10675_),
    .B(_00474_),
    .Y(_03685_));
 XOR2x2_ASAP7_75t_SL _26051_ (.A(_03678_),
    .B(_03676_),
    .Y(_03686_));
 NOR2x1p5_ASAP7_75t_SL _26052_ (.A(_10675_),
    .B(_03686_),
    .Y(_03687_));
 INVx1_ASAP7_75t_R _26053_ (.A(_00933_),
    .Y(_03688_));
 OAI21x1_ASAP7_75t_R _26054_ (.A1(_03685_),
    .A2(_03687_),
    .B(_03688_),
    .Y(_03689_));
 NAND2x2_ASAP7_75t_SL _26055_ (.A(_03689_),
    .B(_03684_),
    .Y(_01279_));
 NOR2x1_ASAP7_75t_SL _26056_ (.A(_00574_),
    .B(_00475_),
    .Y(_03690_));
 XOR2x2_ASAP7_75t_SL _26057_ (.A(_00623_),
    .B(_00662_),
    .Y(_03691_));
 XOR2x2_ASAP7_75t_SL _26058_ (.A(_03691_),
    .B(_00591_),
    .Y(_03692_));
 NAND2x1_ASAP7_75t_R _26059_ (.A(_03677_),
    .B(_03692_),
    .Y(_03693_));
 NOR2x1_ASAP7_75t_L _26060_ (.A(_03677_),
    .B(_03692_),
    .Y(_03694_));
 INVx1_ASAP7_75t_R _26061_ (.A(_03694_),
    .Y(_03695_));
 AOI21x1_ASAP7_75t_SL _26062_ (.A1(_03695_),
    .A2(_03693_),
    .B(_10675_),
    .Y(_03696_));
 OAI21x1_ASAP7_75t_R _26063_ (.A1(_03690_),
    .A2(_03696_),
    .B(_00932_),
    .Y(_03697_));
 INVx1_ASAP7_75t_R _26064_ (.A(_03677_),
    .Y(_03698_));
 XOR2x2_ASAP7_75t_SL _26065_ (.A(_03691_),
    .B(_14914_),
    .Y(_03699_));
 NOR2x1_ASAP7_75t_R _26066_ (.A(_03698_),
    .B(_03699_),
    .Y(_03700_));
 OAI21x1_ASAP7_75t_SL _26067_ (.A1(_03700_),
    .A2(_03694_),
    .B(_00574_),
    .Y(_03701_));
 INVx1_ASAP7_75t_R _26068_ (.A(_00932_),
    .Y(_03702_));
 INVx1_ASAP7_75t_R _26069_ (.A(_03690_),
    .Y(_03703_));
 NAND3x1_ASAP7_75t_R _26070_ (.A(_03701_),
    .B(_03702_),
    .C(_03703_),
    .Y(_03704_));
 NAND2x2_ASAP7_75t_SL _26071_ (.A(_03704_),
    .B(_03697_),
    .Y(_01282_));
 NAND2x1_ASAP7_75t_R _26072_ (.A(_00476_),
    .B(_10675_),
    .Y(_03705_));
 XOR2x2_ASAP7_75t_SL _26073_ (.A(_00593_),
    .B(_00625_),
    .Y(_03706_));
 INVx2_ASAP7_75t_SL _26074_ (.A(_03706_),
    .Y(_03707_));
 INVx1_ASAP7_75t_R _26075_ (.A(_00689_),
    .Y(_03708_));
 XOR2x1_ASAP7_75t_SL _26076_ (.A(_14896_),
    .Y(_03709_),
    .B(_03708_));
 NAND2x1_ASAP7_75t_SL _26077_ (.A(_03707_),
    .B(_03709_),
    .Y(_03710_));
 NOR2x1_ASAP7_75t_R _26078_ (.A(_03708_),
    .B(_14896_),
    .Y(_03711_));
 XNOR2x2_ASAP7_75t_L _26079_ (.A(_00656_),
    .B(_00688_),
    .Y(_03712_));
 NOR2x1_ASAP7_75t_R _26080_ (.A(_00689_),
    .B(_03712_),
    .Y(_03713_));
 OAI21x1_ASAP7_75t_SL _26081_ (.A1(_03711_),
    .A2(_03713_),
    .B(_03706_),
    .Y(_03714_));
 NAND3x1_ASAP7_75t_SL _26082_ (.A(_03710_),
    .B(_00574_),
    .C(_03714_),
    .Y(_03715_));
 AOI21x1_ASAP7_75t_SL _26083_ (.A1(_03705_),
    .A2(_03715_),
    .B(_00903_),
    .Y(_03716_));
 NOR2x1_ASAP7_75t_R _26084_ (.A(_00574_),
    .B(_00476_),
    .Y(_03717_));
 AOI21x1_ASAP7_75t_SL _26085_ (.A1(_03714_),
    .A2(_03710_),
    .B(_10675_),
    .Y(_03718_));
 OAI21x1_ASAP7_75t_R _26086_ (.A1(_03717_),
    .A2(_03718_),
    .B(_00903_),
    .Y(_03719_));
 INVx2_ASAP7_75t_SL _26087_ (.A(_03719_),
    .Y(_03720_));
 NOR2x2_ASAP7_75t_SL _26088_ (.A(_03716_),
    .B(_03720_),
    .Y(_03721_));
 OAI21x1_ASAP7_75t_SL _26091_ (.A1(_03683_),
    .A2(_03675_),
    .B(_03688_),
    .Y(_03723_));
 OAI21x1_ASAP7_75t_SL _26092_ (.A1(_03687_),
    .A2(_03685_),
    .B(_00933_),
    .Y(_03724_));
 NAND2x2_ASAP7_75t_SL _26093_ (.A(_03724_),
    .B(_03723_),
    .Y(_01275_));
 AOI21x1_ASAP7_75t_SL _26094_ (.A1(_03705_),
    .A2(_03715_),
    .B(_08811_),
    .Y(_03725_));
 INVx1_ASAP7_75t_R _26095_ (.A(_03717_),
    .Y(_03726_));
 INVx1_ASAP7_75t_L _26096_ (.A(_03714_),
    .Y(_03727_));
 INVx1_ASAP7_75t_R _26097_ (.A(_03710_),
    .Y(_03728_));
 OAI21x1_ASAP7_75t_R _26098_ (.A1(_03727_),
    .A2(_03728_),
    .B(_00574_),
    .Y(_03729_));
 AOI21x1_ASAP7_75t_SL _26099_ (.A1(_03726_),
    .A2(_03729_),
    .B(_00903_),
    .Y(_03730_));
 NOR2x2_ASAP7_75t_SL _26100_ (.A(_03725_),
    .B(_03730_),
    .Y(_03731_));
 INVx1_ASAP7_75t_R _26103_ (.A(_01286_),
    .Y(_03733_));
 NOR2x1_ASAP7_75t_SL _26104_ (.A(_03733_),
    .B(_03721_),
    .Y(_03734_));
 INVx2_ASAP7_75t_SL _26105_ (.A(_03734_),
    .Y(_03735_));
 OAI21x1_ASAP7_75t_SL _26107_ (.A1(_03696_),
    .A2(_03690_),
    .B(_03702_),
    .Y(_03737_));
 NAND3x1_ASAP7_75t_L _26108_ (.A(_03701_),
    .B(_00932_),
    .C(_03703_),
    .Y(_03738_));
 NAND2x2_ASAP7_75t_SL _26109_ (.A(_03738_),
    .B(_03737_),
    .Y(_01274_));
 XNOR2x2_ASAP7_75t_R _26110_ (.A(_00690_),
    .B(_14945_),
    .Y(_03739_));
 XNOR2x2_ASAP7_75t_SL _26111_ (.A(_00689_),
    .B(_00694_),
    .Y(_03740_));
 XOR2x2_ASAP7_75t_R _26112_ (.A(_00594_),
    .B(_00626_),
    .Y(_03741_));
 XOR2x2_ASAP7_75t_SL _26113_ (.A(_03740_),
    .B(_03741_),
    .Y(_03742_));
 AOI21x1_ASAP7_75t_SL _26114_ (.A1(_03739_),
    .A2(_03742_),
    .B(_10675_),
    .Y(_03743_));
 OR2x2_ASAP7_75t_SL _26115_ (.A(_03742_),
    .B(_03739_),
    .Y(_03744_));
 AND2x2_ASAP7_75t_R _26116_ (.A(_10675_),
    .B(_00528_),
    .Y(_03745_));
 AOI21x1_ASAP7_75t_SL _26117_ (.A1(_03743_),
    .A2(_03744_),
    .B(_03745_),
    .Y(_03746_));
 XOR2x2_ASAP7_75t_SL _26118_ (.A(_03746_),
    .B(_00904_),
    .Y(_03747_));
 AOI21x1_ASAP7_75t_SL _26120_ (.A1(_03721_),
    .A2(_01274_),
    .B(_03747_),
    .Y(_03749_));
 NAND2x1_ASAP7_75t_SL _26121_ (.A(_03735_),
    .B(_03749_),
    .Y(_03750_));
 NAND2x2_ASAP7_75t_SL _26122_ (.A(_03731_),
    .B(_01275_),
    .Y(_03751_));
 INVx2_ASAP7_75t_SL _26123_ (.A(_01280_),
    .Y(_03752_));
 XNOR2x2_ASAP7_75t_SL _26124_ (.A(_00904_),
    .B(_03746_),
    .Y(_03753_));
 AOI21x1_ASAP7_75t_SL _26126_ (.A1(_03752_),
    .A2(_03721_),
    .B(_03753_),
    .Y(_03755_));
 NAND2x1_ASAP7_75t_SL _26127_ (.A(_03751_),
    .B(_03755_),
    .Y(_03756_));
 XOR2x2_ASAP7_75t_R _26128_ (.A(_00690_),
    .B(_00694_),
    .Y(_03757_));
 XOR2x2_ASAP7_75t_SL _26129_ (.A(_12192_),
    .B(_03757_),
    .Y(_03758_));
 XNOR2x2_ASAP7_75t_SL _26130_ (.A(_14966_),
    .B(_03758_),
    .Y(_03759_));
 NOR2x1_ASAP7_75t_R _26131_ (.A(_00574_),
    .B(_00527_),
    .Y(_03760_));
 AOI21x1_ASAP7_75t_SL _26132_ (.A1(_00574_),
    .A2(_03759_),
    .B(_03760_),
    .Y(_03761_));
 XOR2x2_ASAP7_75t_SL _26133_ (.A(_03761_),
    .B(_00905_),
    .Y(_03762_));
 INVx2_ASAP7_75t_SL _26134_ (.A(_03762_),
    .Y(_03763_));
 AO21x1_ASAP7_75t_SL _26137_ (.A1(_03750_),
    .A2(_03756_),
    .B(_03763_),
    .Y(_03766_));
 NOR2x1_ASAP7_75t_SL _26138_ (.A(_01278_),
    .B(_03721_),
    .Y(_03767_));
 NOR2x1_ASAP7_75t_SL _26140_ (.A(_03731_),
    .B(_01279_),
    .Y(_03769_));
 OAI21x1_ASAP7_75t_SL _26143_ (.A1(_03767_),
    .A2(_03769_),
    .B(_03747_),
    .Y(_03772_));
 INVx1_ASAP7_75t_L _26144_ (.A(_01285_),
    .Y(_03773_));
 NAND2x1_ASAP7_75t_SL _26145_ (.A(_03773_),
    .B(_03731_),
    .Y(_03774_));
 NAND2x1_ASAP7_75t_SL _26146_ (.A(_03774_),
    .B(_03749_),
    .Y(_03775_));
 AO21x1_ASAP7_75t_SL _26149_ (.A1(_03772_),
    .A2(_03775_),
    .B(_03762_),
    .Y(_03778_));
 XOR2x2_ASAP7_75t_R _26150_ (.A(_12222_),
    .B(_00692_),
    .Y(_03779_));
 XNOR2x2_ASAP7_75t_L _26151_ (.A(_12159_),
    .B(_03779_),
    .Y(_03780_));
 NOR2x1_ASAP7_75t_SL _26152_ (.A(_00574_),
    .B(_00526_),
    .Y(_03781_));
 AO21x1_ASAP7_75t_SL _26153_ (.A1(_03780_),
    .A2(_00574_),
    .B(_03781_),
    .Y(_03782_));
 INVx1_ASAP7_75t_R _26154_ (.A(_00906_),
    .Y(_03783_));
 XOR2x2_ASAP7_75t_SL _26155_ (.A(_03782_),
    .B(_03783_),
    .Y(_03784_));
 AOI21x1_ASAP7_75t_SL _26158_ (.A1(_03766_),
    .A2(_03778_),
    .B(_03784_),
    .Y(_03787_));
 NOR2x1_ASAP7_75t_SL _26159_ (.A(_03721_),
    .B(_01282_),
    .Y(_03788_));
 INVx2_ASAP7_75t_SL _26160_ (.A(_03788_),
    .Y(_03789_));
 NAND2x1_ASAP7_75t_SL _26161_ (.A(_03755_),
    .B(_03789_),
    .Y(_03790_));
 OAI21x1_ASAP7_75t_SL _26162_ (.A1(_03716_),
    .A2(_03720_),
    .B(_01277_),
    .Y(_03791_));
 AOI21x1_ASAP7_75t_SL _26164_ (.A1(_01286_),
    .A2(_03721_),
    .B(_03747_),
    .Y(_03793_));
 NAND2x1_ASAP7_75t_SL _26165_ (.A(_03791_),
    .B(_03793_),
    .Y(_03794_));
 AND3x1_ASAP7_75t_SL _26166_ (.A(_03790_),
    .B(_03762_),
    .C(_03794_),
    .Y(_03795_));
 AOI21x1_ASAP7_75t_SL _26169_ (.A1(_01281_),
    .A2(_03731_),
    .B(_03747_),
    .Y(_03798_));
 NAND2x1_ASAP7_75t_SL _26170_ (.A(_03752_),
    .B(_03721_),
    .Y(_03799_));
 AOI21x1_ASAP7_75t_R _26171_ (.A1(_03721_),
    .A2(_01274_),
    .B(_03753_),
    .Y(_03800_));
 AO21x1_ASAP7_75t_SL _26172_ (.A1(_03798_),
    .A2(_03799_),
    .B(_03800_),
    .Y(_03801_));
 OAI21x1_ASAP7_75t_SL _26173_ (.A1(_03762_),
    .A2(_03801_),
    .B(_03784_),
    .Y(_03802_));
 XOR2x2_ASAP7_75t_SL _26174_ (.A(_00692_),
    .B(_00693_),
    .Y(_03803_));
 XOR2x2_ASAP7_75t_R _26175_ (.A(_03803_),
    .B(_00660_),
    .Y(_03804_));
 XOR2x2_ASAP7_75t_R _26176_ (.A(_03804_),
    .B(_12267_),
    .Y(_03805_));
 NOR2x1_ASAP7_75t_R _26177_ (.A(_00574_),
    .B(_00525_),
    .Y(_03806_));
 AO21x1_ASAP7_75t_SL _26178_ (.A1(_03805_),
    .A2(_00574_),
    .B(_03806_),
    .Y(_03807_));
 XOR2x2_ASAP7_75t_SL _26179_ (.A(_03807_),
    .B(_00907_),
    .Y(_03808_));
 INVx1_ASAP7_75t_SL _26180_ (.A(_03808_),
    .Y(_03809_));
 OAI21x1_ASAP7_75t_SL _26182_ (.A1(_03795_),
    .A2(_03802_),
    .B(_03809_),
    .Y(_03811_));
 XOR2x2_ASAP7_75t_R _26183_ (.A(_14997_),
    .B(_12268_),
    .Y(_03812_));
 XOR2x2_ASAP7_75t_R _26184_ (.A(_03812_),
    .B(_12098_),
    .Y(_03813_));
 NOR2x1_ASAP7_75t_R _26185_ (.A(_00574_),
    .B(_00524_),
    .Y(_03814_));
 AO21x1_ASAP7_75t_SL _26186_ (.A1(_03813_),
    .A2(_00574_),
    .B(_03814_),
    .Y(_03815_));
 XOR2x2_ASAP7_75t_SL _26187_ (.A(_03815_),
    .B(_00908_),
    .Y(_03816_));
 OAI21x1_ASAP7_75t_SL _26188_ (.A1(_03787_),
    .A2(_03811_),
    .B(_03816_),
    .Y(_03817_));
 NAND2x1_ASAP7_75t_SL _26189_ (.A(_01276_),
    .B(_03721_),
    .Y(_03818_));
 INVx1_ASAP7_75t_SL _26190_ (.A(_01277_),
    .Y(_03819_));
 NAND2x2_ASAP7_75t_L _26191_ (.A(_03819_),
    .B(_03731_),
    .Y(_03820_));
 AO21x1_ASAP7_75t_SL _26193_ (.A1(_03818_),
    .A2(_03820_),
    .B(_03747_),
    .Y(_03822_));
 OAI21x1_ASAP7_75t_SL _26194_ (.A1(_03716_),
    .A2(_03720_),
    .B(_01276_),
    .Y(_03823_));
 OAI21x1_ASAP7_75t_R _26195_ (.A1(_03725_),
    .A2(_03730_),
    .B(_01283_),
    .Y(_03824_));
 AO21x1_ASAP7_75t_SL _26198_ (.A1(_03823_),
    .A2(_03824_),
    .B(_03753_),
    .Y(_03827_));
 AO21x1_ASAP7_75t_SL _26199_ (.A1(_03822_),
    .A2(_03827_),
    .B(_03762_),
    .Y(_03828_));
 OAI21x1_ASAP7_75t_SL _26200_ (.A1(_03725_),
    .A2(_03730_),
    .B(_01277_),
    .Y(_03829_));
 NAND2x1p5_ASAP7_75t_SL _26201_ (.A(_03753_),
    .B(_03829_),
    .Y(_03830_));
 NAND2x1_ASAP7_75t_SL _26202_ (.A(_03747_),
    .B(_03769_),
    .Y(_03831_));
 NAND2x1_ASAP7_75t_SL _26203_ (.A(_03830_),
    .B(_03831_),
    .Y(_03832_));
 OAI21x1_ASAP7_75t_SL _26204_ (.A1(_03791_),
    .A2(_03753_),
    .B(_03762_),
    .Y(_03833_));
 XOR2x2_ASAP7_75t_R _26205_ (.A(_03779_),
    .B(_12159_),
    .Y(_03834_));
 NOR2x1_ASAP7_75t_R _26206_ (.A(_10675_),
    .B(_03834_),
    .Y(_03835_));
 OAI21x1_ASAP7_75t_R _26207_ (.A1(_03781_),
    .A2(_03835_),
    .B(_03783_),
    .Y(_03836_));
 NAND2x1_ASAP7_75t_SL _26208_ (.A(_00574_),
    .B(_03780_),
    .Y(_03837_));
 INVx1_ASAP7_75t_R _26209_ (.A(_03781_),
    .Y(_03838_));
 NAND3x1_ASAP7_75t_R _26210_ (.A(_03837_),
    .B(_00906_),
    .C(_03838_),
    .Y(_03839_));
 NAND2x1_ASAP7_75t_SL _26211_ (.A(_03836_),
    .B(_03839_),
    .Y(_03840_));
 OA21x2_ASAP7_75t_SL _26214_ (.A1(_03832_),
    .A2(_03833_),
    .B(_03840_),
    .Y(_03843_));
 NAND2x1_ASAP7_75t_SL _26215_ (.A(_03828_),
    .B(_03843_),
    .Y(_03844_));
 INVx1_ASAP7_75t_R _26216_ (.A(_01276_),
    .Y(_03845_));
 NOR2x1_ASAP7_75t_SL _26217_ (.A(_03845_),
    .B(_03731_),
    .Y(_03846_));
 INVx1_ASAP7_75t_R _26218_ (.A(_03716_),
    .Y(_03847_));
 INVx1_ASAP7_75t_SL _26219_ (.A(_01283_),
    .Y(_03848_));
 AOI21x1_ASAP7_75t_R _26220_ (.A1(_03719_),
    .A2(_03847_),
    .B(_03848_),
    .Y(_03849_));
 OA21x2_ASAP7_75t_SL _26222_ (.A1(_03846_),
    .A2(_03849_),
    .B(_03753_),
    .Y(_03851_));
 NOR2x1_ASAP7_75t_SL _26223_ (.A(_03773_),
    .B(_03731_),
    .Y(_03852_));
 NOR2x1_ASAP7_75t_SL _26224_ (.A(_01277_),
    .B(_03721_),
    .Y(_03853_));
 OA21x2_ASAP7_75t_SL _26227_ (.A1(_03852_),
    .A2(_03853_),
    .B(_03747_),
    .Y(_03856_));
 OAI21x1_ASAP7_75t_SL _26228_ (.A1(_03851_),
    .A2(_03856_),
    .B(_03763_),
    .Y(_03857_));
 AOI21x1_ASAP7_75t_SL _26229_ (.A1(_03731_),
    .A2(_01282_),
    .B(_03753_),
    .Y(_03858_));
 NOR2x1_ASAP7_75t_SL _26230_ (.A(_01282_),
    .B(_01279_),
    .Y(_03859_));
 INVx2_ASAP7_75t_SL _26231_ (.A(_03859_),
    .Y(_03860_));
 NAND2x1_ASAP7_75t_SL _26232_ (.A(_03858_),
    .B(_03860_),
    .Y(_03861_));
 INVx1_ASAP7_75t_SL _26233_ (.A(_03861_),
    .Y(_03862_));
 NAND2x2_ASAP7_75t_SL _26234_ (.A(_03731_),
    .B(_01282_),
    .Y(_03863_));
 AOI21x1_ASAP7_75t_SL _26235_ (.A1(_03863_),
    .A2(_03860_),
    .B(_03747_),
    .Y(_03864_));
 OAI21x1_ASAP7_75t_SL _26236_ (.A1(_03862_),
    .A2(_03864_),
    .B(_03762_),
    .Y(_03865_));
 NAND3x1_ASAP7_75t_SL _26237_ (.A(_03857_),
    .B(_03865_),
    .C(_03784_),
    .Y(_03866_));
 AOI21x1_ASAP7_75t_SL _26238_ (.A1(_03844_),
    .A2(_03866_),
    .B(_03809_),
    .Y(_03867_));
 NAND2x1_ASAP7_75t_SL _26240_ (.A(_03747_),
    .B(_03767_),
    .Y(_03869_));
 NAND2x1_ASAP7_75t_R _26242_ (.A(_01284_),
    .B(_03721_),
    .Y(_03871_));
 AOI21x1_ASAP7_75t_SL _26243_ (.A1(_03752_),
    .A2(_03731_),
    .B(_03747_),
    .Y(_03872_));
 AOI21x1_ASAP7_75t_SL _26244_ (.A1(_03871_),
    .A2(_03872_),
    .B(_03762_),
    .Y(_03873_));
 NAND2x1_ASAP7_75t_SL _26245_ (.A(_03869_),
    .B(_03873_),
    .Y(_03874_));
 OAI21x1_ASAP7_75t_SL _26246_ (.A1(_03716_),
    .A2(_03720_),
    .B(_01280_),
    .Y(_03875_));
 AO21x1_ASAP7_75t_SL _26248_ (.A1(_03875_),
    .A2(_03824_),
    .B(_03753_),
    .Y(_03877_));
 INVx1_ASAP7_75t_R _26249_ (.A(_01278_),
    .Y(_03878_));
 NAND2x1_ASAP7_75t_SL _26250_ (.A(_03878_),
    .B(_03731_),
    .Y(_03879_));
 OA21x2_ASAP7_75t_SL _26251_ (.A1(_03879_),
    .A2(_03747_),
    .B(_03762_),
    .Y(_03880_));
 AOI21x1_ASAP7_75t_SL _26253_ (.A1(_03877_),
    .A2(_03880_),
    .B(_03840_),
    .Y(_03882_));
 NAND2x1_ASAP7_75t_SL _26254_ (.A(_03874_),
    .B(_03882_),
    .Y(_03883_));
 INVx1_ASAP7_75t_SL _26255_ (.A(_03875_),
    .Y(_03884_));
 AND2x2_ASAP7_75t_R _26256_ (.A(_01278_),
    .B(_01281_),
    .Y(_03885_));
 NOR2x1_ASAP7_75t_SL _26257_ (.A(_03885_),
    .B(_03731_),
    .Y(_03886_));
 OAI21x1_ASAP7_75t_SL _26258_ (.A1(_03884_),
    .A2(_03886_),
    .B(_03747_),
    .Y(_03887_));
 OAI21x1_ASAP7_75t_R _26259_ (.A1(_03747_),
    .A2(_03823_),
    .B(_03763_),
    .Y(_03888_));
 NAND2x1_ASAP7_75t_SL _26260_ (.A(_03753_),
    .B(_03721_),
    .Y(_03889_));
 NOR2x1_ASAP7_75t_R _26261_ (.A(_01274_),
    .B(_03889_),
    .Y(_03890_));
 NOR2x1_ASAP7_75t_SL _26262_ (.A(_03888_),
    .B(_03890_),
    .Y(_03891_));
 NAND2x1_ASAP7_75t_SL _26263_ (.A(_03887_),
    .B(_03891_),
    .Y(_03892_));
 OAI21x1_ASAP7_75t_SL _26265_ (.A1(_03725_),
    .A2(_03730_),
    .B(_03819_),
    .Y(_03894_));
 AND2x2_ASAP7_75t_R _26266_ (.A(_03753_),
    .B(_01291_),
    .Y(_03895_));
 AO21x1_ASAP7_75t_SL _26267_ (.A1(_03894_),
    .A2(_03747_),
    .B(_03895_),
    .Y(_03896_));
 AOI21x1_ASAP7_75t_SL _26269_ (.A1(_03762_),
    .A2(_03896_),
    .B(_03784_),
    .Y(_03898_));
 AOI21x1_ASAP7_75t_SL _26270_ (.A1(_03898_),
    .A2(_03892_),
    .B(_03809_),
    .Y(_03899_));
 NAND2x1_ASAP7_75t_SL _26271_ (.A(_03899_),
    .B(_03883_),
    .Y(_03900_));
 AOI21x1_ASAP7_75t_SL _26272_ (.A1(_03731_),
    .A2(_01279_),
    .B(_03753_),
    .Y(_03901_));
 NAND2x1_ASAP7_75t_SL _26273_ (.A(_03901_),
    .B(_03894_),
    .Y(_03902_));
 NAND2x1_ASAP7_75t_R _26274_ (.A(_03848_),
    .B(_03721_),
    .Y(_03903_));
 AOI21x1_ASAP7_75t_R _26275_ (.A1(_03731_),
    .A2(_01274_),
    .B(_03747_),
    .Y(_03904_));
 AOI21x1_ASAP7_75t_SL _26277_ (.A1(_03903_),
    .A2(_03904_),
    .B(_03762_),
    .Y(_03906_));
 NAND2x1_ASAP7_75t_SL _26278_ (.A(_03902_),
    .B(_03906_),
    .Y(_03907_));
 NOR2x1_ASAP7_75t_SL _26279_ (.A(_03763_),
    .B(_03798_),
    .Y(_03908_));
 OAI21x1_ASAP7_75t_R _26280_ (.A1(_03767_),
    .A2(_03846_),
    .B(_03747_),
    .Y(_03909_));
 AOI21x1_ASAP7_75t_SL _26281_ (.A1(_03908_),
    .A2(_03909_),
    .B(_03840_),
    .Y(_03910_));
 AOI21x1_ASAP7_75t_SL _26283_ (.A1(_03907_),
    .A2(_03910_),
    .B(_03808_),
    .Y(_03912_));
 INVx1_ASAP7_75t_SL _26284_ (.A(_01281_),
    .Y(_03913_));
 OAI21x1_ASAP7_75t_SL _26285_ (.A1(_03725_),
    .A2(_03730_),
    .B(_03913_),
    .Y(_03914_));
 AOI21x1_ASAP7_75t_R _26287_ (.A1(_03774_),
    .A2(_03749_),
    .B(_03762_),
    .Y(_03916_));
 OAI21x1_ASAP7_75t_SL _26288_ (.A1(_03753_),
    .A2(_03914_),
    .B(_03916_),
    .Y(_03917_));
 OA21x2_ASAP7_75t_SL _26289_ (.A1(_03914_),
    .A2(_03753_),
    .B(_03762_),
    .Y(_03918_));
 AND2x4_ASAP7_75t_SL _26290_ (.A(_03753_),
    .B(_03791_),
    .Y(_03919_));
 INVx1_ASAP7_75t_R _26292_ (.A(_01284_),
    .Y(_03921_));
 NAND2x1_ASAP7_75t_SL _26293_ (.A(_03921_),
    .B(_03731_),
    .Y(_03922_));
 NOR2x1_ASAP7_75t_R _26294_ (.A(_03753_),
    .B(_03922_),
    .Y(_03923_));
 NOR2x1_ASAP7_75t_SL _26295_ (.A(_03919_),
    .B(_03923_),
    .Y(_03924_));
 AOI21x1_ASAP7_75t_SL _26296_ (.A1(_03918_),
    .A2(_03924_),
    .B(_03784_),
    .Y(_03925_));
 NAND2x1_ASAP7_75t_SL _26297_ (.A(_03917_),
    .B(_03925_),
    .Y(_03926_));
 AOI21x1_ASAP7_75t_SL _26298_ (.A1(_03926_),
    .A2(_03912_),
    .B(_03816_),
    .Y(_03927_));
 NAND2x1_ASAP7_75t_SL _26299_ (.A(_03927_),
    .B(_03900_),
    .Y(_03928_));
 OAI21x1_ASAP7_75t_SL _26300_ (.A1(_03817_),
    .A2(_03867_),
    .B(_03928_),
    .Y(_00112_));
 INVx1_ASAP7_75t_SL _26301_ (.A(_03816_),
    .Y(_03929_));
 OA21x2_ASAP7_75t_SL _26302_ (.A1(_03788_),
    .A2(_03846_),
    .B(_03747_),
    .Y(_03930_));
 NAND2x1_ASAP7_75t_SL _26303_ (.A(_03721_),
    .B(_01275_),
    .Y(_03931_));
 AO21x1_ASAP7_75t_SL _26305_ (.A1(_03798_),
    .A2(_03931_),
    .B(_03762_),
    .Y(_03933_));
 OAI21x1_ASAP7_75t_SL _26306_ (.A1(_03930_),
    .A2(_03933_),
    .B(_03784_),
    .Y(_03934_));
 NOR2x1_ASAP7_75t_SL _26307_ (.A(_03731_),
    .B(_01274_),
    .Y(_03935_));
 AO21x1_ASAP7_75t_SL _26309_ (.A1(_03935_),
    .A2(_03747_),
    .B(_03763_),
    .Y(_03937_));
 INVx1_ASAP7_75t_R _26311_ (.A(_03823_),
    .Y(_03939_));
 NAND2x1_ASAP7_75t_SL _26312_ (.A(_03753_),
    .B(_03939_),
    .Y(_03940_));
 NAND2x1_ASAP7_75t_SL _26313_ (.A(_03940_),
    .B(_03869_),
    .Y(_03941_));
 NOR2x1p5_ASAP7_75t_SL _26314_ (.A(_03894_),
    .B(_03747_),
    .Y(_03942_));
 NOR3x1_ASAP7_75t_SL _26315_ (.A(_03937_),
    .B(_03941_),
    .C(_03942_),
    .Y(_03943_));
 AOI21x1_ASAP7_75t_SL _26316_ (.A1(_03753_),
    .A2(_03791_),
    .B(_03762_),
    .Y(_03944_));
 NAND2x1_ASAP7_75t_SL _26317_ (.A(_03774_),
    .B(_03800_),
    .Y(_03945_));
 AOI21x1_ASAP7_75t_SL _26318_ (.A1(_03944_),
    .A2(_03945_),
    .B(_03784_),
    .Y(_03946_));
 AOI21x1_ASAP7_75t_SL _26319_ (.A1(_03773_),
    .A2(_03721_),
    .B(_03747_),
    .Y(_03947_));
 AOI21x1_ASAP7_75t_SL _26320_ (.A1(_03820_),
    .A2(_03947_),
    .B(_03763_),
    .Y(_03948_));
 OA21x2_ASAP7_75t_SL _26321_ (.A1(_03731_),
    .A2(_03878_),
    .B(_03747_),
    .Y(_03949_));
 NAND2x1_ASAP7_75t_SL _26322_ (.A(_03735_),
    .B(_03949_),
    .Y(_03950_));
 NAND2x1_ASAP7_75t_SL _26323_ (.A(_03948_),
    .B(_03950_),
    .Y(_03951_));
 NAND2x1_ASAP7_75t_SL _26324_ (.A(_03946_),
    .B(_03951_),
    .Y(_03952_));
 OAI21x1_ASAP7_75t_SL _26325_ (.A1(_03934_),
    .A2(_03943_),
    .B(_03952_),
    .Y(_03953_));
 AOI21x1_ASAP7_75t_SL _26326_ (.A1(_03752_),
    .A2(_03721_),
    .B(_03747_),
    .Y(_03954_));
 AND2x2_ASAP7_75t_SL _26327_ (.A(_03954_),
    .B(_03774_),
    .Y(_03955_));
 AOI21x1_ASAP7_75t_SL _26328_ (.A1(_03845_),
    .A2(_03721_),
    .B(_03753_),
    .Y(_03956_));
 NAND2x1_ASAP7_75t_SL _26329_ (.A(_03762_),
    .B(_03784_),
    .Y(_03957_));
 AO21x1_ASAP7_75t_SL _26330_ (.A1(_03789_),
    .A2(_03956_),
    .B(_03957_),
    .Y(_03958_));
 NOR2x1_ASAP7_75t_SL _26331_ (.A(_03955_),
    .B(_03958_),
    .Y(_03959_));
 NOR2x1_ASAP7_75t_SL _26332_ (.A(_03731_),
    .B(_01275_),
    .Y(_03960_));
 OAI21x1_ASAP7_75t_R _26333_ (.A1(_03721_),
    .A2(_01274_),
    .B(_03747_),
    .Y(_03961_));
 NOR2x1_ASAP7_75t_SL _26334_ (.A(_03960_),
    .B(_03961_),
    .Y(_03962_));
 NAND2x1_ASAP7_75t_SL _26335_ (.A(_03762_),
    .B(_03840_),
    .Y(_03963_));
 AO21x1_ASAP7_75t_SL _26336_ (.A1(_03798_),
    .A2(_03931_),
    .B(_03963_),
    .Y(_03964_));
 NOR2x1_ASAP7_75t_SL _26337_ (.A(_03962_),
    .B(_03964_),
    .Y(_03965_));
 OAI21x1_ASAP7_75t_R _26338_ (.A1(_03716_),
    .A2(_03720_),
    .B(_01285_),
    .Y(_03966_));
 AOI21x1_ASAP7_75t_R _26339_ (.A1(_03824_),
    .A2(_03966_),
    .B(_03753_),
    .Y(_03967_));
 INVx1_ASAP7_75t_SL _26340_ (.A(_01293_),
    .Y(_03968_));
 NAND2x1_ASAP7_75t_SL _26341_ (.A(_03753_),
    .B(_03840_),
    .Y(_03969_));
 OAI21x1_ASAP7_75t_SL _26343_ (.A1(_03968_),
    .A2(_03969_),
    .B(_03763_),
    .Y(_03971_));
 OAI21x1_ASAP7_75t_SL _26344_ (.A1(_03967_),
    .A2(_03971_),
    .B(_03808_),
    .Y(_03972_));
 NOR3x1_ASAP7_75t_SL _26345_ (.A(_03959_),
    .B(_03965_),
    .C(_03972_),
    .Y(_03973_));
 AOI21x1_ASAP7_75t_SL _26346_ (.A1(_03809_),
    .A2(_03953_),
    .B(_03973_),
    .Y(_03974_));
 INVx1_ASAP7_75t_SL _26347_ (.A(_03830_),
    .Y(_03975_));
 NAND2x1_ASAP7_75t_SL _26348_ (.A(_03735_),
    .B(_03975_),
    .Y(_03976_));
 NAND2x1_ASAP7_75t_SL _26349_ (.A(_03914_),
    .B(_03875_),
    .Y(_03977_));
 AOI21x1_ASAP7_75t_SL _26350_ (.A1(_03747_),
    .A2(_03977_),
    .B(_03762_),
    .Y(_03978_));
 NAND2x1_ASAP7_75t_SL _26351_ (.A(_03976_),
    .B(_03978_),
    .Y(_03979_));
 INVx1_ASAP7_75t_SL _26352_ (.A(_03751_),
    .Y(_03980_));
 AND2x2_ASAP7_75t_SL _26353_ (.A(_03753_),
    .B(_01295_),
    .Y(_03981_));
 AOI21x1_ASAP7_75t_SL _26354_ (.A1(_03747_),
    .A2(_03980_),
    .B(_03981_),
    .Y(_03982_));
 AOI21x1_ASAP7_75t_SL _26355_ (.A1(_03918_),
    .A2(_03982_),
    .B(_03784_),
    .Y(_03983_));
 NAND2x1_ASAP7_75t_SL _26356_ (.A(_03979_),
    .B(_03983_),
    .Y(_03984_));
 NAND2x1_ASAP7_75t_SL _26357_ (.A(_01281_),
    .B(_03731_),
    .Y(_03985_));
 OAI21x1_ASAP7_75t_SL _26358_ (.A1(_03731_),
    .A2(_01274_),
    .B(_03747_),
    .Y(_03986_));
 INVx1_ASAP7_75t_SL _26359_ (.A(_03986_),
    .Y(_03987_));
 NAND2x1_ASAP7_75t_SL _26360_ (.A(_03985_),
    .B(_03987_),
    .Y(_03988_));
 AOI21x1_ASAP7_75t_SL _26361_ (.A1(_03791_),
    .A2(_03749_),
    .B(_03763_),
    .Y(_03989_));
 NAND2x1_ASAP7_75t_SL _26362_ (.A(_03988_),
    .B(_03989_),
    .Y(_03990_));
 OA21x2_ASAP7_75t_R _26363_ (.A1(_03730_),
    .A2(_03725_),
    .B(_01280_),
    .Y(_03991_));
 AOI21x1_ASAP7_75t_SL _26364_ (.A1(_03753_),
    .A2(_03991_),
    .B(_03762_),
    .Y(_03992_));
 NAND2x1_ASAP7_75t_SL _26365_ (.A(_03901_),
    .B(_03860_),
    .Y(_03993_));
 AOI21x1_ASAP7_75t_SL _26366_ (.A1(_03992_),
    .A2(_03993_),
    .B(_03840_),
    .Y(_03994_));
 AOI21x1_ASAP7_75t_SL _26367_ (.A1(_03990_),
    .A2(_03994_),
    .B(_03809_),
    .Y(_03995_));
 AOI21x1_ASAP7_75t_SL _26368_ (.A1(_03984_),
    .A2(_03995_),
    .B(_03816_),
    .Y(_03996_));
 NOR2x1_ASAP7_75t_SL _26369_ (.A(_01274_),
    .B(_01275_),
    .Y(_03997_));
 OAI21x1_ASAP7_75t_SL _26370_ (.A1(_03788_),
    .A2(_03997_),
    .B(_03753_),
    .Y(_03998_));
 AO21x1_ASAP7_75t_SL _26371_ (.A1(_03863_),
    .A2(_03829_),
    .B(_03753_),
    .Y(_03999_));
 AOI21x1_ASAP7_75t_SL _26372_ (.A1(_03998_),
    .A2(_03999_),
    .B(_03762_),
    .Y(_04000_));
 OAI21x1_ASAP7_75t_SL _26373_ (.A1(_03939_),
    .A2(_03986_),
    .B(_03762_),
    .Y(_04001_));
 AOI21x1_ASAP7_75t_SL _26374_ (.A1(_03919_),
    .A2(_03914_),
    .B(_04001_),
    .Y(_04002_));
 NOR2x1_ASAP7_75t_SL _26375_ (.A(_04000_),
    .B(_04002_),
    .Y(_04003_));
 NAND2x1_ASAP7_75t_SL _26376_ (.A(_03820_),
    .B(_03947_),
    .Y(_04004_));
 NOR2x1_ASAP7_75t_SL _26377_ (.A(_01281_),
    .B(_03721_),
    .Y(_04005_));
 AOI21x1_ASAP7_75t_SL _26378_ (.A1(_03747_),
    .A2(_04005_),
    .B(_03762_),
    .Y(_04006_));
 AOI21x1_ASAP7_75t_SL _26379_ (.A1(_04004_),
    .A2(_04006_),
    .B(_03840_),
    .Y(_04007_));
 AOI21x1_ASAP7_75t_SL _26380_ (.A1(_03751_),
    .A2(_03793_),
    .B(_03763_),
    .Y(_04008_));
 OAI21x1_ASAP7_75t_SL _26381_ (.A1(_03753_),
    .A2(_03966_),
    .B(_04008_),
    .Y(_04009_));
 AOI21x1_ASAP7_75t_SL _26382_ (.A1(_04007_),
    .A2(_04009_),
    .B(_03808_),
    .Y(_04010_));
 OAI21x1_ASAP7_75t_SL _26383_ (.A1(_03784_),
    .A2(_04003_),
    .B(_04010_),
    .Y(_04011_));
 NAND2x1_ASAP7_75t_SL _26384_ (.A(_03996_),
    .B(_04011_),
    .Y(_04012_));
 OAI21x1_ASAP7_75t_SL _26385_ (.A1(_03929_),
    .A2(_03974_),
    .B(_04012_),
    .Y(_00113_));
 AO21x1_ASAP7_75t_SL _26386_ (.A1(_03721_),
    .A2(_01281_),
    .B(_03747_),
    .Y(_04013_));
 NOR2x1_ASAP7_75t_SL _26387_ (.A(_03980_),
    .B(_04013_),
    .Y(_04014_));
 NOR2x1_ASAP7_75t_SL _26388_ (.A(_01284_),
    .B(_03721_),
    .Y(_04015_));
 INVx2_ASAP7_75t_SL _26389_ (.A(_03914_),
    .Y(_04016_));
 OA21x2_ASAP7_75t_SL _26390_ (.A1(_04015_),
    .A2(_04016_),
    .B(_03747_),
    .Y(_04017_));
 OAI21x1_ASAP7_75t_SL _26391_ (.A1(_04014_),
    .A2(_04017_),
    .B(_03763_),
    .Y(_04018_));
 NOR2x1_ASAP7_75t_SL _26392_ (.A(_03788_),
    .B(_04013_),
    .Y(_04019_));
 NOR2x2_ASAP7_75t_SL _26393_ (.A(_01286_),
    .B(_03731_),
    .Y(_04020_));
 OA21x2_ASAP7_75t_SL _26394_ (.A1(_04020_),
    .A2(_04015_),
    .B(_03747_),
    .Y(_04021_));
 OAI21x1_ASAP7_75t_SL _26395_ (.A1(_04019_),
    .A2(_04021_),
    .B(_03762_),
    .Y(_04022_));
 AOI21x1_ASAP7_75t_SL _26396_ (.A1(_04018_),
    .A2(_04022_),
    .B(_03784_),
    .Y(_04023_));
 OAI21x1_ASAP7_75t_R _26397_ (.A1(_03921_),
    .A2(_03731_),
    .B(_03747_),
    .Y(_04024_));
 NOR2x1_ASAP7_75t_R _26398_ (.A(_03788_),
    .B(_04024_),
    .Y(_04025_));
 AND3x1_ASAP7_75t_SL _26399_ (.A(_03791_),
    .B(_03894_),
    .C(_03753_),
    .Y(_04026_));
 OAI21x1_ASAP7_75t_SL _26400_ (.A1(_04025_),
    .A2(_04026_),
    .B(_03763_),
    .Y(_04027_));
 AO21x1_ASAP7_75t_SL _26401_ (.A1(_01275_),
    .A2(_03721_),
    .B(_03747_),
    .Y(_04028_));
 INVx1_ASAP7_75t_SL _26402_ (.A(_04020_),
    .Y(_04029_));
 AOI21x1_ASAP7_75t_SL _26403_ (.A1(_04029_),
    .A2(_03858_),
    .B(_03763_),
    .Y(_04030_));
 OAI21x1_ASAP7_75t_SL _26404_ (.A1(_04015_),
    .A2(_04028_),
    .B(_04030_),
    .Y(_04031_));
 AOI21x1_ASAP7_75t_SL _26405_ (.A1(_04027_),
    .A2(_04031_),
    .B(_03840_),
    .Y(_04032_));
 NOR3x1_ASAP7_75t_SL _26406_ (.A(_04023_),
    .B(_04032_),
    .C(_03929_),
    .Y(_04033_));
 NAND2x1_ASAP7_75t_SL _26407_ (.A(_03894_),
    .B(_03753_),
    .Y(_04034_));
 NAND2x1_ASAP7_75t_SL _26408_ (.A(_03818_),
    .B(_03901_),
    .Y(_04035_));
 OA21x2_ASAP7_75t_SL _26409_ (.A1(_03849_),
    .A2(_04034_),
    .B(_04035_),
    .Y(_04036_));
 NAND2x1_ASAP7_75t_SL _26410_ (.A(_01293_),
    .B(_03747_),
    .Y(_04037_));
 AOI21x1_ASAP7_75t_R _26411_ (.A1(_03731_),
    .A2(_01279_),
    .B(_03747_),
    .Y(_04038_));
 AOI21x1_ASAP7_75t_SL _26412_ (.A1(_04038_),
    .A2(_03860_),
    .B(_03762_),
    .Y(_04039_));
 AOI21x1_ASAP7_75t_SL _26413_ (.A1(_04037_),
    .A2(_04039_),
    .B(_03784_),
    .Y(_04040_));
 OA21x2_ASAP7_75t_SL _26414_ (.A1(_04036_),
    .A2(_03763_),
    .B(_04040_),
    .Y(_04041_));
 INVx2_ASAP7_75t_SL _26415_ (.A(_03902_),
    .Y(_04042_));
 NAND2x1_ASAP7_75t_SL _26416_ (.A(_03721_),
    .B(_01279_),
    .Y(_04043_));
 AOI21x1_ASAP7_75t_SL _26417_ (.A1(_03863_),
    .A2(_04043_),
    .B(_03747_),
    .Y(_04044_));
 NOR3x1_ASAP7_75t_SL _26418_ (.A(_04042_),
    .B(_03763_),
    .C(_04044_),
    .Y(_04045_));
 NAND2x1_ASAP7_75t_SL _26419_ (.A(_03752_),
    .B(_03731_),
    .Y(_04046_));
 NOR2x1_ASAP7_75t_SL _26420_ (.A(_01291_),
    .B(_03753_),
    .Y(_04047_));
 AO21x1_ASAP7_75t_SL _26421_ (.A1(_03975_),
    .A2(_04046_),
    .B(_04047_),
    .Y(_04048_));
 OAI21x1_ASAP7_75t_SL _26422_ (.A1(_03762_),
    .A2(_04048_),
    .B(_03784_),
    .Y(_04049_));
 OAI21x1_ASAP7_75t_SL _26423_ (.A1(_04045_),
    .A2(_04049_),
    .B(_03929_),
    .Y(_04050_));
 OAI21x1_ASAP7_75t_SL _26424_ (.A1(_04050_),
    .A2(_04041_),
    .B(_03809_),
    .Y(_04051_));
 NAND2x1_ASAP7_75t_SL _26425_ (.A(_03885_),
    .B(_03731_),
    .Y(_04052_));
 AO21x1_ASAP7_75t_SL _26426_ (.A1(_03947_),
    .A2(_04052_),
    .B(_03967_),
    .Y(_04053_));
 OAI21x1_ASAP7_75t_SL _26427_ (.A1(_04016_),
    .A2(_03853_),
    .B(_03753_),
    .Y(_04054_));
 OA21x2_ASAP7_75t_SL _26428_ (.A1(_03823_),
    .A2(_03753_),
    .B(_03763_),
    .Y(_04055_));
 AOI21x1_ASAP7_75t_SL _26429_ (.A1(_04054_),
    .A2(_04055_),
    .B(_03840_),
    .Y(_04056_));
 OAI21x1_ASAP7_75t_SL _26430_ (.A1(_03763_),
    .A2(_04053_),
    .B(_04056_),
    .Y(_04057_));
 OA21x2_ASAP7_75t_SL _26431_ (.A1(_01296_),
    .A2(_03753_),
    .B(_03762_),
    .Y(_04058_));
 NAND2x1_ASAP7_75t_SL _26432_ (.A(_03731_),
    .B(_01279_),
    .Y(_04059_));
 NAND2x1_ASAP7_75t_SL _26433_ (.A(_04059_),
    .B(_03954_),
    .Y(_04060_));
 AOI21x1_ASAP7_75t_SL _26434_ (.A1(_04058_),
    .A2(_04060_),
    .B(_03784_),
    .Y(_04061_));
 AOI21x1_ASAP7_75t_SL _26435_ (.A1(_01290_),
    .A2(_03753_),
    .B(_03755_),
    .Y(_04062_));
 NAND2x1_ASAP7_75t_SL _26436_ (.A(_03763_),
    .B(_04062_),
    .Y(_04063_));
 AOI21x1_ASAP7_75t_SL _26437_ (.A1(_04061_),
    .A2(_04063_),
    .B(_03816_),
    .Y(_04064_));
 AOI21x1_ASAP7_75t_SL _26438_ (.A1(_04057_),
    .A2(_04064_),
    .B(_03809_),
    .Y(_04065_));
 OAI21x1_ASAP7_75t_SL _26439_ (.A1(_04005_),
    .A2(_04020_),
    .B(_03747_),
    .Y(_04066_));
 AOI21x1_ASAP7_75t_SL _26440_ (.A1(_04060_),
    .A2(_04066_),
    .B(_03763_),
    .Y(_04067_));
 OAI21x1_ASAP7_75t_SL _26441_ (.A1(_03747_),
    .A2(_03977_),
    .B(_03763_),
    .Y(_04068_));
 OAI21x1_ASAP7_75t_SL _26442_ (.A1(_04042_),
    .A2(_04068_),
    .B(_03840_),
    .Y(_04069_));
 NOR2x1_ASAP7_75t_SL _26443_ (.A(_04067_),
    .B(_04069_),
    .Y(_04070_));
 INVx1_ASAP7_75t_SL _26444_ (.A(_03947_),
    .Y(_04071_));
 NOR2x1_ASAP7_75t_SL _26445_ (.A(_03762_),
    .B(_03755_),
    .Y(_04072_));
 OAI21x1_ASAP7_75t_SL _26446_ (.A1(_03734_),
    .A2(_04071_),
    .B(_04072_),
    .Y(_04073_));
 NOR2x1_ASAP7_75t_SL _26447_ (.A(_01278_),
    .B(_03731_),
    .Y(_04074_));
 OAI21x1_ASAP7_75t_SL _26448_ (.A1(_03721_),
    .A2(_01274_),
    .B(_03753_),
    .Y(_04075_));
 NOR2x1_ASAP7_75t_SL _26449_ (.A(_04074_),
    .B(_04075_),
    .Y(_04076_));
 AOI21x1_ASAP7_75t_SL _26450_ (.A1(_03791_),
    .A2(_04043_),
    .B(_03753_),
    .Y(_04077_));
 OAI21x1_ASAP7_75t_SL _26451_ (.A1(_04076_),
    .A2(_04077_),
    .B(_03762_),
    .Y(_04078_));
 AOI21x1_ASAP7_75t_SL _26452_ (.A1(_04073_),
    .A2(_04078_),
    .B(_03840_),
    .Y(_04079_));
 OAI21x1_ASAP7_75t_SL _26453_ (.A1(_04079_),
    .A2(_04070_),
    .B(_03816_),
    .Y(_04080_));
 NAND2x1_ASAP7_75t_SL _26454_ (.A(_04080_),
    .B(_04065_),
    .Y(_04081_));
 OAI21x1_ASAP7_75t_SL _26455_ (.A1(_04033_),
    .A2(_04051_),
    .B(_04081_),
    .Y(_00114_));
 NAND2x1_ASAP7_75t_SL _26456_ (.A(_04052_),
    .B(_03793_),
    .Y(_04082_));
 AOI21x1_ASAP7_75t_SL _26457_ (.A1(_03791_),
    .A2(_03800_),
    .B(_03784_),
    .Y(_04083_));
 NAND2x1_ASAP7_75t_SL _26458_ (.A(_04082_),
    .B(_04083_),
    .Y(_04084_));
 INVx1_ASAP7_75t_SL _26459_ (.A(_04025_),
    .Y(_04085_));
 OA21x2_ASAP7_75t_SL _26460_ (.A1(_03922_),
    .A2(_03747_),
    .B(_03784_),
    .Y(_04086_));
 NAND2x1_ASAP7_75t_SL _26461_ (.A(_04085_),
    .B(_04086_),
    .Y(_04087_));
 AOI21x1_ASAP7_75t_SL _26462_ (.A1(_04084_),
    .A2(_04087_),
    .B(_03762_),
    .Y(_04088_));
 OR3x1_ASAP7_75t_SL _26463_ (.A(_03784_),
    .B(_03747_),
    .C(_03829_),
    .Y(_04089_));
 NAND2x1_ASAP7_75t_SL _26464_ (.A(_03880_),
    .B(_04089_),
    .Y(_04090_));
 NAND2x1_ASAP7_75t_SL _26465_ (.A(_03903_),
    .B(_03901_),
    .Y(_04091_));
 OR3x1_ASAP7_75t_SL _26466_ (.A(_03840_),
    .B(_03791_),
    .C(_03753_),
    .Y(_04092_));
 OAI21x1_ASAP7_75t_SL _26467_ (.A1(_03784_),
    .A2(_04091_),
    .B(_04092_),
    .Y(_04093_));
 OAI21x1_ASAP7_75t_SL _26468_ (.A1(_04090_),
    .A2(_04093_),
    .B(_03808_),
    .Y(_04094_));
 NOR2x1_ASAP7_75t_SL _26469_ (.A(_04088_),
    .B(_04094_),
    .Y(_04095_));
 NAND2x1_ASAP7_75t_SL _26470_ (.A(_03993_),
    .B(_03891_),
    .Y(_04096_));
 NOR2x1_ASAP7_75t_R _26471_ (.A(_03731_),
    .B(_01282_),
    .Y(_04097_));
 OAI21x1_ASAP7_75t_SL _26472_ (.A1(_04015_),
    .A2(_04097_),
    .B(_03753_),
    .Y(_04098_));
 OAI21x1_ASAP7_75t_SL _26473_ (.A1(_03853_),
    .A2(_04020_),
    .B(_03747_),
    .Y(_04099_));
 NAND3x1_ASAP7_75t_SL _26474_ (.A(_04098_),
    .B(_04099_),
    .C(_03762_),
    .Y(_04100_));
 NAND2x1_ASAP7_75t_SL _26475_ (.A(_04096_),
    .B(_04100_),
    .Y(_04101_));
 INVx1_ASAP7_75t_SL _26476_ (.A(_03967_),
    .Y(_04102_));
 AOI21x1_ASAP7_75t_SL _26477_ (.A1(_01284_),
    .A2(_03721_),
    .B(_03747_),
    .Y(_04103_));
 NAND2x1_ASAP7_75t_SL _26478_ (.A(_04052_),
    .B(_04103_),
    .Y(_04104_));
 AOI21x1_ASAP7_75t_SL _26479_ (.A1(_04102_),
    .A2(_04104_),
    .B(_03762_),
    .Y(_04105_));
 OAI21x1_ASAP7_75t_SL _26480_ (.A1(_04020_),
    .A2(_03961_),
    .B(_03762_),
    .Y(_04106_));
 NAND2x1_ASAP7_75t_SL _26481_ (.A(_03840_),
    .B(_04106_),
    .Y(_04107_));
 OAI21x1_ASAP7_75t_SL _26482_ (.A1(_04105_),
    .A2(_04107_),
    .B(_03809_),
    .Y(_04108_));
 AOI21x1_ASAP7_75t_SL _26483_ (.A1(_03784_),
    .A2(_04101_),
    .B(_04108_),
    .Y(_04109_));
 OAI21x1_ASAP7_75t_SL _26484_ (.A1(_04095_),
    .A2(_04109_),
    .B(_03816_),
    .Y(_04110_));
 NOR2x1_ASAP7_75t_SL _26485_ (.A(_03939_),
    .B(_03830_),
    .Y(_04111_));
 NOR2x1_ASAP7_75t_SL _26486_ (.A(_03849_),
    .B(_03986_),
    .Y(_04112_));
 OAI21x1_ASAP7_75t_SL _26487_ (.A1(_04111_),
    .A2(_04112_),
    .B(_03762_),
    .Y(_04113_));
 AOI21x1_ASAP7_75t_SL _26488_ (.A1(_03721_),
    .A2(_01275_),
    .B(_03753_),
    .Y(_04114_));
 AOI21x1_ASAP7_75t_SL _26489_ (.A1(_03820_),
    .A2(_04114_),
    .B(_03762_),
    .Y(_04115_));
 OAI21x1_ASAP7_75t_SL _26490_ (.A1(_03734_),
    .A2(_04013_),
    .B(_04115_),
    .Y(_04116_));
 AOI21x1_ASAP7_75t_SL _26492_ (.A1(_04113_),
    .A2(_04116_),
    .B(_03809_),
    .Y(_04118_));
 AO21x1_ASAP7_75t_SL _26493_ (.A1(_03791_),
    .A2(_03824_),
    .B(_03753_),
    .Y(_04119_));
 NOR2x1_ASAP7_75t_R _26494_ (.A(_01282_),
    .B(_01275_),
    .Y(_04120_));
 OAI21x1_ASAP7_75t_SL _26495_ (.A1(_03935_),
    .A2(_04120_),
    .B(_03753_),
    .Y(_04121_));
 AOI21x1_ASAP7_75t_SL _26496_ (.A1(_04119_),
    .A2(_04121_),
    .B(_03763_),
    .Y(_04122_));
 OAI21x1_ASAP7_75t_SL _26497_ (.A1(_03849_),
    .A2(_03991_),
    .B(_03753_),
    .Y(_04123_));
 AO21x1_ASAP7_75t_SL _26498_ (.A1(_03894_),
    .A2(_03966_),
    .B(_03753_),
    .Y(_04124_));
 AOI21x1_ASAP7_75t_SL _26499_ (.A1(_04123_),
    .A2(_04124_),
    .B(_03762_),
    .Y(_04125_));
 NOR3x1_ASAP7_75t_SL _26500_ (.A(_04125_),
    .B(_04122_),
    .C(_03808_),
    .Y(_04126_));
 OAI21x1_ASAP7_75t_SL _26501_ (.A1(_04126_),
    .A2(_04118_),
    .B(_03784_),
    .Y(_04127_));
 OAI21x1_ASAP7_75t_SL _26502_ (.A1(_03935_),
    .A2(_03859_),
    .B(_03747_),
    .Y(_04128_));
 NAND2x1_ASAP7_75t_SL _26503_ (.A(_03763_),
    .B(_04128_),
    .Y(_04129_));
 AOI21x1_ASAP7_75t_R _26504_ (.A1(_01284_),
    .A2(_03721_),
    .B(_03753_),
    .Y(_04130_));
 NAND2x1_ASAP7_75t_SL _26505_ (.A(_03820_),
    .B(_04130_),
    .Y(_04131_));
 AOI21x1_ASAP7_75t_SL _26506_ (.A1(_04131_),
    .A2(_04008_),
    .B(_03808_),
    .Y(_04132_));
 OAI21x1_ASAP7_75t_SL _26507_ (.A1(_03954_),
    .A2(_04129_),
    .B(_04132_),
    .Y(_04133_));
 NAND2x1_ASAP7_75t_SL _26508_ (.A(_03789_),
    .B(_04114_),
    .Y(_04134_));
 AND2x2_ASAP7_75t_SL _26509_ (.A(_03830_),
    .B(_03762_),
    .Y(_04135_));
 AOI21x1_ASAP7_75t_SL _26510_ (.A1(_04134_),
    .A2(_04135_),
    .B(_03809_),
    .Y(_04136_));
 OAI21x1_ASAP7_75t_SL _26511_ (.A1(_03853_),
    .A2(_03960_),
    .B(_03753_),
    .Y(_04137_));
 NAND3x1_ASAP7_75t_SL _26512_ (.A(_04128_),
    .B(_04137_),
    .C(_03763_),
    .Y(_04138_));
 AOI21x1_ASAP7_75t_SL _26513_ (.A1(_04136_),
    .A2(_04138_),
    .B(_03784_),
    .Y(_04139_));
 AOI21x1_ASAP7_75t_SL _26514_ (.A1(_04133_),
    .A2(_04139_),
    .B(_03816_),
    .Y(_04140_));
 NAND2x1_ASAP7_75t_SL _26515_ (.A(_04127_),
    .B(_04140_),
    .Y(_04141_));
 NAND2x1_ASAP7_75t_SL _26516_ (.A(_04110_),
    .B(_04141_),
    .Y(_00115_));
 AND2x2_ASAP7_75t_SL _26517_ (.A(_03872_),
    .B(_03931_),
    .Y(_04142_));
 NAND2x1_ASAP7_75t_SL _26518_ (.A(_03762_),
    .B(_04066_),
    .Y(_04143_));
 AO21x1_ASAP7_75t_SL _26519_ (.A1(_04043_),
    .A2(_03823_),
    .B(_03747_),
    .Y(_04144_));
 AOI21x1_ASAP7_75t_SL _26520_ (.A1(_03978_),
    .A2(_04144_),
    .B(_03784_),
    .Y(_04145_));
 OAI21x1_ASAP7_75t_SL _26521_ (.A1(_04142_),
    .A2(_04143_),
    .B(_04145_),
    .Y(_04146_));
 AOI21x1_ASAP7_75t_R _26522_ (.A1(_01286_),
    .A2(_03731_),
    .B(_03753_),
    .Y(_04147_));
 NAND2x1_ASAP7_75t_SL _26523_ (.A(_03829_),
    .B(_04147_),
    .Y(_04148_));
 AOI21x1_ASAP7_75t_SL _26524_ (.A1(_04148_),
    .A2(_03873_),
    .B(_03840_),
    .Y(_04149_));
 AO21x1_ASAP7_75t_SL _26525_ (.A1(_03922_),
    .A2(_03914_),
    .B(_03753_),
    .Y(_04150_));
 INVx2_ASAP7_75t_SL _26526_ (.A(_03942_),
    .Y(_04151_));
 AOI21x1_ASAP7_75t_SL _26527_ (.A1(_03753_),
    .A2(_04015_),
    .B(_03763_),
    .Y(_04152_));
 NAND3x1_ASAP7_75t_SL _26528_ (.A(_04150_),
    .B(_04151_),
    .C(_04152_),
    .Y(_04153_));
 AOI21x1_ASAP7_75t_SL _26529_ (.A1(_04149_),
    .A2(_04153_),
    .B(_03809_),
    .Y(_04154_));
 NAND2x1_ASAP7_75t_SL _26530_ (.A(_04146_),
    .B(_04154_),
    .Y(_04155_));
 NAND2x1_ASAP7_75t_SL _26531_ (.A(_01282_),
    .B(_01279_),
    .Y(_04156_));
 AOI21x1_ASAP7_75t_SL _26532_ (.A1(_03751_),
    .A2(_04156_),
    .B(_03753_),
    .Y(_04157_));
 AND2x2_ASAP7_75t_SL _26533_ (.A(_04038_),
    .B(_03818_),
    .Y(_04158_));
 OAI21x1_ASAP7_75t_SL _26534_ (.A1(_04157_),
    .A2(_04158_),
    .B(_03762_),
    .Y(_04159_));
 INVx1_ASAP7_75t_SL _26535_ (.A(_03962_),
    .Y(_04160_));
 AOI21x1_ASAP7_75t_SL _26536_ (.A1(_04160_),
    .A2(_04039_),
    .B(_03784_),
    .Y(_04161_));
 NAND2x1_ASAP7_75t_SL _26537_ (.A(_04159_),
    .B(_04161_),
    .Y(_04162_));
 NAND2x1_ASAP7_75t_SL _26538_ (.A(_03762_),
    .B(_03879_),
    .Y(_04163_));
 OA21x2_ASAP7_75t_SL _26539_ (.A1(_04163_),
    .A2(_04103_),
    .B(_03784_),
    .Y(_04164_));
 INVx1_ASAP7_75t_SL _26540_ (.A(_03904_),
    .Y(_04165_));
 AOI21x1_ASAP7_75t_SL _26541_ (.A1(_03956_),
    .A2(_03789_),
    .B(_03762_),
    .Y(_04166_));
 OAI21x1_ASAP7_75t_SL _26542_ (.A1(_03960_),
    .A2(_04165_),
    .B(_04166_),
    .Y(_04167_));
 AOI21x1_ASAP7_75t_SL _26543_ (.A1(_04164_),
    .A2(_04167_),
    .B(_03808_),
    .Y(_04168_));
 AOI21x1_ASAP7_75t_SL _26544_ (.A1(_04162_),
    .A2(_04168_),
    .B(_03816_),
    .Y(_04169_));
 NAND2x1_ASAP7_75t_SL _26545_ (.A(_04155_),
    .B(_04169_),
    .Y(_04170_));
 AND3x1_ASAP7_75t_SL _26546_ (.A(_03985_),
    .B(_03747_),
    .C(_03894_),
    .Y(_04171_));
 INVx1_ASAP7_75t_SL _26547_ (.A(_03916_),
    .Y(_04172_));
 NOR2x1_ASAP7_75t_SL _26548_ (.A(_04171_),
    .B(_04172_),
    .Y(_04173_));
 NOR2x1_ASAP7_75t_SL _26549_ (.A(_03763_),
    .B(_03949_),
    .Y(_04174_));
 AO21x1_ASAP7_75t_SL _26550_ (.A1(_04174_),
    .A2(_04071_),
    .B(_03840_),
    .Y(_04175_));
 AND2x2_ASAP7_75t_SL _26551_ (.A(_03889_),
    .B(_03763_),
    .Y(_04176_));
 NAND2x1_ASAP7_75t_SL _26552_ (.A(_01286_),
    .B(_03721_),
    .Y(_04177_));
 NAND2x1_ASAP7_75t_SL _26553_ (.A(_04177_),
    .B(_03858_),
    .Y(_04178_));
 AOI21x1_ASAP7_75t_SL _26554_ (.A1(_04176_),
    .A2(_04178_),
    .B(_03784_),
    .Y(_04179_));
 OA21x2_ASAP7_75t_SL _26555_ (.A1(_03823_),
    .A2(_03753_),
    .B(_03762_),
    .Y(_04180_));
 NAND2x1_ASAP7_75t_SL _26556_ (.A(_03931_),
    .B(_03798_),
    .Y(_04181_));
 NAND3x1_ASAP7_75t_SL _26557_ (.A(_04180_),
    .B(_04181_),
    .C(_03831_),
    .Y(_04182_));
 AOI21x1_ASAP7_75t_SL _26558_ (.A1(_04179_),
    .A2(_04182_),
    .B(_03808_),
    .Y(_04183_));
 OAI21x1_ASAP7_75t_SL _26559_ (.A1(_04173_),
    .A2(_04175_),
    .B(_04183_),
    .Y(_04184_));
 NAND2x1_ASAP7_75t_SL _26560_ (.A(_03751_),
    .B(_04103_),
    .Y(_04185_));
 OA21x2_ASAP7_75t_R _26561_ (.A1(_03875_),
    .A2(_03753_),
    .B(_03762_),
    .Y(_04186_));
 NAND2x1_ASAP7_75t_SL _26562_ (.A(_04185_),
    .B(_04186_),
    .Y(_04187_));
 NAND2x1_ASAP7_75t_R _26563_ (.A(_01285_),
    .B(_03747_),
    .Y(_04188_));
 NAND2x1_ASAP7_75t_SL _26564_ (.A(_04034_),
    .B(_04188_),
    .Y(_04189_));
 OA21x2_ASAP7_75t_SL _26565_ (.A1(_04189_),
    .A2(_03762_),
    .B(_03784_),
    .Y(_04190_));
 AOI21x1_ASAP7_75t_SL _26566_ (.A1(_04187_),
    .A2(_04190_),
    .B(_03809_),
    .Y(_04191_));
 INVx1_ASAP7_75t_SL _26567_ (.A(_03863_),
    .Y(_04192_));
 OAI21x1_ASAP7_75t_R _26568_ (.A1(_03859_),
    .A2(_04192_),
    .B(_03753_),
    .Y(_04193_));
 AOI21x1_ASAP7_75t_SL _26569_ (.A1(_03909_),
    .A2(_04193_),
    .B(_03762_),
    .Y(_04194_));
 NAND2x1_ASAP7_75t_R _26570_ (.A(_03863_),
    .B(_04103_),
    .Y(_04195_));
 INVx1_ASAP7_75t_R _26571_ (.A(_04157_),
    .Y(_04196_));
 AOI21x1_ASAP7_75t_SL _26572_ (.A1(_04195_),
    .A2(_04196_),
    .B(_03763_),
    .Y(_04197_));
 OAI21x1_ASAP7_75t_SL _26573_ (.A1(_04194_),
    .A2(_04197_),
    .B(_03840_),
    .Y(_04198_));
 AOI21x1_ASAP7_75t_SL _26574_ (.A1(_04198_),
    .A2(_04191_),
    .B(_03929_),
    .Y(_04199_));
 NAND2x1_ASAP7_75t_SL _26575_ (.A(_04199_),
    .B(_04184_),
    .Y(_04200_));
 NAND2x1_ASAP7_75t_SL _26576_ (.A(_04200_),
    .B(_04170_),
    .Y(_00116_));
 AOI21x1_ASAP7_75t_SL _26577_ (.A1(_03753_),
    .A2(_04052_),
    .B(_03762_),
    .Y(_04201_));
 NAND2x1_ASAP7_75t_SL _26578_ (.A(_03774_),
    .B(_03755_),
    .Y(_04202_));
 NAND2x1_ASAP7_75t_SL _26579_ (.A(_04201_),
    .B(_04202_),
    .Y(_04203_));
 INVx1_ASAP7_75t_SL _26580_ (.A(_03793_),
    .Y(_04204_));
 AOI21x1_ASAP7_75t_SL _26581_ (.A1(_04204_),
    .A2(_03918_),
    .B(_03809_),
    .Y(_04205_));
 AOI21x1_ASAP7_75t_SL _26582_ (.A1(_04203_),
    .A2(_04205_),
    .B(_03840_),
    .Y(_04206_));
 NAND2x1_ASAP7_75t_SL _26583_ (.A(_03751_),
    .B(_04130_),
    .Y(_04207_));
 NAND2x1_ASAP7_75t_SL _26584_ (.A(_03791_),
    .B(_03954_),
    .Y(_04208_));
 AOI21x1_ASAP7_75t_SL _26585_ (.A1(_04207_),
    .A2(_04208_),
    .B(_03763_),
    .Y(_04209_));
 NAND2x1_ASAP7_75t_SL _26586_ (.A(_03753_),
    .B(_01282_),
    .Y(_04210_));
 AOI21x1_ASAP7_75t_SL _26587_ (.A1(_04210_),
    .A2(_03861_),
    .B(_03762_),
    .Y(_04211_));
 OAI21x1_ASAP7_75t_SL _26588_ (.A1(_04209_),
    .A2(_04211_),
    .B(_03809_),
    .Y(_04212_));
 NAND2x1_ASAP7_75t_SL _26589_ (.A(_04206_),
    .B(_04212_),
    .Y(_04213_));
 OA21x2_ASAP7_75t_SL _26590_ (.A1(_04192_),
    .A2(_04016_),
    .B(_03747_),
    .Y(_04214_));
 INVx1_ASAP7_75t_R _26591_ (.A(_03966_),
    .Y(_04215_));
 OAI21x1_ASAP7_75t_SL _26592_ (.A1(_04215_),
    .A2(_04020_),
    .B(_03747_),
    .Y(_04216_));
 OA21x2_ASAP7_75t_SL _26593_ (.A1(_03824_),
    .A2(_03747_),
    .B(_03762_),
    .Y(_04217_));
 AOI21x1_ASAP7_75t_SL _26594_ (.A1(_04216_),
    .A2(_04217_),
    .B(_03808_),
    .Y(_04218_));
 OAI21x1_ASAP7_75t_SL _26595_ (.A1(_04172_),
    .A2(_04214_),
    .B(_04218_),
    .Y(_04219_));
 AO21x1_ASAP7_75t_SL _26596_ (.A1(_03731_),
    .A2(_03773_),
    .B(_03753_),
    .Y(_04220_));
 OA21x2_ASAP7_75t_SL _26597_ (.A1(_03848_),
    .A2(_03747_),
    .B(_03763_),
    .Y(_04221_));
 AOI21x1_ASAP7_75t_SL _26598_ (.A1(_04220_),
    .A2(_04221_),
    .B(_03809_),
    .Y(_04222_));
 NAND2x1_ASAP7_75t_SL _26599_ (.A(_03903_),
    .B(_03919_),
    .Y(_04223_));
 AOI21x1_ASAP7_75t_SL _26600_ (.A1(_03747_),
    .A2(_04020_),
    .B(_03833_),
    .Y(_04224_));
 NAND2x1_ASAP7_75t_SL _26601_ (.A(_04223_),
    .B(_04224_),
    .Y(_04225_));
 AOI21x1_ASAP7_75t_SL _26602_ (.A1(_04222_),
    .A2(_04225_),
    .B(_03784_),
    .Y(_04226_));
 NAND2x1_ASAP7_75t_SL _26603_ (.A(_04219_),
    .B(_04226_),
    .Y(_04227_));
 AOI21x1_ASAP7_75t_SL _26604_ (.A1(_04213_),
    .A2(_04227_),
    .B(_03929_),
    .Y(_04228_));
 AO21x1_ASAP7_75t_SL _26605_ (.A1(_03949_),
    .A2(_04059_),
    .B(_03942_),
    .Y(_04229_));
 AOI21x1_ASAP7_75t_SL _26606_ (.A1(_03762_),
    .A2(_04229_),
    .B(_03809_),
    .Y(_04230_));
 AO221x1_ASAP7_75t_SL _26607_ (.A1(_03747_),
    .A2(_04029_),
    .B1(_03818_),
    .B2(_03919_),
    .C(_03762_),
    .Y(_04231_));
 AOI21x1_ASAP7_75t_SL _26608_ (.A1(_03747_),
    .A2(_03985_),
    .B(_03991_),
    .Y(_04232_));
 OAI21x1_ASAP7_75t_SL _26609_ (.A1(_03763_),
    .A2(_04232_),
    .B(_03809_),
    .Y(_04233_));
 NAND2x1_ASAP7_75t_SL _26610_ (.A(_03747_),
    .B(_03791_),
    .Y(_04234_));
 AOI21x1_ASAP7_75t_SL _26611_ (.A1(_04234_),
    .A2(_04098_),
    .B(_03762_),
    .Y(_04235_));
 OAI21x1_ASAP7_75t_SL _26612_ (.A1(_04233_),
    .A2(_04235_),
    .B(_03840_),
    .Y(_04236_));
 AOI21x1_ASAP7_75t_SL _26613_ (.A1(_04231_),
    .A2(_04230_),
    .B(_04236_),
    .Y(_04237_));
 AO21x1_ASAP7_75t_SL _26614_ (.A1(_03966_),
    .A2(_03824_),
    .B(_03747_),
    .Y(_04238_));
 OAI21x1_ASAP7_75t_SL _26615_ (.A1(_04097_),
    .A2(_03997_),
    .B(_03747_),
    .Y(_04239_));
 AOI21x1_ASAP7_75t_SL _26616_ (.A1(_04238_),
    .A2(_04239_),
    .B(_03763_),
    .Y(_04240_));
 AO21x1_ASAP7_75t_SL _26617_ (.A1(_01275_),
    .A2(_03753_),
    .B(_03762_),
    .Y(_04241_));
 OAI21x1_ASAP7_75t_SL _26618_ (.A1(_04241_),
    .A2(_04157_),
    .B(_03808_),
    .Y(_04242_));
 OAI21x1_ASAP7_75t_SL _26619_ (.A1(_04240_),
    .A2(_04242_),
    .B(_03784_),
    .Y(_04243_));
 NAND2x1_ASAP7_75t_SL _26620_ (.A(_04046_),
    .B(_04130_),
    .Y(_04244_));
 AO21x1_ASAP7_75t_SL _26621_ (.A1(_03731_),
    .A2(_03878_),
    .B(_03913_),
    .Y(_04245_));
 AOI21x1_ASAP7_75t_SL _26622_ (.A1(_03753_),
    .A2(_04245_),
    .B(_03763_),
    .Y(_04246_));
 NAND2x1_ASAP7_75t_SL _26623_ (.A(_04244_),
    .B(_04246_),
    .Y(_04247_));
 NAND2x1_ASAP7_75t_SL _26624_ (.A(_03985_),
    .B(_03793_),
    .Y(_04248_));
 NAND3x1_ASAP7_75t_SL _26625_ (.A(_03772_),
    .B(_04248_),
    .C(_03763_),
    .Y(_04249_));
 AOI21x1_ASAP7_75t_SL _26626_ (.A1(_04247_),
    .A2(_04249_),
    .B(_03808_),
    .Y(_04250_));
 OAI21x1_ASAP7_75t_SL _26627_ (.A1(_04243_),
    .A2(_04250_),
    .B(_03929_),
    .Y(_04251_));
 NOR2x1_ASAP7_75t_SL _26628_ (.A(_04251_),
    .B(_04237_),
    .Y(_04252_));
 NOR2x1_ASAP7_75t_SL _26629_ (.A(_04228_),
    .B(_04252_),
    .Y(_00117_));
 INVx1_ASAP7_75t_SL _26630_ (.A(_03981_),
    .Y(_04253_));
 AOI21x1_ASAP7_75t_SL _26631_ (.A1(_04253_),
    .A2(_03790_),
    .B(_03763_),
    .Y(_04254_));
 NAND2x1_ASAP7_75t_SL _26632_ (.A(_03747_),
    .B(_03853_),
    .Y(_04255_));
 AOI21x1_ASAP7_75t_SL _26633_ (.A1(_04255_),
    .A2(_04098_),
    .B(_03762_),
    .Y(_04256_));
 OAI21x1_ASAP7_75t_SL _26634_ (.A1(_04254_),
    .A2(_04256_),
    .B(_03840_),
    .Y(_04257_));
 NAND2x1_ASAP7_75t_SL _26635_ (.A(_04059_),
    .B(_03755_),
    .Y(_04258_));
 OAI21x1_ASAP7_75t_SL _26636_ (.A1(_03935_),
    .A2(_03859_),
    .B(_03753_),
    .Y(_04259_));
 AOI21x1_ASAP7_75t_SL _26637_ (.A1(_04258_),
    .A2(_04259_),
    .B(_03762_),
    .Y(_04260_));
 INVx1_ASAP7_75t_SL _26638_ (.A(_03935_),
    .Y(_04261_));
 NAND2x1_ASAP7_75t_SL _26639_ (.A(_04147_),
    .B(_04261_),
    .Y(_04262_));
 OAI21x1_ASAP7_75t_SL _26640_ (.A1(_04120_),
    .A2(_04192_),
    .B(_03753_),
    .Y(_04263_));
 AOI21x1_ASAP7_75t_SL _26641_ (.A1(_04262_),
    .A2(_04263_),
    .B(_03763_),
    .Y(_04264_));
 OAI21x1_ASAP7_75t_SL _26642_ (.A1(_04260_),
    .A2(_04264_),
    .B(_03784_),
    .Y(_04265_));
 NAND2x1_ASAP7_75t_SL _26643_ (.A(_04257_),
    .B(_04265_),
    .Y(_04266_));
 INVx1_ASAP7_75t_SL _26644_ (.A(_04068_),
    .Y(_04267_));
 AO21x1_ASAP7_75t_SL _26645_ (.A1(_03721_),
    .A2(_03848_),
    .B(_03753_),
    .Y(_04268_));
 AOI21x1_ASAP7_75t_SL _26646_ (.A1(_04268_),
    .A2(_04185_),
    .B(_03763_),
    .Y(_04269_));
 OAI21x1_ASAP7_75t_SL _26647_ (.A1(_04267_),
    .A2(_04269_),
    .B(_03840_),
    .Y(_04270_));
 AOI21x1_ASAP7_75t_SL _26648_ (.A1(_01289_),
    .A2(_03753_),
    .B(_03762_),
    .Y(_04271_));
 AOI21x1_ASAP7_75t_SL _26649_ (.A1(_04271_),
    .A2(_04207_),
    .B(_03840_),
    .Y(_04272_));
 AOI21x1_ASAP7_75t_SL _26650_ (.A1(_03820_),
    .A2(_04177_),
    .B(_03747_),
    .Y(_04273_));
 OAI21x1_ASAP7_75t_SL _26651_ (.A1(_03987_),
    .A2(_04273_),
    .B(_03762_),
    .Y(_04274_));
 AOI21x1_ASAP7_75t_SL _26652_ (.A1(_04272_),
    .A2(_04274_),
    .B(_03809_),
    .Y(_04275_));
 AOI21x1_ASAP7_75t_SL _26653_ (.A1(_04270_),
    .A2(_04275_),
    .B(_03929_),
    .Y(_04276_));
 OAI21x1_ASAP7_75t_SL _26654_ (.A1(_03808_),
    .A2(_04266_),
    .B(_04276_),
    .Y(_04277_));
 NAND2x1_ASAP7_75t_SL _26655_ (.A(_03872_),
    .B(_04261_),
    .Y(_04278_));
 NAND3x1_ASAP7_75t_SL _26656_ (.A(_03894_),
    .B(_03747_),
    .C(_04052_),
    .Y(_04279_));
 AOI21x1_ASAP7_75t_SL _26657_ (.A1(_04278_),
    .A2(_04279_),
    .B(_03762_),
    .Y(_04280_));
 NOR2x1_ASAP7_75t_SL _26658_ (.A(_03753_),
    .B(_03824_),
    .Y(_04281_));
 AOI21x1_ASAP7_75t_SL _26659_ (.A1(_04043_),
    .A2(_03872_),
    .B(_04281_),
    .Y(_04282_));
 OAI21x1_ASAP7_75t_SL _26660_ (.A1(_03763_),
    .A2(_04282_),
    .B(_03840_),
    .Y(_04283_));
 NOR2x1_ASAP7_75t_SL _26661_ (.A(_04280_),
    .B(_04283_),
    .Y(_04284_));
 NAND2x1_ASAP7_75t_SL _26662_ (.A(_03751_),
    .B(_03954_),
    .Y(_04285_));
 INVx1_ASAP7_75t_SL _26663_ (.A(_03791_),
    .Y(_04286_));
 OAI21x1_ASAP7_75t_SL _26664_ (.A1(_04286_),
    .A2(_04074_),
    .B(_03747_),
    .Y(_04287_));
 AOI21x1_ASAP7_75t_SL _26665_ (.A1(_04285_),
    .A2(_04287_),
    .B(_03762_),
    .Y(_04288_));
 OAI21x1_ASAP7_75t_SL _26666_ (.A1(_03833_),
    .A2(_04062_),
    .B(_03784_),
    .Y(_04289_));
 OAI21x1_ASAP7_75t_SL _26667_ (.A1(_04288_),
    .A2(_04289_),
    .B(_03808_),
    .Y(_04290_));
 NOR2x1_ASAP7_75t_SL _26668_ (.A(_04284_),
    .B(_04290_),
    .Y(_04291_));
 OAI21x1_ASAP7_75t_SL _26669_ (.A1(_04015_),
    .A2(_04074_),
    .B(_03753_),
    .Y(_04292_));
 AOI21x1_ASAP7_75t_SL _26670_ (.A1(_04180_),
    .A2(_04292_),
    .B(_03840_),
    .Y(_04293_));
 AO21x1_ASAP7_75t_SL _26671_ (.A1(_01288_),
    .A2(_01294_),
    .B(_03753_),
    .Y(_04294_));
 AND2x2_ASAP7_75t_SL _26672_ (.A(_04294_),
    .B(_03763_),
    .Y(_04295_));
 AO21x1_ASAP7_75t_SL _26673_ (.A1(_03751_),
    .A2(_04156_),
    .B(_03747_),
    .Y(_04296_));
 NAND2x1_ASAP7_75t_SL _26674_ (.A(_04295_),
    .B(_04296_),
    .Y(_04297_));
 NAND2x1_ASAP7_75t_SL _26675_ (.A(_04293_),
    .B(_04297_),
    .Y(_04298_));
 NAND2x1_ASAP7_75t_SL _26676_ (.A(_04130_),
    .B(_03735_),
    .Y(_04299_));
 OAI21x1_ASAP7_75t_SL _26677_ (.A1(_03767_),
    .A2(_03852_),
    .B(_03753_),
    .Y(_04300_));
 AOI21x1_ASAP7_75t_SL _26678_ (.A1(_04299_),
    .A2(_04300_),
    .B(_03762_),
    .Y(_04301_));
 NAND2x1_ASAP7_75t_SL _26679_ (.A(_03858_),
    .B(_03894_),
    .Y(_04302_));
 OAI21x1_ASAP7_75t_SL _26680_ (.A1(_04015_),
    .A2(_03886_),
    .B(_03753_),
    .Y(_04303_));
 AOI21x1_ASAP7_75t_SL _26681_ (.A1(_04303_),
    .A2(_04302_),
    .B(_03763_),
    .Y(_04304_));
 OAI21x1_ASAP7_75t_SL _26682_ (.A1(_04304_),
    .A2(_04301_),
    .B(_03840_),
    .Y(_04305_));
 AOI21x1_ASAP7_75t_SL _26683_ (.A1(_04298_),
    .A2(_04305_),
    .B(_03808_),
    .Y(_04306_));
 OAI21x1_ASAP7_75t_SL _26684_ (.A1(_04306_),
    .A2(_04291_),
    .B(_03929_),
    .Y(_04307_));
 NAND2x1_ASAP7_75t_SL _26685_ (.A(_04277_),
    .B(_04307_),
    .Y(_00118_));
 NAND2x1_ASAP7_75t_SL _26686_ (.A(_03753_),
    .B(_04215_),
    .Y(_04308_));
 OA21x2_ASAP7_75t_SL _26687_ (.A1(_03791_),
    .A2(_03753_),
    .B(_03763_),
    .Y(_04309_));
 AOI21x1_ASAP7_75t_SL _26688_ (.A1(_04308_),
    .A2(_04309_),
    .B(_03784_),
    .Y(_04310_));
 NOR2x1_ASAP7_75t_SL _26689_ (.A(_03763_),
    .B(_03872_),
    .Y(_04311_));
 OA21x2_ASAP7_75t_SL _26690_ (.A1(_03731_),
    .A2(_01285_),
    .B(_03747_),
    .Y(_04312_));
 NAND2x1_ASAP7_75t_SL _26691_ (.A(_03820_),
    .B(_04312_),
    .Y(_04313_));
 NAND2x1_ASAP7_75t_SL _26692_ (.A(_04311_),
    .B(_04313_),
    .Y(_04314_));
 AOI21x1_ASAP7_75t_SL _26693_ (.A1(_04310_),
    .A2(_04314_),
    .B(_03809_),
    .Y(_04315_));
 NOR2x1_ASAP7_75t_R _26694_ (.A(_03753_),
    .B(_01282_),
    .Y(_04316_));
 AO21x1_ASAP7_75t_SL _26695_ (.A1(_03904_),
    .A2(_04043_),
    .B(_04316_),
    .Y(_04317_));
 NAND2x1_ASAP7_75t_SL _26696_ (.A(_03762_),
    .B(_04317_),
    .Y(_04318_));
 NAND2x1_ASAP7_75t_SL _26697_ (.A(_03751_),
    .B(_04312_),
    .Y(_04319_));
 AOI21x1_ASAP7_75t_SL _26698_ (.A1(_04319_),
    .A2(_04039_),
    .B(_03840_),
    .Y(_04320_));
 NAND2x1_ASAP7_75t_SL _26699_ (.A(_04318_),
    .B(_04320_),
    .Y(_04321_));
 AOI21x1_ASAP7_75t_SL _26700_ (.A1(_04315_),
    .A2(_04321_),
    .B(_03929_),
    .Y(_04322_));
 NAND2x1_ASAP7_75t_SL _26701_ (.A(_03976_),
    .B(_04083_),
    .Y(_04323_));
 NAND2x1_ASAP7_75t_SL _26702_ (.A(_04046_),
    .B(_03800_),
    .Y(_04324_));
 OAI21x1_ASAP7_75t_R _26703_ (.A1(_03747_),
    .A2(_03823_),
    .B(_03784_),
    .Y(_04325_));
 NOR2x1_ASAP7_75t_R _26704_ (.A(_03773_),
    .B(_03889_),
    .Y(_04326_));
 NOR2x1_ASAP7_75t_SL _26705_ (.A(_04325_),
    .B(_04326_),
    .Y(_04327_));
 NAND2x1_ASAP7_75t_SL _26706_ (.A(_04324_),
    .B(_04327_),
    .Y(_04328_));
 AOI21x1_ASAP7_75t_SL _26707_ (.A1(_04323_),
    .A2(_04328_),
    .B(_03763_),
    .Y(_04329_));
 INVx1_ASAP7_75t_SL _26708_ (.A(_04147_),
    .Y(_04330_));
 AOI21x1_ASAP7_75t_SL _26709_ (.A1(_04330_),
    .A2(_04185_),
    .B(_03840_),
    .Y(_04331_));
 AND3x1_ASAP7_75t_SL _26710_ (.A(_03904_),
    .B(_03840_),
    .C(_03931_),
    .Y(_04332_));
 AO21x1_ASAP7_75t_SL _26711_ (.A1(_03735_),
    .A2(_04130_),
    .B(_03762_),
    .Y(_04333_));
 NOR3x1_ASAP7_75t_SL _26712_ (.A(_04331_),
    .B(_04332_),
    .C(_04333_),
    .Y(_04334_));
 OAI21x1_ASAP7_75t_SL _26713_ (.A1(_04329_),
    .A2(_04334_),
    .B(_03809_),
    .Y(_04335_));
 NAND2x1_ASAP7_75t_SL _26714_ (.A(_04322_),
    .B(_04335_),
    .Y(_04336_));
 AO21x1_ASAP7_75t_SL _26715_ (.A1(_03894_),
    .A2(_03791_),
    .B(_03747_),
    .Y(_04337_));
 NAND2x1_ASAP7_75t_SL _26716_ (.A(_03751_),
    .B(_03800_),
    .Y(_04338_));
 AOI21x1_ASAP7_75t_SL _26717_ (.A1(_04338_),
    .A2(_04337_),
    .B(_03763_),
    .Y(_04339_));
 AO21x1_ASAP7_75t_SL _26718_ (.A1(_01294_),
    .A2(_03753_),
    .B(_03762_),
    .Y(_04340_));
 AND3x1_ASAP7_75t_SL _26719_ (.A(_03922_),
    .B(_03747_),
    .C(_03829_),
    .Y(_04341_));
 OAI21x1_ASAP7_75t_SL _26720_ (.A1(_04340_),
    .A2(_04341_),
    .B(_03840_),
    .Y(_04342_));
 NOR2x1_ASAP7_75t_SL _26721_ (.A(_04342_),
    .B(_04339_),
    .Y(_04343_));
 AOI21x1_ASAP7_75t_SL _26722_ (.A1(_03747_),
    .A2(_04074_),
    .B(_03762_),
    .Y(_04344_));
 OAI21x1_ASAP7_75t_SL _26723_ (.A1(_03773_),
    .A2(_03747_),
    .B(_04344_),
    .Y(_04345_));
 NAND3x1_ASAP7_75t_SL _26724_ (.A(_04186_),
    .B(_04181_),
    .C(_03831_),
    .Y(_04346_));
 AOI21x1_ASAP7_75t_SL _26725_ (.A1(_04345_),
    .A2(_04346_),
    .B(_03840_),
    .Y(_04347_));
 OAI21x1_ASAP7_75t_SL _26726_ (.A1(_04347_),
    .A2(_04343_),
    .B(_03808_),
    .Y(_04348_));
 AO21x1_ASAP7_75t_SL _26727_ (.A1(_03791_),
    .A2(_03824_),
    .B(_03747_),
    .Y(_04349_));
 OAI21x1_ASAP7_75t_SL _26728_ (.A1(_03939_),
    .A2(_03852_),
    .B(_03747_),
    .Y(_04350_));
 AOI21x1_ASAP7_75t_SL _26729_ (.A1(_04349_),
    .A2(_04350_),
    .B(_03762_),
    .Y(_04351_));
 NAND2x1_ASAP7_75t_SL _26730_ (.A(_04059_),
    .B(_04312_),
    .Y(_04352_));
 AOI21x1_ASAP7_75t_SL _26731_ (.A1(_04104_),
    .A2(_04352_),
    .B(_03763_),
    .Y(_04353_));
 OAI21x1_ASAP7_75t_SL _26732_ (.A1(_04351_),
    .A2(_04353_),
    .B(_03784_),
    .Y(_04354_));
 OA21x2_ASAP7_75t_SL _26733_ (.A1(_01281_),
    .A2(_03753_),
    .B(_03762_),
    .Y(_04355_));
 NAND2x1_ASAP7_75t_SL _26734_ (.A(_04355_),
    .B(_04296_),
    .Y(_04356_));
 OA21x2_ASAP7_75t_SL _26735_ (.A1(_03889_),
    .A2(_01279_),
    .B(_03823_),
    .Y(_04357_));
 AOI21x1_ASAP7_75t_SL _26736_ (.A1(_04344_),
    .A2(_04357_),
    .B(_03784_),
    .Y(_04358_));
 AOI21x1_ASAP7_75t_SL _26737_ (.A1(_04356_),
    .A2(_04358_),
    .B(_03808_),
    .Y(_04359_));
 AOI21x1_ASAP7_75t_SL _26738_ (.A1(_04354_),
    .A2(_04359_),
    .B(_03816_),
    .Y(_04360_));
 NAND2x1_ASAP7_75t_SL _26739_ (.A(_04348_),
    .B(_04360_),
    .Y(_04361_));
 NAND2x1_ASAP7_75t_SL _26740_ (.A(_04336_),
    .B(_04361_),
    .Y(_00119_));
 AND2x2_ASAP7_75t_R _26741_ (.A(_10675_),
    .B(_00477_),
    .Y(_04362_));
 XOR2x2_ASAP7_75t_SL _26742_ (.A(_12805_),
    .B(_01585_),
    .Y(_04363_));
 XOR2x2_ASAP7_75t_SL _26743_ (.A(_00695_),
    .B(_00569_),
    .Y(_04364_));
 XOR2x2_ASAP7_75t_SL _26744_ (.A(_12772_),
    .B(_04364_),
    .Y(_04365_));
 XOR2x2_ASAP7_75t_SL _26745_ (.A(_04363_),
    .B(_04365_),
    .Y(_04366_));
 NOR2x1p5_ASAP7_75t_L _26746_ (.A(_10675_),
    .B(_04366_),
    .Y(_04367_));
 INVx1_ASAP7_75t_R _26747_ (.A(_00486_),
    .Y(_04368_));
 OAI21x1_ASAP7_75t_R _26748_ (.A1(_04362_),
    .A2(_04367_),
    .B(_04368_),
    .Y(_04369_));
 NOR2x1_ASAP7_75t_L _26749_ (.A(_00574_),
    .B(_00477_),
    .Y(_04370_));
 XNOR2x2_ASAP7_75t_SL _26750_ (.A(_04365_),
    .B(_04363_),
    .Y(_04371_));
 NOR2x1_ASAP7_75t_L _26751_ (.A(_10675_),
    .B(_04371_),
    .Y(_04372_));
 OAI21x1_ASAP7_75t_R _26752_ (.A1(_04370_),
    .A2(_04372_),
    .B(_00486_),
    .Y(_04373_));
 NAND2x2_ASAP7_75t_SL _26753_ (.A(_04369_),
    .B(_04373_),
    .Y(_01302_));
 NOR2x1_ASAP7_75t_L _26754_ (.A(_00574_),
    .B(_00478_),
    .Y(_04374_));
 XOR2x2_ASAP7_75t_SL _26755_ (.A(_00631_),
    .B(_00670_),
    .Y(_04375_));
 XOR2x2_ASAP7_75t_SL _26756_ (.A(_04375_),
    .B(_00599_),
    .Y(_04376_));
 NAND2x1_ASAP7_75t_R _26757_ (.A(_04364_),
    .B(_04376_),
    .Y(_04377_));
 INVx2_ASAP7_75t_R _26758_ (.A(_04364_),
    .Y(_04378_));
 INVx1_ASAP7_75t_R _26759_ (.A(_04376_),
    .Y(_04379_));
 NAND2x1_ASAP7_75t_R _26760_ (.A(_04378_),
    .B(_04379_),
    .Y(_04380_));
 AOI21x1_ASAP7_75t_SL _26761_ (.A1(_04377_),
    .A2(_04380_),
    .B(_10675_),
    .Y(_04381_));
 OAI21x1_ASAP7_75t_R _26762_ (.A1(_04374_),
    .A2(_04381_),
    .B(_00964_),
    .Y(_04382_));
 AND2x2_ASAP7_75t_R _26763_ (.A(_10675_),
    .B(_00478_),
    .Y(_04383_));
 XOR2x2_ASAP7_75t_SL _26764_ (.A(_04376_),
    .B(_04378_),
    .Y(_04384_));
 NOR2x1_ASAP7_75t_R _26765_ (.A(_10675_),
    .B(_04384_),
    .Y(_04385_));
 OAI21x1_ASAP7_75t_R _26766_ (.A1(_04383_),
    .A2(_04385_),
    .B(_08903_),
    .Y(_04386_));
 NAND2x1_ASAP7_75t_SL _26767_ (.A(_04382_),
    .B(_04386_),
    .Y(_01305_));
 NOR2x1_ASAP7_75t_R _26768_ (.A(_00574_),
    .B(_00479_),
    .Y(_04387_));
 INVx1_ASAP7_75t_SL _26769_ (.A(_04387_),
    .Y(_04388_));
 XOR2x2_ASAP7_75t_SL _26770_ (.A(_00601_),
    .B(_00633_),
    .Y(_04389_));
 INVx1_ASAP7_75t_SL _26771_ (.A(_04389_),
    .Y(_04390_));
 INVx1_ASAP7_75t_R _26772_ (.A(_00697_),
    .Y(_04391_));
 XOR2x2_ASAP7_75t_SL _26773_ (.A(_01581_),
    .B(_04391_),
    .Y(_04392_));
 NOR2x1_ASAP7_75t_R _26774_ (.A(_04390_),
    .B(_04392_),
    .Y(_04393_));
 AND2x2_ASAP7_75t_L _26775_ (.A(_04392_),
    .B(_04390_),
    .Y(_04394_));
 OAI21x1_ASAP7_75t_SL _26776_ (.A1(_04393_),
    .A2(_04394_),
    .B(_00574_),
    .Y(_04395_));
 INVx1_ASAP7_75t_R _26777_ (.A(_00935_),
    .Y(_04396_));
 AOI21x1_ASAP7_75t_R _26778_ (.A1(_04388_),
    .A2(_04395_),
    .B(_04396_),
    .Y(_04397_));
 NAND2x1_ASAP7_75t_R _26779_ (.A(_00479_),
    .B(_10675_),
    .Y(_04398_));
 XOR2x2_ASAP7_75t_SL _26780_ (.A(_04392_),
    .B(_04390_),
    .Y(_04399_));
 NAND2x1_ASAP7_75t_L _26781_ (.A(_00574_),
    .B(_04399_),
    .Y(_04400_));
 AOI21x1_ASAP7_75t_R _26782_ (.A1(_04398_),
    .A2(_04400_),
    .B(_00935_),
    .Y(_04401_));
 NOR2x1_ASAP7_75t_SL _26783_ (.A(_04397_),
    .B(_04401_),
    .Y(_04402_));
 OAI21x1_ASAP7_75t_SL _26786_ (.A1(_04367_),
    .A2(_04362_),
    .B(_00486_),
    .Y(_04404_));
 OAI21x1_ASAP7_75t_SL _26787_ (.A1(_04370_),
    .A2(_04372_),
    .B(_04368_),
    .Y(_04405_));
 NAND2x2_ASAP7_75t_SL _26788_ (.A(_04405_),
    .B(_04404_),
    .Y(_01298_));
 AOI21x1_ASAP7_75t_SL _26789_ (.A1(_04388_),
    .A2(_04395_),
    .B(_00935_),
    .Y(_04406_));
 AOI21x1_ASAP7_75t_SL _26790_ (.A1(_04398_),
    .A2(_04400_),
    .B(_04396_),
    .Y(_04407_));
 NOR2x1_ASAP7_75t_SL _26791_ (.A(_04406_),
    .B(_04407_),
    .Y(_04408_));
 NAND2x1_ASAP7_75t_R _26794_ (.A(_01299_),
    .B(_04402_),
    .Y(_04410_));
 NAND2x1_ASAP7_75t_SL _26796_ (.A(_01306_),
    .B(_04408_),
    .Y(_04412_));
 XNOR2x2_ASAP7_75t_SL _26797_ (.A(_00698_),
    .B(_01646_),
    .Y(_04413_));
 XNOR2x2_ASAP7_75t_L _26798_ (.A(_00569_),
    .B(_00697_),
    .Y(_04414_));
 XOR2x2_ASAP7_75t_R _26799_ (.A(_00602_),
    .B(_00634_),
    .Y(_04415_));
 XOR2x2_ASAP7_75t_SL _26800_ (.A(_04414_),
    .B(_04415_),
    .Y(_04416_));
 AOI21x1_ASAP7_75t_R _26801_ (.A1(_04413_),
    .A2(_04416_),
    .B(_10675_),
    .Y(_04417_));
 OR2x2_ASAP7_75t_SL _26802_ (.A(_04416_),
    .B(_04413_),
    .Y(_04418_));
 AND2x2_ASAP7_75t_R _26803_ (.A(_10675_),
    .B(_00554_),
    .Y(_04419_));
 AOI21x1_ASAP7_75t_SL _26804_ (.A1(_04417_),
    .A2(_04418_),
    .B(_04419_),
    .Y(_04420_));
 XOR2x2_ASAP7_75t_SL _26805_ (.A(_04420_),
    .B(_00936_),
    .Y(_04421_));
 AO21x1_ASAP7_75t_SL _26808_ (.A1(_04410_),
    .A2(_04412_),
    .B(_04421_),
    .Y(_04424_));
 NOR2x1_ASAP7_75t_SL _26809_ (.A(_10675_),
    .B(_04399_),
    .Y(_04425_));
 OAI21x1_ASAP7_75t_SL _26810_ (.A1(_04387_),
    .A2(_04425_),
    .B(_00935_),
    .Y(_04426_));
 NAND3x1_ASAP7_75t_SL _26811_ (.A(_04395_),
    .B(_04396_),
    .C(_04388_),
    .Y(_04427_));
 INVx2_ASAP7_75t_SL _26812_ (.A(_01300_),
    .Y(_04428_));
 AOI21x1_ASAP7_75t_SL _26813_ (.A1(_04426_),
    .A2(_04427_),
    .B(_04428_),
    .Y(_04429_));
 INVx2_ASAP7_75t_SL _26814_ (.A(_04429_),
    .Y(_04430_));
 INVx1_ASAP7_75t_SL _26815_ (.A(_01308_),
    .Y(_04431_));
 XOR2x2_ASAP7_75t_SL _26817_ (.A(_04420_),
    .B(_08920_),
    .Y(_04433_));
 AOI21x1_ASAP7_75t_R _26818_ (.A1(_04431_),
    .A2(_04402_),
    .B(_04433_),
    .Y(_04434_));
 NAND2x1_ASAP7_75t_SL _26819_ (.A(_04430_),
    .B(_04434_),
    .Y(_04435_));
 XOR2x2_ASAP7_75t_R _26820_ (.A(_00569_),
    .B(_00698_),
    .Y(_04436_));
 XOR2x2_ASAP7_75t_SL _26821_ (.A(_12872_),
    .B(_04436_),
    .Y(_04437_));
 XOR2x2_ASAP7_75t_SL _26822_ (.A(_04437_),
    .B(_01666_),
    .Y(_04438_));
 OR2x2_ASAP7_75t_R _26823_ (.A(_00574_),
    .B(_00548_),
    .Y(_04439_));
 OAI21x1_ASAP7_75t_R _26824_ (.A1(_10675_),
    .A2(_04438_),
    .B(_04439_),
    .Y(_04440_));
 XNOR2x2_ASAP7_75t_SL _26825_ (.A(_00937_),
    .B(_04440_),
    .Y(_04441_));
 AO21x1_ASAP7_75t_SL _26828_ (.A1(_04435_),
    .A2(_04424_),
    .B(_04441_),
    .Y(_04444_));
 NAND2x1_ASAP7_75t_SL _26829_ (.A(_01305_),
    .B(_04408_),
    .Y(_04445_));
 OAI21x1_ASAP7_75t_R _26830_ (.A1(_04374_),
    .A2(_04381_),
    .B(_08903_),
    .Y(_04446_));
 OAI21x1_ASAP7_75t_R _26831_ (.A1(_04383_),
    .A2(_04385_),
    .B(_00964_),
    .Y(_04447_));
 NAND2x1_ASAP7_75t_SL _26832_ (.A(_04446_),
    .B(_04447_),
    .Y(_04448_));
 NAND2x1_ASAP7_75t_SL _26833_ (.A(_04448_),
    .B(_01298_),
    .Y(_04449_));
 AOI21x1_ASAP7_75t_SL _26835_ (.A1(_04445_),
    .A2(_04449_),
    .B(_04421_),
    .Y(_04451_));
 INVx1_ASAP7_75t_SL _26836_ (.A(_04451_),
    .Y(_04452_));
 AOI21x1_ASAP7_75t_SL _26838_ (.A1(_01305_),
    .A2(_04408_),
    .B(_04433_),
    .Y(_04454_));
 NAND2x1_ASAP7_75t_SL _26839_ (.A(_04449_),
    .B(_04454_),
    .Y(_04455_));
 XOR2x2_ASAP7_75t_SL _26840_ (.A(_04440_),
    .B(_00937_),
    .Y(_04456_));
 AO21x1_ASAP7_75t_SL _26843_ (.A1(_04452_),
    .A2(_04455_),
    .B(_04456_),
    .Y(_04459_));
 XOR2x2_ASAP7_75t_R _26844_ (.A(_12905_),
    .B(_01713_),
    .Y(_04460_));
 XOR2x2_ASAP7_75t_R _26845_ (.A(_04460_),
    .B(_12848_),
    .Y(_04461_));
 NOR2x1_ASAP7_75t_R _26846_ (.A(_00574_),
    .B(_00547_),
    .Y(_04462_));
 AO21x1_ASAP7_75t_R _26847_ (.A1(_04461_),
    .A2(_00574_),
    .B(_04462_),
    .Y(_04463_));
 XOR2x2_ASAP7_75t_SL _26848_ (.A(_04463_),
    .B(_00938_),
    .Y(_04464_));
 AOI21x1_ASAP7_75t_SL _26851_ (.A1(_04444_),
    .A2(_04459_),
    .B(_04464_),
    .Y(_04467_));
 XNOR2x2_ASAP7_75t_SL _26852_ (.A(_00938_),
    .B(_04463_),
    .Y(_04468_));
 NAND2x2_ASAP7_75t_SL _26856_ (.A(_04402_),
    .B(_01298_),
    .Y(_04472_));
 NAND2x1p5_ASAP7_75t_L _26857_ (.A(_04430_),
    .B(_04472_),
    .Y(_04473_));
 NOR2x1_ASAP7_75t_SL _26859_ (.A(_04428_),
    .B(_04408_),
    .Y(_04475_));
 OAI21x1_ASAP7_75t_R _26860_ (.A1(_04421_),
    .A2(_04475_),
    .B(_04441_),
    .Y(_04476_));
 AOI21x1_ASAP7_75t_SL _26861_ (.A1(_04421_),
    .A2(_04473_),
    .B(_04476_),
    .Y(_04477_));
 INVx1_ASAP7_75t_SL _26862_ (.A(_01306_),
    .Y(_04478_));
 NAND2x1_ASAP7_75t_SL _26863_ (.A(_04478_),
    .B(_04402_),
    .Y(_04479_));
 INVx1_ASAP7_75t_SL _26864_ (.A(_01299_),
    .Y(_04480_));
 AOI21x1_ASAP7_75t_R _26866_ (.A1(_04480_),
    .A2(_04408_),
    .B(_04433_),
    .Y(_04482_));
 NAND2x1_ASAP7_75t_R _26867_ (.A(_04479_),
    .B(_04482_),
    .Y(_04483_));
 NAND2x1_ASAP7_75t_SL _26868_ (.A(_04480_),
    .B(_04402_),
    .Y(_04484_));
 NOR2x1p5_ASAP7_75t_SL _26869_ (.A(_04429_),
    .B(_04421_),
    .Y(_04485_));
 NAND2x1_ASAP7_75t_L _26870_ (.A(_04484_),
    .B(_04485_),
    .Y(_04486_));
 AOI21x1_ASAP7_75t_SL _26873_ (.A1(_04483_),
    .A2(_04486_),
    .B(_04441_),
    .Y(_04489_));
 NOR2x1_ASAP7_75t_SL _26874_ (.A(_04477_),
    .B(_04489_),
    .Y(_04490_));
 XOR2x2_ASAP7_75t_SL _26875_ (.A(_00700_),
    .B(_00701_),
    .Y(_04491_));
 XOR2x2_ASAP7_75t_R _26876_ (.A(_04491_),
    .B(_00668_),
    .Y(_04492_));
 XNOR2x2_ASAP7_75t_R _26877_ (.A(_12916_),
    .B(_04492_),
    .Y(_04493_));
 NOR2x1_ASAP7_75t_R _26878_ (.A(_00574_),
    .B(_00546_),
    .Y(_04494_));
 AO21x1_ASAP7_75t_SL _26879_ (.A1(_04493_),
    .A2(_00574_),
    .B(_04494_),
    .Y(_04495_));
 XOR2x2_ASAP7_75t_SL _26880_ (.A(_04495_),
    .B(_00939_),
    .Y(_04496_));
 OAI21x1_ASAP7_75t_SL _26882_ (.A1(_04490_),
    .A2(_04468_),
    .B(_04496_),
    .Y(_04498_));
 NOR2x1_ASAP7_75t_SL _26883_ (.A(_04467_),
    .B(_04498_),
    .Y(_04499_));
 NAND2x2_ASAP7_75t_SL _26884_ (.A(_04408_),
    .B(_01298_),
    .Y(_04500_));
 OAI21x1_ASAP7_75t_SL _26886_ (.A1(_04387_),
    .A2(_04425_),
    .B(_04396_),
    .Y(_04502_));
 NAND3x1_ASAP7_75t_SL _26887_ (.A(_04395_),
    .B(_00935_),
    .C(_04388_),
    .Y(_04503_));
 AOI21x1_ASAP7_75t_R _26889_ (.A1(_04502_),
    .A2(_04503_),
    .B(_01303_),
    .Y(_04505_));
 INVx1_ASAP7_75t_R _26890_ (.A(_04505_),
    .Y(_04506_));
 AND3x1_ASAP7_75t_SL _26891_ (.A(_04500_),
    .B(_04421_),
    .C(_04506_),
    .Y(_04507_));
 AOI21x1_ASAP7_75t_SL _26893_ (.A1(_04448_),
    .A2(_04402_),
    .B(_04421_),
    .Y(_04508_));
 NAND2x1_ASAP7_75t_SL _26895_ (.A(_01309_),
    .B(_04408_),
    .Y(_04510_));
 AO21x1_ASAP7_75t_SL _26897_ (.A1(_04508_),
    .A2(_04510_),
    .B(_04456_),
    .Y(_04512_));
 NOR2x1_ASAP7_75t_SL _26898_ (.A(_04507_),
    .B(_04512_),
    .Y(_04513_));
 AOI21x1_ASAP7_75t_SL _26900_ (.A1(_04426_),
    .A2(_04427_),
    .B(_01301_),
    .Y(_04515_));
 INVx1_ASAP7_75t_R _26901_ (.A(_04515_),
    .Y(_04516_));
 AOI21x1_ASAP7_75t_SL _26902_ (.A1(_04516_),
    .A2(_04472_),
    .B(_04433_),
    .Y(_04517_));
 NAND2x1_ASAP7_75t_SL _26903_ (.A(_04431_),
    .B(_04408_),
    .Y(_04518_));
 AO21x1_ASAP7_75t_SL _26904_ (.A1(_04508_),
    .A2(_04518_),
    .B(_04441_),
    .Y(_04519_));
 OAI21x1_ASAP7_75t_SL _26905_ (.A1(_04517_),
    .A2(_04519_),
    .B(_04464_),
    .Y(_04520_));
 INVx2_ASAP7_75t_SL _26906_ (.A(_04496_),
    .Y(_04521_));
 OAI21x1_ASAP7_75t_SL _26908_ (.A1(_04513_),
    .A2(_04520_),
    .B(_04521_),
    .Y(_04523_));
 INVx2_ASAP7_75t_SL _26909_ (.A(_04485_),
    .Y(_04524_));
 INVx1_ASAP7_75t_R _26910_ (.A(_01309_),
    .Y(_04525_));
 NOR2x1_ASAP7_75t_SL _26911_ (.A(_04525_),
    .B(_04408_),
    .Y(_04526_));
 NAND2x1_ASAP7_75t_R _26912_ (.A(_01303_),
    .B(_04402_),
    .Y(_04527_));
 AO21x1_ASAP7_75t_SL _26914_ (.A1(_04445_),
    .A2(_04527_),
    .B(_04433_),
    .Y(_04529_));
 OA21x2_ASAP7_75t_SL _26915_ (.A1(_04524_),
    .A2(_04526_),
    .B(_04529_),
    .Y(_04530_));
 AOI21x1_ASAP7_75t_R _26916_ (.A1(_01304_),
    .A2(_04408_),
    .B(_04421_),
    .Y(_04531_));
 AOI21x1_ASAP7_75t_R _26917_ (.A1(_04448_),
    .A2(_04402_),
    .B(_04433_),
    .Y(_04532_));
 AO21x1_ASAP7_75t_SL _26918_ (.A1(_04531_),
    .A2(_04506_),
    .B(_04532_),
    .Y(_04533_));
 OAI21x1_ASAP7_75t_SL _26919_ (.A1(_04441_),
    .A2(_04533_),
    .B(_04468_),
    .Y(_04534_));
 AOI21x1_ASAP7_75t_SL _26920_ (.A1(_04441_),
    .A2(_04530_),
    .B(_04534_),
    .Y(_04535_));
 XOR2x2_ASAP7_75t_R _26921_ (.A(_12787_),
    .B(_01748_),
    .Y(_04536_));
 INVx1_ASAP7_75t_R _26922_ (.A(_00569_),
    .Y(_04537_));
 XOR2x2_ASAP7_75t_L _26923_ (.A(_04536_),
    .B(_04537_),
    .Y(_04538_));
 NOR2x1_ASAP7_75t_SL _26924_ (.A(_00574_),
    .B(_00545_),
    .Y(_04539_));
 AO21x1_ASAP7_75t_SL _26925_ (.A1(_04538_),
    .A2(_00574_),
    .B(_04539_),
    .Y(_04540_));
 XOR2x2_ASAP7_75t_SL _26926_ (.A(_04540_),
    .B(_00940_),
    .Y(_04541_));
 OAI21x1_ASAP7_75t_SL _26928_ (.A1(_04523_),
    .A2(_04535_),
    .B(_04541_),
    .Y(_04543_));
 AND2x2_ASAP7_75t_SL _26929_ (.A(_01301_),
    .B(_01304_),
    .Y(_04544_));
 NOR2x1_ASAP7_75t_SL _26930_ (.A(_04544_),
    .B(_04408_),
    .Y(_04545_));
 INVx2_ASAP7_75t_SL _26931_ (.A(_01303_),
    .Y(_04546_));
 AOI21x1_ASAP7_75t_SL _26932_ (.A1(_04426_),
    .A2(_04427_),
    .B(_04546_),
    .Y(_04547_));
 OA21x2_ASAP7_75t_SL _26933_ (.A1(_04545_),
    .A2(_04547_),
    .B(_04421_),
    .Y(_04548_));
 NAND2x1_ASAP7_75t_SL _26934_ (.A(_04480_),
    .B(_04408_),
    .Y(_04549_));
 AOI21x1_ASAP7_75t_SL _26936_ (.A1(_04549_),
    .A2(_04508_),
    .B(_04441_),
    .Y(_04551_));
 INVx1_ASAP7_75t_SL _26937_ (.A(_04551_),
    .Y(_04552_));
 NOR2x1_ASAP7_75t_SL _26940_ (.A(_01300_),
    .B(_04408_),
    .Y(_04555_));
 NAND2x1_ASAP7_75t_R _26942_ (.A(_01314_),
    .B(_04433_),
    .Y(_04557_));
 OAI21x1_ASAP7_75t_SL _26943_ (.A1(_04433_),
    .A2(_04555_),
    .B(_04557_),
    .Y(_04558_));
 AOI21x1_ASAP7_75t_SL _26945_ (.A1(_04441_),
    .A2(_04558_),
    .B(_04468_),
    .Y(_04560_));
 OAI21x1_ASAP7_75t_SL _26946_ (.A1(_04548_),
    .A2(_04552_),
    .B(_04560_),
    .Y(_04561_));
 AOI21x1_ASAP7_75t_SL _26948_ (.A1(_04433_),
    .A2(_04515_),
    .B(_04456_),
    .Y(_04563_));
 OAI21x1_ASAP7_75t_SL _26949_ (.A1(_04406_),
    .A2(_04407_),
    .B(_01306_),
    .Y(_04564_));
 OAI21x1_ASAP7_75t_SL _26950_ (.A1(_04397_),
    .A2(_04401_),
    .B(_01303_),
    .Y(_04565_));
 AO21x1_ASAP7_75t_SL _26951_ (.A1(_04564_),
    .A2(_04565_),
    .B(_04433_),
    .Y(_04566_));
 AOI21x1_ASAP7_75t_SL _26953_ (.A1(_04563_),
    .A2(_04566_),
    .B(_04464_),
    .Y(_04568_));
 INVx1_ASAP7_75t_SL _26954_ (.A(_01307_),
    .Y(_04569_));
 OAI21x1_ASAP7_75t_SL _26955_ (.A1(_04406_),
    .A2(_04407_),
    .B(_04569_),
    .Y(_04570_));
 INVx1_ASAP7_75t_R _26956_ (.A(_04570_),
    .Y(_04571_));
 OAI21x1_ASAP7_75t_SL _26957_ (.A1(_04547_),
    .A2(_04571_),
    .B(_04433_),
    .Y(_04572_));
 NAND2x1_ASAP7_75t_SL _26959_ (.A(_04421_),
    .B(_04515_),
    .Y(_04574_));
 NAND3x1_ASAP7_75t_SL _26960_ (.A(_04572_),
    .B(_04456_),
    .C(_04574_),
    .Y(_04575_));
 AOI21x1_ASAP7_75t_SL _26961_ (.A1(_04568_),
    .A2(_04575_),
    .B(_04521_),
    .Y(_04576_));
 AOI21x1_ASAP7_75t_SL _26962_ (.A1(_04561_),
    .A2(_04576_),
    .B(_04541_),
    .Y(_04577_));
 AOI21x1_ASAP7_75t_R _26963_ (.A1(_04426_),
    .A2(_04427_),
    .B(_01307_),
    .Y(_04578_));
 NAND2x1_ASAP7_75t_SL _26965_ (.A(_04421_),
    .B(_04578_),
    .Y(_04580_));
 NAND3x1_ASAP7_75t_SL _26966_ (.A(_04524_),
    .B(_04441_),
    .C(_04580_),
    .Y(_04581_));
 INVx1_ASAP7_75t_SL _26967_ (.A(_01304_),
    .Y(_04582_));
 OAI21x1_ASAP7_75t_SL _26968_ (.A1(_04406_),
    .A2(_04407_),
    .B(_04582_),
    .Y(_04583_));
 INVx2_ASAP7_75t_SL _26969_ (.A(_04583_),
    .Y(_04584_));
 AO21x1_ASAP7_75t_SL _26970_ (.A1(_04584_),
    .A2(_04421_),
    .B(_04468_),
    .Y(_04585_));
 AOI21x1_ASAP7_75t_SL _26971_ (.A1(_04519_),
    .A2(_04581_),
    .B(_04585_),
    .Y(_04586_));
 NOR2x1_ASAP7_75t_SL _26972_ (.A(_04456_),
    .B(_04531_),
    .Y(_04587_));
 AO21x1_ASAP7_75t_SL _26974_ (.A1(_04410_),
    .A2(_04516_),
    .B(_04433_),
    .Y(_04589_));
 NAND2x1_ASAP7_75t_SL _26975_ (.A(_04587_),
    .B(_04589_),
    .Y(_04590_));
 NAND2x1_ASAP7_75t_SL _26976_ (.A(_01300_),
    .B(_04402_),
    .Y(_04591_));
 AOI21x1_ASAP7_75t_SL _26977_ (.A1(_04591_),
    .A2(_04500_),
    .B(_04433_),
    .Y(_04592_));
 INVx1_ASAP7_75t_SL _26978_ (.A(_04592_),
    .Y(_04593_));
 AOI21x1_ASAP7_75t_R _26979_ (.A1(_04448_),
    .A2(_04408_),
    .B(_04421_),
    .Y(_04594_));
 AOI21x1_ASAP7_75t_SL _26980_ (.A1(_04479_),
    .A2(_04594_),
    .B(_04441_),
    .Y(_04595_));
 NAND2x1_ASAP7_75t_SL _26981_ (.A(_04593_),
    .B(_04595_),
    .Y(_04596_));
 AOI21x1_ASAP7_75t_SL _26982_ (.A1(_04590_),
    .A2(_04596_),
    .B(_04464_),
    .Y(_04597_));
 OAI21x1_ASAP7_75t_SL _26983_ (.A1(_04586_),
    .A2(_04597_),
    .B(_04521_),
    .Y(_04598_));
 NAND2x1_ASAP7_75t_SL _26984_ (.A(_04577_),
    .B(_04598_),
    .Y(_04599_));
 OAI21x1_ASAP7_75t_SL _26985_ (.A1(_04499_),
    .A2(_04543_),
    .B(_04599_),
    .Y(_00120_));
 NAND2x1_ASAP7_75t_SL _26986_ (.A(_04430_),
    .B(_04508_),
    .Y(_04600_));
 NAND2x1_ASAP7_75t_SL _26987_ (.A(_01305_),
    .B(_04402_),
    .Y(_04601_));
 AOI21x1_ASAP7_75t_SL _26988_ (.A1(_01304_),
    .A2(_04408_),
    .B(_04433_),
    .Y(_04602_));
 AOI21x1_ASAP7_75t_SL _26989_ (.A1(_04601_),
    .A2(_04602_),
    .B(_04456_),
    .Y(_04603_));
 NAND2x1_ASAP7_75t_SL _26990_ (.A(_04600_),
    .B(_04603_),
    .Y(_04604_));
 NOR2x1_ASAP7_75t_SL _26991_ (.A(_04421_),
    .B(_04408_),
    .Y(_04605_));
 AOI21x1_ASAP7_75t_SL _26992_ (.A1(_01303_),
    .A2(_04605_),
    .B(_04441_),
    .Y(_04606_));
 AOI21x1_ASAP7_75t_R _26993_ (.A1(_04408_),
    .A2(_01302_),
    .B(_04433_),
    .Y(_04607_));
 NAND2x1_ASAP7_75t_SL _26994_ (.A(_04449_),
    .B(_04607_),
    .Y(_04608_));
 AOI21x1_ASAP7_75t_SL _26995_ (.A1(_04606_),
    .A2(_04608_),
    .B(_04464_),
    .Y(_04609_));
 AOI21x1_ASAP7_75t_SL _26996_ (.A1(_04604_),
    .A2(_04609_),
    .B(_04521_),
    .Y(_04610_));
 NOR2x1_ASAP7_75t_R _26997_ (.A(_04433_),
    .B(_04565_),
    .Y(_04611_));
 OAI21x1_ASAP7_75t_R _26998_ (.A1(_04433_),
    .A2(_04583_),
    .B(_04456_),
    .Y(_04612_));
 NOR2x1_ASAP7_75t_SL _26999_ (.A(_04611_),
    .B(_04612_),
    .Y(_04613_));
 NOR2x1p5_ASAP7_75t_SL _27000_ (.A(_04421_),
    .B(_04475_),
    .Y(_04614_));
 NAND2x1_ASAP7_75t_SL _27001_ (.A(_04510_),
    .B(_04614_),
    .Y(_04615_));
 NAND2x1_ASAP7_75t_SL _27002_ (.A(_04613_),
    .B(_04615_),
    .Y(_04616_));
 OA21x2_ASAP7_75t_SL _27003_ (.A1(_04583_),
    .A2(_04433_),
    .B(_04441_),
    .Y(_04617_));
 NAND2x1_ASAP7_75t_R _27004_ (.A(_01318_),
    .B(_04433_),
    .Y(_04618_));
 OA21x2_ASAP7_75t_SL _27005_ (.A1(_04500_),
    .A2(_04433_),
    .B(_04618_),
    .Y(_04619_));
 AOI21x1_ASAP7_75t_SL _27006_ (.A1(_04617_),
    .A2(_04619_),
    .B(_04468_),
    .Y(_04620_));
 NAND2x1_ASAP7_75t_SL _27007_ (.A(_04616_),
    .B(_04620_),
    .Y(_04621_));
 AOI21x1_ASAP7_75t_SL _27008_ (.A1(_04610_),
    .A2(_04621_),
    .B(_04541_),
    .Y(_04622_));
 AOI21x1_ASAP7_75t_SL _27009_ (.A1(_04426_),
    .A2(_04427_),
    .B(_01300_),
    .Y(_04623_));
 INVx2_ASAP7_75t_SL _27010_ (.A(_04623_),
    .Y(_04624_));
 AOI21x1_ASAP7_75t_SL _27011_ (.A1(_04431_),
    .A2(_04402_),
    .B(_04421_),
    .Y(_04625_));
 NAND2x1_ASAP7_75t_SL _27012_ (.A(_04624_),
    .B(_04625_),
    .Y(_04626_));
 NAND2x1_ASAP7_75t_R _27013_ (.A(_04582_),
    .B(_04421_),
    .Y(_04627_));
 OA21x2_ASAP7_75t_SL _27014_ (.A1(_04627_),
    .A2(_04402_),
    .B(_04456_),
    .Y(_04628_));
 AOI21x1_ASAP7_75t_SL _27015_ (.A1(_04626_),
    .A2(_04628_),
    .B(_04464_),
    .Y(_04629_));
 AOI21x1_ASAP7_75t_R _27016_ (.A1(_04426_),
    .A2(_04427_),
    .B(_04431_),
    .Y(_04630_));
 NAND2x1_ASAP7_75t_SL _27017_ (.A(_04421_),
    .B(_04630_),
    .Y(_04631_));
 NOR2x1_ASAP7_75t_R _27018_ (.A(_04421_),
    .B(_04526_),
    .Y(_04632_));
 AOI21x1_ASAP7_75t_SL _27019_ (.A1(_04500_),
    .A2(_04632_),
    .B(_04456_),
    .Y(_04633_));
 NAND2x1_ASAP7_75t_SL _27020_ (.A(_04631_),
    .B(_04633_),
    .Y(_04634_));
 AOI21x1_ASAP7_75t_SL _27021_ (.A1(_04629_),
    .A2(_04634_),
    .B(_04496_),
    .Y(_04635_));
 AO21x1_ASAP7_75t_SL _27022_ (.A1(_04583_),
    .A2(_04430_),
    .B(_04421_),
    .Y(_04636_));
 AOI21x1_ASAP7_75t_R _27023_ (.A1(_04426_),
    .A2(_04427_),
    .B(_04480_),
    .Y(_04637_));
 INVx1_ASAP7_75t_R _27024_ (.A(_04637_),
    .Y(_04638_));
 AO21x1_ASAP7_75t_SL _27025_ (.A1(_04601_),
    .A2(_04638_),
    .B(_04433_),
    .Y(_04639_));
 AOI21x1_ASAP7_75t_SL _27026_ (.A1(_04636_),
    .A2(_04639_),
    .B(_04456_),
    .Y(_04640_));
 AO21x1_ASAP7_75t_SL _27027_ (.A1(_04445_),
    .A2(_04591_),
    .B(_04433_),
    .Y(_04641_));
 NAND2x1_ASAP7_75t_R _27028_ (.A(_01305_),
    .B(_01302_),
    .Y(_04642_));
 NAND2x2_ASAP7_75t_SL _27029_ (.A(_04448_),
    .B(_04408_),
    .Y(_04643_));
 AO21x1_ASAP7_75t_SL _27030_ (.A1(_04642_),
    .A2(_04643_),
    .B(_04421_),
    .Y(_04644_));
 AOI21x1_ASAP7_75t_SL _27031_ (.A1(_04641_),
    .A2(_04644_),
    .B(_04441_),
    .Y(_04645_));
 OAI21x1_ASAP7_75t_SL _27032_ (.A1(_04640_),
    .A2(_04645_),
    .B(_04464_),
    .Y(_04646_));
 NAND2x1_ASAP7_75t_SL _27033_ (.A(_04635_),
    .B(_04646_),
    .Y(_04647_));
 NAND2x1_ASAP7_75t_SL _27034_ (.A(_04622_),
    .B(_04647_),
    .Y(_04648_));
 NOR2x1_ASAP7_75t_SL _27035_ (.A(_04408_),
    .B(_01298_),
    .Y(_04649_));
 OAI21x1_ASAP7_75t_SL _27036_ (.A1(_04448_),
    .A2(_04402_),
    .B(_04421_),
    .Y(_04650_));
 NOR2x1_ASAP7_75t_SL _27037_ (.A(_04649_),
    .B(_04650_),
    .Y(_04651_));
 AOI211x1_ASAP7_75t_SL _27038_ (.A1(_04472_),
    .A2(_04531_),
    .B(_04651_),
    .C(_04468_),
    .Y(_04652_));
 AOI21x1_ASAP7_75t_SL _27040_ (.A1(_04410_),
    .A2(_04445_),
    .B(_04433_),
    .Y(_04654_));
 NOR2x1_ASAP7_75t_SL _27041_ (.A(_04421_),
    .B(_04505_),
    .Y(_04655_));
 AO21x1_ASAP7_75t_SL _27042_ (.A1(_04655_),
    .A2(_04518_),
    .B(_04464_),
    .Y(_04656_));
 OAI21x1_ASAP7_75t_SL _27043_ (.A1(_04654_),
    .A2(_04656_),
    .B(_04441_),
    .Y(_04657_));
 INVx1_ASAP7_75t_SL _27044_ (.A(_01316_),
    .Y(_04658_));
 NOR2x1_ASAP7_75t_R _27045_ (.A(_04421_),
    .B(_04468_),
    .Y(_04659_));
 INVx1_ASAP7_75t_SL _27046_ (.A(_04659_),
    .Y(_04660_));
 INVx1_ASAP7_75t_SL _27047_ (.A(_04564_),
    .Y(_04661_));
 OAI21x1_ASAP7_75t_SL _27048_ (.A1(_04630_),
    .A2(_04661_),
    .B(_04421_),
    .Y(_04662_));
 OAI21x1_ASAP7_75t_SL _27049_ (.A1(_04658_),
    .A2(_04660_),
    .B(_04662_),
    .Y(_04663_));
 AOI21x1_ASAP7_75t_SL _27050_ (.A1(_04456_),
    .A2(_04663_),
    .B(_04521_),
    .Y(_04664_));
 OAI21x1_ASAP7_75t_SL _27051_ (.A1(_04652_),
    .A2(_04657_),
    .B(_04664_),
    .Y(_04665_));
 OAI21x1_ASAP7_75t_SL _27052_ (.A1(_04433_),
    .A2(_04601_),
    .B(_04441_),
    .Y(_04666_));
 INVx1_ASAP7_75t_SL _27053_ (.A(_04574_),
    .Y(_04667_));
 AO21x1_ASAP7_75t_SL _27054_ (.A1(_04614_),
    .A2(_04549_),
    .B(_04667_),
    .Y(_04668_));
 NAND2x1_ASAP7_75t_SL _27055_ (.A(_04472_),
    .B(_04531_),
    .Y(_04669_));
 AOI21x1_ASAP7_75t_SL _27056_ (.A1(_04484_),
    .A2(_04454_),
    .B(_04441_),
    .Y(_04670_));
 AOI21x1_ASAP7_75t_SL _27057_ (.A1(_04669_),
    .A2(_04670_),
    .B(_04464_),
    .Y(_04671_));
 OAI21x1_ASAP7_75t_SL _27058_ (.A1(_04666_),
    .A2(_04668_),
    .B(_04671_),
    .Y(_04672_));
 NAND2x1_ASAP7_75t_SL _27059_ (.A(_04518_),
    .B(_04532_),
    .Y(_04673_));
 NOR2x1_ASAP7_75t_SL _27060_ (.A(_04441_),
    .B(_04485_),
    .Y(_04674_));
 AOI21x1_ASAP7_75t_SL _27061_ (.A1(_04673_),
    .A2(_04674_),
    .B(_04468_),
    .Y(_04675_));
 AOI21x1_ASAP7_75t_SL _27062_ (.A1(_01301_),
    .A2(_04402_),
    .B(_04433_),
    .Y(_04676_));
 NAND2x1_ASAP7_75t_SL _27063_ (.A(_04510_),
    .B(_04676_),
    .Y(_04677_));
 NAND3x1_ASAP7_75t_SL _27064_ (.A(_04626_),
    .B(_04677_),
    .C(_04441_),
    .Y(_04678_));
 AOI21x1_ASAP7_75t_SL _27065_ (.A1(_04675_),
    .A2(_04678_),
    .B(_04496_),
    .Y(_04679_));
 INVx1_ASAP7_75t_SL _27066_ (.A(_04541_),
    .Y(_04680_));
 AOI21x1_ASAP7_75t_SL _27067_ (.A1(_04672_),
    .A2(_04679_),
    .B(_04680_),
    .Y(_04681_));
 NAND2x1_ASAP7_75t_SL _27068_ (.A(_04665_),
    .B(_04681_),
    .Y(_04682_));
 NAND2x1_ASAP7_75t_SL _27069_ (.A(_04648_),
    .B(_04682_),
    .Y(_00121_));
 NAND2x1_ASAP7_75t_SL _27070_ (.A(_04472_),
    .B(_04594_),
    .Y(_04683_));
 AO21x1_ASAP7_75t_SL _27071_ (.A1(_04593_),
    .A2(_04683_),
    .B(_04456_),
    .Y(_04684_));
 NAND2x1_ASAP7_75t_SL _27072_ (.A(_04546_),
    .B(_04408_),
    .Y(_04685_));
 NOR2x1_ASAP7_75t_SL _27073_ (.A(_01314_),
    .B(_04433_),
    .Y(_04686_));
 AO21x1_ASAP7_75t_SL _27074_ (.A1(_04614_),
    .A2(_04685_),
    .B(_04686_),
    .Y(_04687_));
 NAND2x1_ASAP7_75t_SL _27075_ (.A(_04456_),
    .B(_04687_),
    .Y(_04688_));
 AOI21x1_ASAP7_75t_SL _27076_ (.A1(_04684_),
    .A2(_04688_),
    .B(_04464_),
    .Y(_04689_));
 AOI21x1_ASAP7_75t_R _27077_ (.A1(_04408_),
    .A2(_01302_),
    .B(_04421_),
    .Y(_04690_));
 AOI21x1_ASAP7_75t_SL _27078_ (.A1(_04449_),
    .A2(_04690_),
    .B(_04441_),
    .Y(_04691_));
 NAND2x1_ASAP7_75t_SL _27079_ (.A(_01316_),
    .B(_04421_),
    .Y(_04692_));
 AO21x1_ASAP7_75t_SL _27080_ (.A1(_04691_),
    .A2(_04692_),
    .B(_04468_),
    .Y(_04693_));
 NAND2x1_ASAP7_75t_R _27081_ (.A(_04408_),
    .B(_01302_),
    .Y(_04694_));
 AO21x1_ASAP7_75t_SL _27082_ (.A1(_04694_),
    .A2(_04410_),
    .B(_04433_),
    .Y(_04695_));
 NAND2x1p5_ASAP7_75t_SL _27083_ (.A(_04428_),
    .B(_04402_),
    .Y(_04696_));
 AO21x1_ASAP7_75t_SL _27084_ (.A1(_04412_),
    .A2(_04696_),
    .B(_04421_),
    .Y(_04697_));
 AND3x1_ASAP7_75t_SL _27085_ (.A(_04695_),
    .B(_04441_),
    .C(_04697_),
    .Y(_04698_));
 OAI21x1_ASAP7_75t_SL _27086_ (.A1(_04693_),
    .A2(_04698_),
    .B(_04680_),
    .Y(_04699_));
 NOR2x1_ASAP7_75t_SL _27087_ (.A(_04689_),
    .B(_04699_),
    .Y(_04700_));
 OAI21x1_ASAP7_75t_SL _27088_ (.A1(_04578_),
    .A2(_04584_),
    .B(_04421_),
    .Y(_04701_));
 AOI21x1_ASAP7_75t_SL _27089_ (.A1(_01304_),
    .A2(_04402_),
    .B(_04421_),
    .Y(_04702_));
 NAND2x1_ASAP7_75t_SL _27090_ (.A(_04500_),
    .B(_04702_),
    .Y(_04703_));
 AOI21x1_ASAP7_75t_SL _27091_ (.A1(_04701_),
    .A2(_04703_),
    .B(_04441_),
    .Y(_04704_));
 AOI21x1_ASAP7_75t_SL _27092_ (.A1(_04502_),
    .A2(_04503_),
    .B(_01309_),
    .Y(_04705_));
 OAI21x1_ASAP7_75t_SL _27093_ (.A1(_04578_),
    .A2(_04705_),
    .B(_04421_),
    .Y(_04706_));
 NAND2x1_ASAP7_75t_SL _27094_ (.A(_04643_),
    .B(_04702_),
    .Y(_04707_));
 AOI21x1_ASAP7_75t_SL _27095_ (.A1(_04706_),
    .A2(_04707_),
    .B(_04456_),
    .Y(_04708_));
 OAI21x1_ASAP7_75t_SL _27096_ (.A1(_04704_),
    .A2(_04708_),
    .B(_04464_),
    .Y(_04709_));
 AOI21x1_ASAP7_75t_SL _27097_ (.A1(_01307_),
    .A2(_04402_),
    .B(_04433_),
    .Y(_04710_));
 NAND2x1_ASAP7_75t_SL _27098_ (.A(_04643_),
    .B(_04710_),
    .Y(_04711_));
 OAI21x1_ASAP7_75t_SL _27099_ (.A1(_04623_),
    .A2(_04475_),
    .B(_04433_),
    .Y(_04712_));
 AOI21x1_ASAP7_75t_SL _27100_ (.A1(_04711_),
    .A2(_04712_),
    .B(_04441_),
    .Y(_04713_));
 AOI211x1_ASAP7_75t_SL _27101_ (.A1(_01298_),
    .A2(_04402_),
    .B(_04578_),
    .C(_04421_),
    .Y(_04714_));
 OAI21x1_ASAP7_75t_SL _27102_ (.A1(_04705_),
    .A2(_04650_),
    .B(_04441_),
    .Y(_04715_));
 NOR2x1_ASAP7_75t_SL _27103_ (.A(_04714_),
    .B(_04715_),
    .Y(_04716_));
 OAI21x1_ASAP7_75t_SL _27104_ (.A1(_04713_),
    .A2(_04716_),
    .B(_04468_),
    .Y(_04717_));
 NAND2x1_ASAP7_75t_SL _27105_ (.A(_04709_),
    .B(_04717_),
    .Y(_04718_));
 OAI21x1_ASAP7_75t_SL _27106_ (.A1(_04680_),
    .A2(_04718_),
    .B(_04521_),
    .Y(_04719_));
 NAND2x1_ASAP7_75t_SL _27107_ (.A(_01309_),
    .B(_04402_),
    .Y(_04720_));
 NAND2x1_ASAP7_75t_SL _27108_ (.A(_04720_),
    .B(_04602_),
    .Y(_04721_));
 NAND2x1_ASAP7_75t_SL _27109_ (.A(_04694_),
    .B(_04655_),
    .Y(_04722_));
 AOI21x1_ASAP7_75t_SL _27110_ (.A1(_04721_),
    .A2(_04722_),
    .B(_04456_),
    .Y(_04723_));
 NAND2x1_ASAP7_75t_SL _27111_ (.A(_04433_),
    .B(_04565_),
    .Y(_04724_));
 OAI21x1_ASAP7_75t_SL _27112_ (.A1(_04584_),
    .A2(_04724_),
    .B(_04456_),
    .Y(_04725_));
 OAI21x1_ASAP7_75t_SL _27113_ (.A1(_04592_),
    .A2(_04725_),
    .B(_04464_),
    .Y(_04726_));
 NOR2x1_ASAP7_75t_SL _27114_ (.A(_04723_),
    .B(_04726_),
    .Y(_04727_));
 AO21x1_ASAP7_75t_SL _27115_ (.A1(_04402_),
    .A2(_04546_),
    .B(_04433_),
    .Y(_04728_));
 NAND2x1_ASAP7_75t_SL _27116_ (.A(_04510_),
    .B(_04625_),
    .Y(_04729_));
 AOI21x1_ASAP7_75t_SL _27117_ (.A1(_04728_),
    .A2(_04729_),
    .B(_04441_),
    .Y(_04730_));
 NOR2x1_ASAP7_75t_SL _27118_ (.A(_01301_),
    .B(_04408_),
    .Y(_04731_));
 OAI21x1_ASAP7_75t_SL _27119_ (.A1(_04448_),
    .A2(_04402_),
    .B(_04433_),
    .Y(_04732_));
 NOR2x1_ASAP7_75t_SL _27120_ (.A(_04731_),
    .B(_04732_),
    .Y(_04733_));
 OAI21x1_ASAP7_75t_SL _27121_ (.A1(_04408_),
    .A2(_01302_),
    .B(_04421_),
    .Y(_04734_));
 OAI21x1_ASAP7_75t_SL _27122_ (.A1(_04623_),
    .A2(_04734_),
    .B(_04441_),
    .Y(_04735_));
 OAI21x1_ASAP7_75t_SL _27123_ (.A1(_04733_),
    .A2(_04735_),
    .B(_04468_),
    .Y(_04736_));
 NOR2x1_ASAP7_75t_SL _27124_ (.A(_04730_),
    .B(_04736_),
    .Y(_04737_));
 OAI21x1_ASAP7_75t_SL _27125_ (.A1(_04727_),
    .A2(_04737_),
    .B(_04541_),
    .Y(_04738_));
 NAND2x1_ASAP7_75t_SL _27126_ (.A(_04421_),
    .B(_04637_),
    .Y(_04739_));
 OAI21x1_ASAP7_75t_SL _27127_ (.A1(_04623_),
    .A2(_04584_),
    .B(_04433_),
    .Y(_04740_));
 AOI21x1_ASAP7_75t_SL _27128_ (.A1(_04739_),
    .A2(_04740_),
    .B(_04441_),
    .Y(_04741_));
 NAND2x1_ASAP7_75t_R _27129_ (.A(_04544_),
    .B(_04408_),
    .Y(_04742_));
 NAND2x1_ASAP7_75t_SL _27130_ (.A(_04742_),
    .B(_04625_),
    .Y(_04743_));
 AOI21x1_ASAP7_75t_SL _27131_ (.A1(_04662_),
    .A2(_04743_),
    .B(_04456_),
    .Y(_04744_));
 OAI21x1_ASAP7_75t_SL _27132_ (.A1(_04741_),
    .A2(_04744_),
    .B(_04468_),
    .Y(_04745_));
 NAND2x1_ASAP7_75t_SL _27133_ (.A(_01313_),
    .B(_04433_),
    .Y(_04746_));
 OAI21x1_ASAP7_75t_SL _27134_ (.A1(_04433_),
    .A2(_04505_),
    .B(_04746_),
    .Y(_04747_));
 OR2x2_ASAP7_75t_SL _27135_ (.A(_04747_),
    .B(_04441_),
    .Y(_04748_));
 OA21x2_ASAP7_75t_SL _27136_ (.A1(_01319_),
    .A2(_04433_),
    .B(_04441_),
    .Y(_04749_));
 AOI21x1_ASAP7_75t_SL _27137_ (.A1(_04749_),
    .A2(_04722_),
    .B(_04468_),
    .Y(_04750_));
 AOI21x1_ASAP7_75t_SL _27138_ (.A1(_04748_),
    .A2(_04750_),
    .B(_04541_),
    .Y(_04751_));
 AOI21x1_ASAP7_75t_SL _27139_ (.A1(_04745_),
    .A2(_04751_),
    .B(_04521_),
    .Y(_04752_));
 NAND2x1_ASAP7_75t_SL _27140_ (.A(_04738_),
    .B(_04752_),
    .Y(_04753_));
 OAI21x1_ASAP7_75t_SL _27141_ (.A1(_04700_),
    .A2(_04719_),
    .B(_04753_),
    .Y(_00122_));
 AND2x2_ASAP7_75t_SL _27142_ (.A(_04710_),
    .B(_04624_),
    .Y(_04754_));
 NOR2x1_ASAP7_75t_R _27143_ (.A(_04402_),
    .B(_01302_),
    .Y(_04755_));
 AO21x1_ASAP7_75t_SL _27144_ (.A1(_04402_),
    .A2(_01309_),
    .B(_04421_),
    .Y(_04756_));
 OAI21x1_ASAP7_75t_SL _27145_ (.A1(_04755_),
    .A2(_04756_),
    .B(_04441_),
    .Y(_04757_));
 OAI21x1_ASAP7_75t_SL _27146_ (.A1(_04754_),
    .A2(_04757_),
    .B(_04521_),
    .Y(_04758_));
 AND2x2_ASAP7_75t_SL _27147_ (.A(_04449_),
    .B(_04601_),
    .Y(_04759_));
 OAI21x1_ASAP7_75t_SL _27148_ (.A1(_04433_),
    .A2(_04759_),
    .B(_04456_),
    .Y(_04760_));
 NOR2x1_ASAP7_75t_SL _27149_ (.A(_04655_),
    .B(_04760_),
    .Y(_04761_));
 NOR2x1_ASAP7_75t_SL _27150_ (.A(_04758_),
    .B(_04761_),
    .Y(_04762_));
 AND3x1_ASAP7_75t_SL _27151_ (.A(_04472_),
    .B(_04643_),
    .C(_04421_),
    .Y(_04763_));
 OAI21x1_ASAP7_75t_SL _27152_ (.A1(_04476_),
    .A2(_04763_),
    .B(_04496_),
    .Y(_04764_));
 NOR2x1_ASAP7_75t_SL _27153_ (.A(_04421_),
    .B(_04473_),
    .Y(_04765_));
 NOR2x1_ASAP7_75t_SL _27154_ (.A(_04765_),
    .B(_04760_),
    .Y(_04766_));
 OAI21x1_ASAP7_75t_SL _27155_ (.A1(_04766_),
    .A2(_04764_),
    .B(_04464_),
    .Y(_04767_));
 OAI21x1_ASAP7_75t_SL _27156_ (.A1(_04762_),
    .A2(_04767_),
    .B(_04680_),
    .Y(_04768_));
 OAI21x1_ASAP7_75t_SL _27157_ (.A1(_04623_),
    .A2(_04734_),
    .B(_04456_),
    .Y(_04769_));
 AOI21x1_ASAP7_75t_SL _27158_ (.A1(_04510_),
    .A2(_04702_),
    .B(_04769_),
    .Y(_04770_));
 NAND2x1_ASAP7_75t_SL _27159_ (.A(_04638_),
    .B(_04614_),
    .Y(_04771_));
 AND2x2_ASAP7_75t_SL _27160_ (.A(_04601_),
    .B(_04421_),
    .Y(_04772_));
 NAND2x1_ASAP7_75t_SL _27161_ (.A(_04412_),
    .B(_04772_),
    .Y(_04773_));
 AOI21x1_ASAP7_75t_SL _27162_ (.A1(_04771_),
    .A2(_04773_),
    .B(_04456_),
    .Y(_04774_));
 OAI21x1_ASAP7_75t_SL _27163_ (.A1(_04770_),
    .A2(_04774_),
    .B(_04496_),
    .Y(_04775_));
 OR3x1_ASAP7_75t_SL _27164_ (.A(_04661_),
    .B(_04433_),
    .C(_04429_),
    .Y(_04776_));
 NOR2x1_ASAP7_75t_SL _27165_ (.A(_04456_),
    .B(_04451_),
    .Y(_04777_));
 NAND2x1_ASAP7_75t_SL _27166_ (.A(_04776_),
    .B(_04777_),
    .Y(_04778_));
 INVx1_ASAP7_75t_SL _27167_ (.A(_04630_),
    .Y(_04779_));
 AOI21x1_ASAP7_75t_SL _27168_ (.A1(_04779_),
    .A2(_04696_),
    .B(_04433_),
    .Y(_04780_));
 AOI21x1_ASAP7_75t_SL _27169_ (.A1(_04412_),
    .A2(_04527_),
    .B(_04421_),
    .Y(_04781_));
 OAI21x1_ASAP7_75t_SL _27170_ (.A1(_04780_),
    .A2(_04781_),
    .B(_04456_),
    .Y(_04782_));
 NAND3x1_ASAP7_75t_SL _27171_ (.A(_04778_),
    .B(_04521_),
    .C(_04782_),
    .Y(_04783_));
 AOI21x1_ASAP7_75t_SL _27172_ (.A1(_04775_),
    .A2(_04783_),
    .B(_04464_),
    .Y(_04784_));
 OAI21x1_ASAP7_75t_SL _27173_ (.A1(_04591_),
    .A2(_04660_),
    .B(_04563_),
    .Y(_04785_));
 AO21x1_ASAP7_75t_SL _27174_ (.A1(_04402_),
    .A2(_04478_),
    .B(_04433_),
    .Y(_04786_));
 NAND2x1_ASAP7_75t_SL _27175_ (.A(_04464_),
    .B(_04694_),
    .Y(_04787_));
 NAND3x1_ASAP7_75t_SL _27176_ (.A(_04429_),
    .B(_04468_),
    .C(_04421_),
    .Y(_04788_));
 OAI21x1_ASAP7_75t_SL _27177_ (.A1(_04786_),
    .A2(_04787_),
    .B(_04788_),
    .Y(_04789_));
 OAI21x1_ASAP7_75t_SL _27178_ (.A1(_04785_),
    .A2(_04789_),
    .B(_04496_),
    .Y(_04790_));
 AOI21x1_ASAP7_75t_SL _27179_ (.A1(_04433_),
    .A2(_04578_),
    .B(_04464_),
    .Y(_04791_));
 NAND2x1_ASAP7_75t_SL _27180_ (.A(_04791_),
    .B(_04711_),
    .Y(_04792_));
 NAND2x1p5_ASAP7_75t_SL _27181_ (.A(_04430_),
    .B(_04532_),
    .Y(_04793_));
 AOI21x1_ASAP7_75t_SL _27182_ (.A1(_04544_),
    .A2(_04408_),
    .B(_04421_),
    .Y(_04794_));
 AOI21x1_ASAP7_75t_SL _27183_ (.A1(_04720_),
    .A2(_04794_),
    .B(_04468_),
    .Y(_04795_));
 NAND2x1_ASAP7_75t_SL _27184_ (.A(_04793_),
    .B(_04795_),
    .Y(_04796_));
 AOI21x1_ASAP7_75t_SL _27185_ (.A1(_04792_),
    .A2(_04796_),
    .B(_04441_),
    .Y(_04797_));
 NOR2x1_ASAP7_75t_SL _27186_ (.A(_04790_),
    .B(_04797_),
    .Y(_04798_));
 AOI21x1_ASAP7_75t_R _27187_ (.A1(_01307_),
    .A2(_04402_),
    .B(_04421_),
    .Y(_04799_));
 NAND2x1_ASAP7_75t_SL _27188_ (.A(_04742_),
    .B(_04799_),
    .Y(_04800_));
 AOI21x1_ASAP7_75t_SL _27189_ (.A1(_04662_),
    .A2(_04800_),
    .B(_04441_),
    .Y(_04801_));
 NAND2x1_ASAP7_75t_SL _27190_ (.A(_04464_),
    .B(_04715_),
    .Y(_04802_));
 OAI21x1_ASAP7_75t_SL _27191_ (.A1(_04801_),
    .A2(_04802_),
    .B(_04521_),
    .Y(_04803_));
 NAND2x1_ASAP7_75t_SL _27192_ (.A(_04608_),
    .B(_04551_),
    .Y(_04804_));
 OAI21x1_ASAP7_75t_SL _27193_ (.A1(_04623_),
    .A2(_04705_),
    .B(_04421_),
    .Y(_04805_));
 NAND2x1_ASAP7_75t_SL _27194_ (.A(_04448_),
    .B(_04605_),
    .Y(_04806_));
 AOI21x1_ASAP7_75t_SL _27195_ (.A1(_04433_),
    .A2(_04578_),
    .B(_04456_),
    .Y(_04807_));
 NAND3x1_ASAP7_75t_SL _27196_ (.A(_04805_),
    .B(_04806_),
    .C(_04807_),
    .Y(_04808_));
 AOI21x1_ASAP7_75t_SL _27197_ (.A1(_04804_),
    .A2(_04808_),
    .B(_04464_),
    .Y(_04809_));
 NOR2x1_ASAP7_75t_SL _27198_ (.A(_04803_),
    .B(_04809_),
    .Y(_04810_));
 OAI21x1_ASAP7_75t_SL _27199_ (.A1(_04798_),
    .A2(_04810_),
    .B(_04541_),
    .Y(_04811_));
 OAI21x1_ASAP7_75t_SL _27200_ (.A1(_04768_),
    .A2(_04784_),
    .B(_04811_),
    .Y(_00123_));
 NAND2x1_ASAP7_75t_R _27201_ (.A(_04410_),
    .B(_04690_),
    .Y(_04812_));
 AO21x1_ASAP7_75t_R _27202_ (.A1(_04500_),
    .A2(_04642_),
    .B(_04433_),
    .Y(_04813_));
 AOI21x1_ASAP7_75t_R _27203_ (.A1(_04812_),
    .A2(_04813_),
    .B(_04456_),
    .Y(_04814_));
 INVx1_ASAP7_75t_R _27204_ (.A(_04691_),
    .Y(_04815_));
 OAI21x1_ASAP7_75t_R _27205_ (.A1(_04651_),
    .A2(_04815_),
    .B(_04464_),
    .Y(_04816_));
 NOR2x1_ASAP7_75t_SL _27206_ (.A(_04814_),
    .B(_04816_),
    .Y(_04817_));
 OAI21x1_ASAP7_75t_R _27207_ (.A1(_04515_),
    .A2(_04799_),
    .B(_04441_),
    .Y(_04818_));
 AOI21x1_ASAP7_75t_SL _27208_ (.A1(_04445_),
    .A2(_04472_),
    .B(_04421_),
    .Y(_04819_));
 OAI21x1_ASAP7_75t_R _27209_ (.A1(_04654_),
    .A2(_04819_),
    .B(_04456_),
    .Y(_04820_));
 AOI21x1_ASAP7_75t_R _27210_ (.A1(_04818_),
    .A2(_04820_),
    .B(_04464_),
    .Y(_04821_));
 NOR3x1_ASAP7_75t_SL _27211_ (.A(_04817_),
    .B(_04496_),
    .C(_04821_),
    .Y(_04822_));
 OAI21x1_ASAP7_75t_R _27212_ (.A1(_04637_),
    .A2(_04649_),
    .B(_04433_),
    .Y(_04823_));
 AOI21x1_ASAP7_75t_SL _27213_ (.A1(_04823_),
    .A2(_04613_),
    .B(_04468_),
    .Y(_04824_));
 AOI21x1_ASAP7_75t_R _27214_ (.A1(_04546_),
    .A2(_04408_),
    .B(_04421_),
    .Y(_04825_));
 NAND2x1_ASAP7_75t_R _27215_ (.A(_04472_),
    .B(_04825_),
    .Y(_04826_));
 NAND3x1_ASAP7_75t_R _27216_ (.A(_04721_),
    .B(_04826_),
    .C(_04441_),
    .Y(_04827_));
 NAND2x1_ASAP7_75t_SL _27217_ (.A(_04824_),
    .B(_04827_),
    .Y(_04828_));
 AOI21x1_ASAP7_75t_SL _27218_ (.A1(_01309_),
    .A2(_04408_),
    .B(_04433_),
    .Y(_04829_));
 NAND2x1_ASAP7_75t_L _27219_ (.A(_04591_),
    .B(_04829_),
    .Y(_04830_));
 AOI21x1_ASAP7_75t_R _27220_ (.A1(_04572_),
    .A2(_04830_),
    .B(_04441_),
    .Y(_04831_));
 OAI21x1_ASAP7_75t_R _27221_ (.A1(_04578_),
    .A2(_04555_),
    .B(_04433_),
    .Y(_04832_));
 AOI21x1_ASAP7_75t_R _27222_ (.A1(_04701_),
    .A2(_04832_),
    .B(_04456_),
    .Y(_04833_));
 OAI21x1_ASAP7_75t_R _27223_ (.A1(_04831_),
    .A2(_04833_),
    .B(_04468_),
    .Y(_04834_));
 NAND2x1_ASAP7_75t_SL _27224_ (.A(_04828_),
    .B(_04834_),
    .Y(_04835_));
 OAI21x1_ASAP7_75t_R _27225_ (.A1(_04521_),
    .A2(_04835_),
    .B(_04680_),
    .Y(_04836_));
 AND2x2_ASAP7_75t_R _27226_ (.A(_04799_),
    .B(_04445_),
    .Y(_04837_));
 NOR2x1_ASAP7_75t_R _27227_ (.A(_04448_),
    .B(_01298_),
    .Y(_04838_));
 OA21x2_ASAP7_75t_SL _27228_ (.A1(_04755_),
    .A2(_04838_),
    .B(_04421_),
    .Y(_04839_));
 OAI21x1_ASAP7_75t_R _27229_ (.A1(_04837_),
    .A2(_04839_),
    .B(_04441_),
    .Y(_04840_));
 INVx1_ASAP7_75t_R _27230_ (.A(_04589_),
    .Y(_04841_));
 OAI21x1_ASAP7_75t_R _27231_ (.A1(_04451_),
    .A2(_04841_),
    .B(_04456_),
    .Y(_04842_));
 AOI21x1_ASAP7_75t_R _27232_ (.A1(_04840_),
    .A2(_04842_),
    .B(_04521_),
    .Y(_04843_));
 INVx1_ASAP7_75t_R _27233_ (.A(_04605_),
    .Y(_04844_));
 NAND2x1_ASAP7_75t_SL _27234_ (.A(_04720_),
    .B(_04454_),
    .Y(_04845_));
 AOI21x1_ASAP7_75t_R _27235_ (.A1(_04844_),
    .A2(_04845_),
    .B(_04441_),
    .Y(_04846_));
 INVx1_ASAP7_75t_SL _27236_ (.A(_04649_),
    .Y(_04847_));
 NAND2x1_ASAP7_75t_R _27237_ (.A(_04482_),
    .B(_04847_),
    .Y(_04848_));
 AOI21x1_ASAP7_75t_R _27238_ (.A1(_04669_),
    .A2(_04848_),
    .B(_04456_),
    .Y(_04849_));
 NOR2x1_ASAP7_75t_SL _27239_ (.A(_04846_),
    .B(_04849_),
    .Y(_04850_));
 OAI21x1_ASAP7_75t_R _27240_ (.A1(_04496_),
    .A2(_04850_),
    .B(_04464_),
    .Y(_04851_));
 AND2x2_ASAP7_75t_R _27241_ (.A(_04602_),
    .B(_04696_),
    .Y(_04852_));
 OAI21x1_ASAP7_75t_R _27242_ (.A1(_04406_),
    .A2(_04407_),
    .B(_01301_),
    .Y(_04853_));
 AOI21x1_ASAP7_75t_R _27243_ (.A1(_04421_),
    .A2(_04853_),
    .B(_04456_),
    .Y(_04854_));
 INVx1_ASAP7_75t_R _27244_ (.A(_04625_),
    .Y(_04855_));
 AOI21x1_ASAP7_75t_R _27245_ (.A1(_04854_),
    .A2(_04855_),
    .B(_04496_),
    .Y(_04856_));
 OAI21x1_ASAP7_75t_R _27246_ (.A1(_04852_),
    .A2(_04519_),
    .B(_04856_),
    .Y(_04857_));
 OA21x2_ASAP7_75t_R _27247_ (.A1(_04431_),
    .A2(_04433_),
    .B(_04456_),
    .Y(_04858_));
 AO21x1_ASAP7_75t_R _27248_ (.A1(_04402_),
    .A2(_04428_),
    .B(_04421_),
    .Y(_04859_));
 AOI21x1_ASAP7_75t_R _27249_ (.A1(_04858_),
    .A2(_04859_),
    .B(_04521_),
    .Y(_04860_));
 NAND2x1_ASAP7_75t_SL _27250_ (.A(_04500_),
    .B(_04799_),
    .Y(_04861_));
 NOR2x1_ASAP7_75t_SL _27251_ (.A(_04456_),
    .B(_04611_),
    .Y(_04862_));
 NAND2x1_ASAP7_75t_R _27252_ (.A(_04861_),
    .B(_04862_),
    .Y(_04863_));
 AOI21x1_ASAP7_75t_R _27253_ (.A1(_04860_),
    .A2(_04863_),
    .B(_04464_),
    .Y(_04864_));
 AOI21x1_ASAP7_75t_R _27254_ (.A1(_04857_),
    .A2(_04864_),
    .B(_04680_),
    .Y(_04865_));
 OAI21x1_ASAP7_75t_SL _27255_ (.A1(_04843_),
    .A2(_04851_),
    .B(_04865_),
    .Y(_04866_));
 OAI21x1_ASAP7_75t_SL _27256_ (.A1(_04822_),
    .A2(_04836_),
    .B(_04866_),
    .Y(_00124_));
 AOI21x1_ASAP7_75t_SL _27257_ (.A1(_04756_),
    .A2(_04617_),
    .B(_04521_),
    .Y(_04867_));
 NOR2x1_ASAP7_75t_SL _27258_ (.A(_04441_),
    .B(_04794_),
    .Y(_04868_));
 AO21x1_ASAP7_75t_SL _27259_ (.A1(_04527_),
    .A2(_04779_),
    .B(_04433_),
    .Y(_04869_));
 NAND2x1_ASAP7_75t_SL _27260_ (.A(_04868_),
    .B(_04869_),
    .Y(_04870_));
 AOI21x1_ASAP7_75t_SL _27261_ (.A1(_04867_),
    .A2(_04870_),
    .B(_04464_),
    .Y(_04871_));
 NAND2x1_ASAP7_75t_SL _27262_ (.A(_04433_),
    .B(_01305_),
    .Y(_04872_));
 AOI21x1_ASAP7_75t_SL _27263_ (.A1(_04872_),
    .A2(_04455_),
    .B(_04441_),
    .Y(_04873_));
 NAND2x1_ASAP7_75t_SL _27264_ (.A(_04500_),
    .B(_04710_),
    .Y(_04874_));
 NAND2x1_ASAP7_75t_SL _27265_ (.A(_04430_),
    .B(_04655_),
    .Y(_04875_));
 AOI21x1_ASAP7_75t_SL _27266_ (.A1(_04874_),
    .A2(_04875_),
    .B(_04456_),
    .Y(_04876_));
 OAI21x1_ASAP7_75t_SL _27267_ (.A1(_04873_),
    .A2(_04876_),
    .B(_04521_),
    .Y(_04877_));
 AOI21x1_ASAP7_75t_SL _27268_ (.A1(_04877_),
    .A2(_04871_),
    .B(_04680_),
    .Y(_04878_));
 AND2x2_ASAP7_75t_SL _27269_ (.A(_04518_),
    .B(_04421_),
    .Y(_04879_));
 AO21x1_ASAP7_75t_SL _27270_ (.A1(_01306_),
    .A2(_04433_),
    .B(_04441_),
    .Y(_04880_));
 OA21x2_ASAP7_75t_SL _27271_ (.A1(_04879_),
    .A2(_04880_),
    .B(_04496_),
    .Y(_04881_));
 NAND2x1_ASAP7_75t_SL _27272_ (.A(_04479_),
    .B(_04485_),
    .Y(_04882_));
 NOR2x1_ASAP7_75t_SL _27273_ (.A(_04705_),
    .B(_04429_),
    .Y(_04883_));
 OA21x2_ASAP7_75t_SL _27274_ (.A1(_04883_),
    .A2(_04433_),
    .B(_04441_),
    .Y(_04884_));
 NAND2x1_ASAP7_75t_SL _27275_ (.A(_04882_),
    .B(_04884_),
    .Y(_04885_));
 AOI21x1_ASAP7_75t_SL _27276_ (.A1(_04881_),
    .A2(_04885_),
    .B(_04468_),
    .Y(_04886_));
 AOI21x1_ASAP7_75t_SL _27277_ (.A1(_04583_),
    .A2(_04445_),
    .B(_04433_),
    .Y(_04887_));
 OA21x2_ASAP7_75t_SL _27278_ (.A1(_04564_),
    .A2(_04421_),
    .B(_04441_),
    .Y(_04888_));
 NAND2x1_ASAP7_75t_SL _27279_ (.A(_04720_),
    .B(_04879_),
    .Y(_04889_));
 AOI21x1_ASAP7_75t_SL _27280_ (.A1(_04888_),
    .A2(_04889_),
    .B(_04496_),
    .Y(_04890_));
 OAI21x1_ASAP7_75t_SL _27281_ (.A1(_04519_),
    .A2(_04887_),
    .B(_04890_),
    .Y(_04891_));
 NAND2x1_ASAP7_75t_SL _27282_ (.A(_04886_),
    .B(_04891_),
    .Y(_04892_));
 NAND2x1_ASAP7_75t_SL _27283_ (.A(_04878_),
    .B(_04892_),
    .Y(_04893_));
 AO21x1_ASAP7_75t_SL _27284_ (.A1(_04402_),
    .A2(_01303_),
    .B(_04456_),
    .Y(_04894_));
 OA21x2_ASAP7_75t_SL _27285_ (.A1(_04894_),
    .A2(_04602_),
    .B(_04521_),
    .Y(_04895_));
 OA21x2_ASAP7_75t_SL _27286_ (.A1(_04433_),
    .A2(_04429_),
    .B(_04456_),
    .Y(_04896_));
 AOI22x1_ASAP7_75t_SL _27287_ (.A1(_04433_),
    .A2(_04578_),
    .B1(_04605_),
    .B2(_04448_),
    .Y(_04897_));
 NAND2x1_ASAP7_75t_SL _27288_ (.A(_04896_),
    .B(_04897_),
    .Y(_04898_));
 AOI21x1_ASAP7_75t_SL _27289_ (.A1(_04895_),
    .A2(_04898_),
    .B(_04468_),
    .Y(_04899_));
 NAND2x1_ASAP7_75t_SL _27290_ (.A(_04428_),
    .B(_04605_),
    .Y(_04900_));
 NAND2x1_ASAP7_75t_SL _27291_ (.A(_04694_),
    .B(_04676_),
    .Y(_04901_));
 AOI21x1_ASAP7_75t_SL _27292_ (.A1(_04900_),
    .A2(_04901_),
    .B(_04456_),
    .Y(_04902_));
 NOR2x1_ASAP7_75t_SL _27293_ (.A(_04433_),
    .B(_04705_),
    .Y(_04903_));
 AOI211x1_ASAP7_75t_SL _27294_ (.A1(_04485_),
    .A2(_04410_),
    .B(_04441_),
    .C(_04903_),
    .Y(_04904_));
 OAI21x1_ASAP7_75t_SL _27295_ (.A1(_04902_),
    .A2(_04904_),
    .B(_04496_),
    .Y(_04905_));
 AOI21x1_ASAP7_75t_SL _27296_ (.A1(_04899_),
    .A2(_04905_),
    .B(_04541_),
    .Y(_04906_));
 AND2x2_ASAP7_75t_SL _27297_ (.A(_04532_),
    .B(_04642_),
    .Y(_04907_));
 NOR2x1_ASAP7_75t_SL _27298_ (.A(_04421_),
    .B(_04630_),
    .Y(_04908_));
 AO21x1_ASAP7_75t_SL _27299_ (.A1(_04908_),
    .A2(_04564_),
    .B(_04456_),
    .Y(_04909_));
 NOR2x1_ASAP7_75t_SL _27300_ (.A(_04907_),
    .B(_04909_),
    .Y(_04910_));
 AO21x1_ASAP7_75t_SL _27301_ (.A1(_01298_),
    .A2(_04433_),
    .B(_04441_),
    .Y(_04911_));
 OAI21x1_ASAP7_75t_SL _27302_ (.A1(_04911_),
    .A2(_04839_),
    .B(_04496_),
    .Y(_04912_));
 NOR2x1_ASAP7_75t_SL _27303_ (.A(_04910_),
    .B(_04912_),
    .Y(_04913_));
 NAND2x1_ASAP7_75t_SL _27304_ (.A(_04720_),
    .B(_04531_),
    .Y(_04914_));
 INVx1_ASAP7_75t_SL _27305_ (.A(_04517_),
    .Y(_04915_));
 AOI21x1_ASAP7_75t_SL _27306_ (.A1(_04914_),
    .A2(_04915_),
    .B(_04441_),
    .Y(_04916_));
 INVx1_ASAP7_75t_SL _27307_ (.A(_04544_),
    .Y(_04917_));
 AOI21x1_ASAP7_75t_SL _27308_ (.A1(_04565_),
    .A2(_04570_),
    .B(_04433_),
    .Y(_04918_));
 AOI21x1_ASAP7_75t_SL _27309_ (.A1(_04917_),
    .A2(_04702_),
    .B(_04918_),
    .Y(_04919_));
 OAI21x1_ASAP7_75t_SL _27310_ (.A1(_04456_),
    .A2(_04919_),
    .B(_04521_),
    .Y(_04920_));
 NOR2x1_ASAP7_75t_SL _27311_ (.A(_04916_),
    .B(_04920_),
    .Y(_04921_));
 OAI21x1_ASAP7_75t_SL _27312_ (.A1(_04913_),
    .A2(_04921_),
    .B(_04468_),
    .Y(_04922_));
 NAND2x1_ASAP7_75t_SL _27313_ (.A(_04906_),
    .B(_04922_),
    .Y(_04923_));
 NAND2x1_ASAP7_75t_SL _27314_ (.A(_04893_),
    .B(_04923_),
    .Y(_00125_));
 AND2x2_ASAP7_75t_SL _27315_ (.A(_04618_),
    .B(_04464_),
    .Y(_04924_));
 AO21x1_ASAP7_75t_SL _27316_ (.A1(_04529_),
    .A2(_04924_),
    .B(_04456_),
    .Y(_04925_));
 AND2x2_ASAP7_75t_SL _27317_ (.A(_04829_),
    .B(_04601_),
    .Y(_04926_));
 AOI211x1_ASAP7_75t_SL _27318_ (.A1(_04759_),
    .A2(_04433_),
    .B(_04926_),
    .C(_04464_),
    .Y(_04927_));
 OAI21x1_ASAP7_75t_SL _27319_ (.A1(_04925_),
    .A2(_04927_),
    .B(_04521_),
    .Y(_04928_));
 AND3x1_ASAP7_75t_SL _27320_ (.A(_04500_),
    .B(_04421_),
    .C(_04527_),
    .Y(_04929_));
 AO21x1_ASAP7_75t_SL _27321_ (.A1(_04433_),
    .A2(_04759_),
    .B(_04929_),
    .Y(_04930_));
 OA21x2_ASAP7_75t_SL _27322_ (.A1(_04624_),
    .A2(_04433_),
    .B(_04464_),
    .Y(_04931_));
 AO21x1_ASAP7_75t_SL _27323_ (.A1(_04897_),
    .A2(_04931_),
    .B(_04441_),
    .Y(_04932_));
 AOI21x1_ASAP7_75t_SL _27324_ (.A1(_04468_),
    .A2(_04930_),
    .B(_04932_),
    .Y(_04933_));
 NOR2x1_ASAP7_75t_SL _27325_ (.A(_04928_),
    .B(_04933_),
    .Y(_04934_));
 NAND2x1_ASAP7_75t_SL _27326_ (.A(_04464_),
    .B(_04725_),
    .Y(_04935_));
 AOI21x1_ASAP7_75t_SL _27327_ (.A1(_04786_),
    .A2(_04861_),
    .B(_04456_),
    .Y(_04936_));
 NOR2x1_ASAP7_75t_SL _27328_ (.A(_04935_),
    .B(_04936_),
    .Y(_04937_));
 AO21x1_ASAP7_75t_SL _27329_ (.A1(_01312_),
    .A2(_04433_),
    .B(_04441_),
    .Y(_04938_));
 AO21x1_ASAP7_75t_SL _27330_ (.A1(_04500_),
    .A2(_04710_),
    .B(_04938_),
    .Y(_04939_));
 AOI21x1_ASAP7_75t_SL _27331_ (.A1(_04624_),
    .A2(_04720_),
    .B(_04421_),
    .Y(_04940_));
 OAI21x1_ASAP7_75t_SL _27332_ (.A1(_04772_),
    .A2(_04940_),
    .B(_04441_),
    .Y(_04941_));
 AOI21x1_ASAP7_75t_SL _27333_ (.A1(_04939_),
    .A2(_04941_),
    .B(_04464_),
    .Y(_04942_));
 OAI21x1_ASAP7_75t_SL _27334_ (.A1(_04937_),
    .A2(_04942_),
    .B(_04496_),
    .Y(_04943_));
 NAND2x1_ASAP7_75t_SL _27335_ (.A(_04541_),
    .B(_04943_),
    .Y(_04944_));
 AND2x2_ASAP7_75t_SL _27336_ (.A(_04825_),
    .B(_04601_),
    .Y(_04945_));
 NOR2x1_ASAP7_75t_SL _27337_ (.A(_04433_),
    .B(_04555_),
    .Y(_04946_));
 AO21x1_ASAP7_75t_SL _27338_ (.A1(_04946_),
    .A2(_04742_),
    .B(_04468_),
    .Y(_04947_));
 NAND2x1_ASAP7_75t_SL _27339_ (.A(_04500_),
    .B(_04655_),
    .Y(_04948_));
 AOI21x1_ASAP7_75t_SL _27340_ (.A1(_04624_),
    .A2(_04676_),
    .B(_04464_),
    .Y(_04949_));
 AOI21x1_ASAP7_75t_SL _27341_ (.A1(_04948_),
    .A2(_04949_),
    .B(_04441_),
    .Y(_04950_));
 OAI21x1_ASAP7_75t_SL _27342_ (.A1(_04945_),
    .A2(_04947_),
    .B(_04950_),
    .Y(_04951_));
 AOI21x1_ASAP7_75t_R _27343_ (.A1(_04402_),
    .A2(_01302_),
    .B(_04421_),
    .Y(_04952_));
 NOR2x1_ASAP7_75t_SL _27344_ (.A(_04433_),
    .B(_04564_),
    .Y(_04953_));
 AOI21x1_ASAP7_75t_SL _27345_ (.A1(_04685_),
    .A2(_04952_),
    .B(_04953_),
    .Y(_04954_));
 AOI21x1_ASAP7_75t_SL _27346_ (.A1(_04421_),
    .A2(_04429_),
    .B(_04464_),
    .Y(_04955_));
 NAND2x1_ASAP7_75t_SL _27347_ (.A(_04747_),
    .B(_04955_),
    .Y(_04956_));
 OAI21x1_ASAP7_75t_SL _27348_ (.A1(_04468_),
    .A2(_04954_),
    .B(_04956_),
    .Y(_04957_));
 AOI21x1_ASAP7_75t_SL _27349_ (.A1(_04441_),
    .A2(_04957_),
    .B(_04521_),
    .Y(_04958_));
 NAND2x1_ASAP7_75t_SL _27350_ (.A(_04951_),
    .B(_04958_),
    .Y(_04959_));
 AOI21x1_ASAP7_75t_R _27351_ (.A1(_04502_),
    .A2(_04503_),
    .B(_04431_),
    .Y(_04960_));
 OAI21x1_ASAP7_75t_SL _27352_ (.A1(_04960_),
    .A2(_04515_),
    .B(_04433_),
    .Y(_04961_));
 NAND2x1_ASAP7_75t_SL _27353_ (.A(_04510_),
    .B(_04710_),
    .Y(_04962_));
 AOI21x1_ASAP7_75t_SL _27354_ (.A1(_04961_),
    .A2(_04962_),
    .B(_04441_),
    .Y(_04963_));
 OAI21x1_ASAP7_75t_SL _27355_ (.A1(_04578_),
    .A2(_04545_),
    .B(_04433_),
    .Y(_04964_));
 NAND2x1_ASAP7_75t_SL _27356_ (.A(_04696_),
    .B(_04454_),
    .Y(_04965_));
 AOI21x1_ASAP7_75t_SL _27357_ (.A1(_04964_),
    .A2(_04965_),
    .B(_04456_),
    .Y(_04966_));
 OAI21x1_ASAP7_75t_SL _27358_ (.A1(_04963_),
    .A2(_04966_),
    .B(_04464_),
    .Y(_04967_));
 INVx1_ASAP7_75t_R _27359_ (.A(_01301_),
    .Y(_04968_));
 NAND2x1_ASAP7_75t_SL _27360_ (.A(_04968_),
    .B(_04605_),
    .Y(_04969_));
 NAND3x1_ASAP7_75t_SL _27361_ (.A(_04969_),
    .B(_04807_),
    .C(_04739_),
    .Y(_04970_));
 AND2x2_ASAP7_75t_SL _27362_ (.A(_01311_),
    .B(_01317_),
    .Y(_04971_));
 OA21x2_ASAP7_75t_SL _27363_ (.A1(_04433_),
    .A2(_04971_),
    .B(_04456_),
    .Y(_04972_));
 OAI21x1_ASAP7_75t_SL _27364_ (.A1(_04755_),
    .A2(_04838_),
    .B(_04433_),
    .Y(_04973_));
 AOI21x1_ASAP7_75t_SL _27365_ (.A1(_04972_),
    .A2(_04973_),
    .B(_04464_),
    .Y(_04974_));
 AOI21x1_ASAP7_75t_SL _27366_ (.A1(_04970_),
    .A2(_04974_),
    .B(_04496_),
    .Y(_04975_));
 AOI21x1_ASAP7_75t_SL _27367_ (.A1(_04967_),
    .A2(_04975_),
    .B(_04541_),
    .Y(_04976_));
 NAND2x1_ASAP7_75t_SL _27368_ (.A(_04959_),
    .B(_04976_),
    .Y(_04977_));
 OAI21x1_ASAP7_75t_SL _27369_ (.A1(_04934_),
    .A2(_04944_),
    .B(_04977_),
    .Y(_00126_));
 AOI211x1_ASAP7_75t_SL _27370_ (.A1(_04430_),
    .A2(_04421_),
    .B(_04908_),
    .C(_04441_),
    .Y(_04978_));
 NOR2x1_ASAP7_75t_SL _27371_ (.A(_04434_),
    .B(_04825_),
    .Y(_04979_));
 AO21x1_ASAP7_75t_SL _27372_ (.A1(_04623_),
    .A2(_04421_),
    .B(_04456_),
    .Y(_04980_));
 OAI21x1_ASAP7_75t_SL _27373_ (.A1(_04979_),
    .A2(_04980_),
    .B(_04464_),
    .Y(_04981_));
 OAI21x1_ASAP7_75t_SL _27374_ (.A1(_04978_),
    .A2(_04981_),
    .B(_04541_),
    .Y(_04982_));
 NAND2x1_ASAP7_75t_SL _27375_ (.A(_04500_),
    .B(_04434_),
    .Y(_04983_));
 NAND2x1_ASAP7_75t_SL _27376_ (.A(_04983_),
    .B(_04691_),
    .Y(_04984_));
 NOR2x1_ASAP7_75t_SL _27377_ (.A(_04433_),
    .B(_01305_),
    .Y(_04985_));
 OAI21x1_ASAP7_75t_SL _27378_ (.A1(_04985_),
    .A2(_04819_),
    .B(_04441_),
    .Y(_04986_));
 AOI21x1_ASAP7_75t_SL _27379_ (.A1(_04984_),
    .A2(_04986_),
    .B(_04464_),
    .Y(_04987_));
 OAI21x1_ASAP7_75t_SL _27380_ (.A1(_04982_),
    .A2(_04987_),
    .B(_04496_),
    .Y(_04988_));
 INVx1_ASAP7_75t_SL _27381_ (.A(_04862_),
    .Y(_04989_));
 OAI21x1_ASAP7_75t_SL _27382_ (.A1(_04433_),
    .A2(_04472_),
    .B(_04669_),
    .Y(_04990_));
 AND3x1_ASAP7_75t_SL _27383_ (.A(_04402_),
    .B(_04968_),
    .C(_04421_),
    .Y(_04991_));
 AO21x1_ASAP7_75t_SL _27384_ (.A1(_01308_),
    .A2(_04433_),
    .B(_04441_),
    .Y(_04992_));
 OA21x2_ASAP7_75t_SL _27385_ (.A1(_04991_),
    .A2(_04992_),
    .B(_04468_),
    .Y(_04993_));
 OAI21x1_ASAP7_75t_SL _27386_ (.A1(_04989_),
    .A2(_04990_),
    .B(_04993_),
    .Y(_04994_));
 AND3x1_ASAP7_75t_SL _27387_ (.A(_04591_),
    .B(_04624_),
    .C(_04433_),
    .Y(_04995_));
 AO21x1_ASAP7_75t_SL _27388_ (.A1(_04532_),
    .A2(_04500_),
    .B(_04456_),
    .Y(_04996_));
 NAND2x1_ASAP7_75t_SL _27389_ (.A(_04421_),
    .B(_04475_),
    .Y(_04997_));
 OAI21x1_ASAP7_75t_R _27390_ (.A1(_01317_),
    .A2(_04421_),
    .B(_04456_),
    .Y(_04998_));
 AOI21x1_ASAP7_75t_SL _27391_ (.A1(_04421_),
    .A2(_04578_),
    .B(_04998_),
    .Y(_04999_));
 AOI21x1_ASAP7_75t_SL _27392_ (.A1(_04997_),
    .A2(_04999_),
    .B(_04468_),
    .Y(_05000_));
 OAI21x1_ASAP7_75t_SL _27393_ (.A1(_04995_),
    .A2(_04996_),
    .B(_05000_),
    .Y(_05001_));
 AOI21x1_ASAP7_75t_SL _27394_ (.A1(_04994_),
    .A2(_05001_),
    .B(_04541_),
    .Y(_05002_));
 NOR2x1_ASAP7_75t_SL _27395_ (.A(_04988_),
    .B(_05002_),
    .Y(_05003_));
 OAI21x1_ASAP7_75t_SL _27396_ (.A1(_04960_),
    .A2(_04637_),
    .B(_04421_),
    .Y(_05004_));
 OAI21x1_ASAP7_75t_SL _27397_ (.A1(_04429_),
    .A2(_04661_),
    .B(_04433_),
    .Y(_05005_));
 AOI21x1_ASAP7_75t_SL _27398_ (.A1(_05004_),
    .A2(_05005_),
    .B(_04441_),
    .Y(_05006_));
 NAND2x1_ASAP7_75t_SL _27399_ (.A(_04694_),
    .B(_04434_),
    .Y(_05007_));
 AOI21x1_ASAP7_75t_SL _27400_ (.A1(_04800_),
    .A2(_05007_),
    .B(_04456_),
    .Y(_05008_));
 OAI21x1_ASAP7_75t_SL _27401_ (.A1(_05006_),
    .A2(_05008_),
    .B(_04468_),
    .Y(_05009_));
 OAI21x1_ASAP7_75t_SL _27402_ (.A1(_04676_),
    .A2(_04952_),
    .B(_04549_),
    .Y(_05010_));
 NAND2x1_ASAP7_75t_SL _27403_ (.A(_04456_),
    .B(_05010_),
    .Y(_05011_));
 AND2x2_ASAP7_75t_SL _27404_ (.A(_04627_),
    .B(_04441_),
    .Y(_05012_));
 AOI21x1_ASAP7_75t_SL _27405_ (.A1(_05012_),
    .A2(_04973_),
    .B(_04468_),
    .Y(_05013_));
 AOI21x1_ASAP7_75t_SL _27406_ (.A1(_05011_),
    .A2(_05013_),
    .B(_04541_),
    .Y(_05014_));
 NAND2x1_ASAP7_75t_SL _27407_ (.A(_05009_),
    .B(_05014_),
    .Y(_05015_));
 NAND2x1_ASAP7_75t_SL _27408_ (.A(_04793_),
    .B(_04615_),
    .Y(_05016_));
 AOI21x1_ASAP7_75t_SL _27409_ (.A1(_04510_),
    .A2(_04710_),
    .B(_04441_),
    .Y(_05017_));
 AOI21x1_ASAP7_75t_SL _27410_ (.A1(_04683_),
    .A2(_05017_),
    .B(_04468_),
    .Y(_05018_));
 OAI21x1_ASAP7_75t_SL _27411_ (.A1(_04456_),
    .A2(_05016_),
    .B(_05018_),
    .Y(_05019_));
 NAND2x1_ASAP7_75t_SL _27412_ (.A(_04685_),
    .B(_04532_),
    .Y(_05020_));
 OAI21x1_ASAP7_75t_SL _27413_ (.A1(_04960_),
    .A2(_04637_),
    .B(_04433_),
    .Y(_05021_));
 NAND3x1_ASAP7_75t_SL _27414_ (.A(_05020_),
    .B(_04441_),
    .C(_05021_),
    .Y(_05022_));
 AOI21x1_ASAP7_75t_SL _27415_ (.A1(_04500_),
    .A2(_04799_),
    .B(_04829_),
    .Y(_05023_));
 AOI21x1_ASAP7_75t_SL _27416_ (.A1(_04456_),
    .A2(_05023_),
    .B(_04464_),
    .Y(_05024_));
 AOI21x1_ASAP7_75t_SL _27417_ (.A1(_05022_),
    .A2(_05024_),
    .B(_04680_),
    .Y(_05025_));
 NAND2x1_ASAP7_75t_SL _27418_ (.A(_05019_),
    .B(_05025_),
    .Y(_05026_));
 AOI21x1_ASAP7_75t_SL _27419_ (.A1(_05015_),
    .A2(_05026_),
    .B(_04496_),
    .Y(_05027_));
 NOR2x1_ASAP7_75t_SL _27420_ (.A(_05003_),
    .B(_05027_),
    .Y(_00127_));
 NOR2x1_ASAP7_75t_R _27421_ (.A(_00574_),
    .B(_00480_),
    .Y(_05028_));
 XOR2x2_ASAP7_75t_SL _27422_ (.A(_10706_),
    .B(_02307_),
    .Y(_05029_));
 XOR2x2_ASAP7_75t_SL _27423_ (.A(_00575_),
    .B(_00582_),
    .Y(_05030_));
 XOR2x2_ASAP7_75t_SL _27424_ (.A(_05030_),
    .B(_00640_),
    .Y(_05031_));
 XOR2x2_ASAP7_75t_SL _27425_ (.A(_05029_),
    .B(_05031_),
    .Y(_05032_));
 NOR2x1p5_ASAP7_75t_L _27426_ (.A(_10675_),
    .B(_05032_),
    .Y(_05033_));
 OAI21x1_ASAP7_75t_R _27427_ (.A1(_05028_),
    .A2(_05033_),
    .B(_00849_),
    .Y(_05034_));
 AND2x2_ASAP7_75t_R _27428_ (.A(_10675_),
    .B(_00480_),
    .Y(_05035_));
 XNOR2x2_ASAP7_75t_SL _27429_ (.A(_05031_),
    .B(_05029_),
    .Y(_05036_));
 NOR2x1p5_ASAP7_75t_SL _27430_ (.A(_10675_),
    .B(_05036_),
    .Y(_05037_));
 INVx1_ASAP7_75t_R _27431_ (.A(_00849_),
    .Y(_05038_));
 OAI21x1_ASAP7_75t_R _27432_ (.A1(_05035_),
    .A2(_05037_),
    .B(_05038_),
    .Y(_05039_));
 NAND2x2_ASAP7_75t_SL _27433_ (.A(_05039_),
    .B(_05034_),
    .Y(_05040_));
 NAND2x1p5_ASAP7_75t_L _27435_ (.A(_00481_),
    .B(_10675_),
    .Y(_05041_));
 XOR2x2_ASAP7_75t_SL _27436_ (.A(_10696_),
    .B(_10879_),
    .Y(_05042_));
 XOR2x2_ASAP7_75t_L _27437_ (.A(_05042_),
    .B(_10666_),
    .Y(_05043_));
 NAND2x1_ASAP7_75t_L _27438_ (.A(_00574_),
    .B(_05043_),
    .Y(_05044_));
 INVx1_ASAP7_75t_R _27439_ (.A(_00838_),
    .Y(_05045_));
 AOI21x1_ASAP7_75t_SL _27440_ (.A1(_05041_),
    .A2(_05044_),
    .B(_05045_),
    .Y(_05046_));
 OR2x2_ASAP7_75t_L _27441_ (.A(_00574_),
    .B(_00481_),
    .Y(_05047_));
 XOR2x2_ASAP7_75t_L _27442_ (.A(_05042_),
    .B(_05030_),
    .Y(_05048_));
 NAND2x1p5_ASAP7_75t_L _27443_ (.A(_00574_),
    .B(_05048_),
    .Y(_05049_));
 AOI21x1_ASAP7_75t_R _27444_ (.A1(_05047_),
    .A2(_05049_),
    .B(_00838_),
    .Y(_05050_));
 NOR2x2_ASAP7_75t_SL _27445_ (.A(_05046_),
    .B(_05050_),
    .Y(_05051_));
 NOR2x1_ASAP7_75t_R _27447_ (.A(_00574_),
    .B(_00482_),
    .Y(_05052_));
 XOR2x2_ASAP7_75t_SL _27448_ (.A(_00576_),
    .B(_00641_),
    .Y(_05053_));
 NAND2x1_ASAP7_75t_L _27449_ (.A(_02308_),
    .B(_05053_),
    .Y(_05054_));
 XNOR2x2_ASAP7_75t_SL _27450_ (.A(_00576_),
    .B(_00641_),
    .Y(_05055_));
 NAND2x1_ASAP7_75t_R _27451_ (.A(_00672_),
    .B(_05055_),
    .Y(_05056_));
 AOI21x1_ASAP7_75t_SL _27452_ (.A1(_05054_),
    .A2(_05056_),
    .B(_02338_),
    .Y(_05057_));
 INVx1_ASAP7_75t_SL _27453_ (.A(_05057_),
    .Y(_05058_));
 NAND3x1_ASAP7_75t_R _27454_ (.A(_05056_),
    .B(_05054_),
    .C(_02338_),
    .Y(_05059_));
 AOI21x1_ASAP7_75t_SL _27455_ (.A1(_05058_),
    .A2(_05059_),
    .B(_10675_),
    .Y(_05060_));
 INVx1_ASAP7_75t_R _27456_ (.A(_00860_),
    .Y(_05061_));
 OAI21x1_ASAP7_75t_SL _27457_ (.A1(_05052_),
    .A2(_05060_),
    .B(_05061_),
    .Y(_05062_));
 XOR2x2_ASAP7_75t_SL _27458_ (.A(_05053_),
    .B(_00672_),
    .Y(_05063_));
 NOR2x1_ASAP7_75t_SL _27459_ (.A(_02337_),
    .B(_05063_),
    .Y(_05064_));
 OAI21x1_ASAP7_75t_SL _27460_ (.A1(_05057_),
    .A2(_05064_),
    .B(_00574_),
    .Y(_05065_));
 INVx1_ASAP7_75t_L _27461_ (.A(_05052_),
    .Y(_05066_));
 NAND3x1_ASAP7_75t_SL _27462_ (.A(_05065_),
    .B(_00860_),
    .C(_05066_),
    .Y(_05067_));
 NAND2x2_ASAP7_75t_SL _27463_ (.A(_05062_),
    .B(_05067_),
    .Y(_05068_));
 AOI21x1_ASAP7_75t_SL _27465_ (.A1(_05049_),
    .A2(_05047_),
    .B(_05045_),
    .Y(_05069_));
 AOI21x1_ASAP7_75t_SL _27466_ (.A1(_05041_),
    .A2(_05044_),
    .B(_00838_),
    .Y(_05070_));
 NOR2x2_ASAP7_75t_SL _27467_ (.A(_05070_),
    .B(_05069_),
    .Y(_05071_));
 OAI21x1_ASAP7_75t_SL _27469_ (.A1(_05052_),
    .A2(_05060_),
    .B(_00860_),
    .Y(_05072_));
 NAND3x2_ASAP7_75t_SL _27470_ (.B(_05061_),
    .C(_05066_),
    .Y(_05073_),
    .A(_05065_));
 NAND2x2_ASAP7_75t_SL _27471_ (.A(_05072_),
    .B(_05073_),
    .Y(_05074_));
 XNOR2x2_ASAP7_75t_R _27473_ (.A(_00642_),
    .B(_10761_),
    .Y(_05075_));
 NOR2x1_ASAP7_75t_R _27474_ (.A(_05075_),
    .B(_02367_),
    .Y(_05076_));
 AO21x1_ASAP7_75t_SL _27475_ (.A1(_02367_),
    .A2(_05075_),
    .B(_10675_),
    .Y(_05077_));
 NAND2x1_ASAP7_75t_R _27476_ (.A(_00489_),
    .B(_10675_),
    .Y(_05078_));
 OAI21x1_ASAP7_75t_SL _27477_ (.A1(_05076_),
    .A2(_05077_),
    .B(_05078_),
    .Y(_05079_));
 XOR2x2_ASAP7_75t_SL _27478_ (.A(_05079_),
    .B(_00863_),
    .Y(_05080_));
 AOI21x1_ASAP7_75t_SL _27484_ (.A1(_05062_),
    .A2(_05067_),
    .B(_01326_),
    .Y(_05086_));
 AOI21x1_ASAP7_75t_SL _27486_ (.A1(_05071_),
    .A2(_05040_),
    .B(_05068_),
    .Y(_05088_));
 NOR2x1_ASAP7_75t_L _27487_ (.A(_05086_),
    .B(_05088_),
    .Y(_05089_));
 XNOR2x2_ASAP7_75t_SL _27488_ (.A(_00863_),
    .B(_05079_),
    .Y(_05090_));
 NOR2x1_ASAP7_75t_SL _27491_ (.A(_01324_),
    .B(_05074_),
    .Y(_05093_));
 NAND2x1_ASAP7_75t_R _27492_ (.A(_05090_),
    .B(_05093_),
    .Y(_05094_));
 OAI21x1_ASAP7_75t_SL _27493_ (.A1(_05080_),
    .A2(_05089_),
    .B(_05094_),
    .Y(_05095_));
 AO21x1_ASAP7_75t_R _27495_ (.A1(_05073_),
    .A2(_05072_),
    .B(_01322_),
    .Y(_05097_));
 AOI21x1_ASAP7_75t_R _27496_ (.A1(_05068_),
    .A2(_05071_),
    .B(_05090_),
    .Y(_05098_));
 XOR2x2_ASAP7_75t_R _27497_ (.A(_10748_),
    .B(_00643_),
    .Y(_05099_));
 XOR2x2_ASAP7_75t_SL _27498_ (.A(_02384_),
    .B(_05099_),
    .Y(_05100_));
 NOR2x1_ASAP7_75t_R _27499_ (.A(_00574_),
    .B(_00568_),
    .Y(_05101_));
 AOI21x1_ASAP7_75t_R _27500_ (.A1(_00574_),
    .A2(_05100_),
    .B(_05101_),
    .Y(_05102_));
 XNOR2x2_ASAP7_75t_SL _27501_ (.A(_00864_),
    .B(_05102_),
    .Y(_05103_));
 INVx3_ASAP7_75t_SL _27502_ (.A(_05103_),
    .Y(_05104_));
 AOI21x1_ASAP7_75t_R _27504_ (.A1(_05097_),
    .A2(_05098_),
    .B(_05104_),
    .Y(_05106_));
 INVx1_ASAP7_75t_R _27505_ (.A(_05106_),
    .Y(_05107_));
 INVx1_ASAP7_75t_R _27507_ (.A(_01336_),
    .Y(_05109_));
 AO21x1_ASAP7_75t_SL _27510_ (.A1(_05067_),
    .A2(_05062_),
    .B(_01323_),
    .Y(_05112_));
 NAND2x1p5_ASAP7_75t_SL _27512_ (.A(_05112_),
    .B(_05090_),
    .Y(_05114_));
 OAI21x1_ASAP7_75t_R _27513_ (.A1(_05109_),
    .A2(_05090_),
    .B(_05114_),
    .Y(_05115_));
 XOR2x2_ASAP7_75t_R _27514_ (.A(_00580_),
    .B(_00581_),
    .Y(_05116_));
 XOR2x2_ASAP7_75t_R _27515_ (.A(_05116_),
    .B(_13574_),
    .Y(_05117_));
 XOR2x2_ASAP7_75t_R _27516_ (.A(_05117_),
    .B(_10730_),
    .Y(_05118_));
 NOR2x1_ASAP7_75t_R _27517_ (.A(_00574_),
    .B(_00566_),
    .Y(_05119_));
 AO21x1_ASAP7_75t_SL _27518_ (.A1(_05118_),
    .A2(_00574_),
    .B(_05119_),
    .Y(_05120_));
 XOR2x2_ASAP7_75t_SL _27519_ (.A(_05120_),
    .B(_00866_),
    .Y(_05121_));
 INVx1_ASAP7_75t_SL _27520_ (.A(_05121_),
    .Y(_05122_));
 AOI21x1_ASAP7_75t_R _27521_ (.A1(_05104_),
    .A2(_05115_),
    .B(_05122_),
    .Y(_05123_));
 OAI21x1_ASAP7_75t_R _27522_ (.A1(_05095_),
    .A2(_05107_),
    .B(_05123_),
    .Y(_05124_));
 INVx1_ASAP7_75t_R _27523_ (.A(_05072_),
    .Y(_05125_));
 NAND2x1_ASAP7_75t_R _27524_ (.A(_00482_),
    .B(_10675_),
    .Y(_05126_));
 NAND3x1_ASAP7_75t_R _27525_ (.A(_05059_),
    .B(_05058_),
    .C(_00574_),
    .Y(_05127_));
 AOI21x1_ASAP7_75t_R _27526_ (.A1(_05126_),
    .A2(_05127_),
    .B(_00860_),
    .Y(_05128_));
 INVx1_ASAP7_75t_R _27527_ (.A(_01329_),
    .Y(_05129_));
 OAI21x1_ASAP7_75t_R _27528_ (.A1(_05125_),
    .A2(_05128_),
    .B(_05129_),
    .Y(_05130_));
 AOI21x1_ASAP7_75t_R _27529_ (.A1(_05066_),
    .A2(_05065_),
    .B(_00860_),
    .Y(_05131_));
 AOI21x1_ASAP7_75t_R _27530_ (.A1(_05126_),
    .A2(_05127_),
    .B(_05061_),
    .Y(_05132_));
 INVx2_ASAP7_75t_R _27531_ (.A(_01326_),
    .Y(_05133_));
 OAI21x1_ASAP7_75t_R _27532_ (.A1(_05131_),
    .A2(_05132_),
    .B(_05133_),
    .Y(_05134_));
 AO21x1_ASAP7_75t_R _27533_ (.A1(_05130_),
    .A2(_05134_),
    .B(_05080_),
    .Y(_05135_));
 INVx1_ASAP7_75t_SL _27535_ (.A(_01323_),
    .Y(_05137_));
 NOR2x1p5_ASAP7_75t_SL _27536_ (.A(_05137_),
    .B(_05068_),
    .Y(_05138_));
 NOR2x1p5_ASAP7_75t_SL _27537_ (.A(_05090_),
    .B(_05138_),
    .Y(_05139_));
 NOR2x1_ASAP7_75t_L _27538_ (.A(_05103_),
    .B(_05139_),
    .Y(_05140_));
 AOI21x1_ASAP7_75t_R _27540_ (.A1(_05135_),
    .A2(_05140_),
    .B(_05121_),
    .Y(_05142_));
 NAND2x1_ASAP7_75t_SL _27541_ (.A(_05051_),
    .B(_05040_),
    .Y(_05143_));
 OAI21x1_ASAP7_75t_SL _27542_ (.A1(_05068_),
    .A2(_05143_),
    .B(_05098_),
    .Y(_05144_));
 NAND2x1_ASAP7_75t_R _27544_ (.A(_05090_),
    .B(_05086_),
    .Y(_05146_));
 NAND3x1_ASAP7_75t_R _27546_ (.A(_05144_),
    .B(_05146_),
    .C(_05103_),
    .Y(_05148_));
 XOR2x2_ASAP7_75t_SL _27547_ (.A(_00579_),
    .B(_00580_),
    .Y(_05149_));
 XOR2x2_ASAP7_75t_R _27548_ (.A(_05149_),
    .B(_13550_),
    .Y(_05150_));
 XOR2x2_ASAP7_75t_SL _27549_ (.A(_05150_),
    .B(_10826_),
    .Y(_05151_));
 NOR2x1_ASAP7_75t_R _27550_ (.A(_00574_),
    .B(_00567_),
    .Y(_05152_));
 AO21x1_ASAP7_75t_R _27551_ (.A1(_05151_),
    .A2(_00574_),
    .B(_05152_),
    .Y(_05153_));
 XOR2x2_ASAP7_75t_SL _27552_ (.A(_05153_),
    .B(_00865_),
    .Y(_05154_));
 INVx1_ASAP7_75t_SL _27553_ (.A(_05154_),
    .Y(_05155_));
 AOI21x1_ASAP7_75t_R _27555_ (.A1(_05142_),
    .A2(_05148_),
    .B(_05155_),
    .Y(_05157_));
 NAND2x1_ASAP7_75t_L _27556_ (.A(_05124_),
    .B(_05157_),
    .Y(_05158_));
 AOI21x1_ASAP7_75t_SL _27557_ (.A1(_05072_),
    .A2(_05073_),
    .B(_05133_),
    .Y(_05159_));
 NOR2x1p5_ASAP7_75t_SL _27558_ (.A(_05159_),
    .B(_05090_),
    .Y(_05160_));
 NOR2x1_ASAP7_75t_R _27559_ (.A(_05103_),
    .B(_05160_),
    .Y(_05161_));
 NOR2x1_ASAP7_75t_L _27560_ (.A(_01324_),
    .B(_05068_),
    .Y(_05162_));
 INVx1_ASAP7_75t_R _27561_ (.A(_01322_),
    .Y(_05163_));
 AO21x1_ASAP7_75t_SL _27562_ (.A1(_05067_),
    .A2(_05062_),
    .B(_05163_),
    .Y(_05164_));
 INVx1_ASAP7_75t_R _27563_ (.A(_05164_),
    .Y(_05165_));
 OAI21x1_ASAP7_75t_R _27565_ (.A1(_05162_),
    .A2(_05165_),
    .B(_05090_),
    .Y(_05167_));
 AOI21x1_ASAP7_75t_R _27566_ (.A1(_05161_),
    .A2(_05167_),
    .B(_05121_),
    .Y(_05168_));
 AOI21x1_ASAP7_75t_SL _27567_ (.A1(_05074_),
    .A2(_05040_),
    .B(_05080_),
    .Y(_05169_));
 AOI21x1_ASAP7_75t_SL _27568_ (.A1(_05112_),
    .A2(_05169_),
    .B(_05104_),
    .Y(_05170_));
 NAND2x1_ASAP7_75t_L _27569_ (.A(_05074_),
    .B(_05051_),
    .Y(_05171_));
 INVx1_ASAP7_75t_SL _27570_ (.A(_01328_),
    .Y(_05172_));
 AO21x1_ASAP7_75t_R _27571_ (.A1(_05067_),
    .A2(_05062_),
    .B(_05172_),
    .Y(_05173_));
 AO21x1_ASAP7_75t_R _27572_ (.A1(_05171_),
    .A2(_05173_),
    .B(_05090_),
    .Y(_05174_));
 NAND2x1_ASAP7_75t_R _27573_ (.A(_05170_),
    .B(_05174_),
    .Y(_05175_));
 AOI21x1_ASAP7_75t_R _27576_ (.A1(_05168_),
    .A2(_05175_),
    .B(_05154_),
    .Y(_05178_));
 NAND2x1_ASAP7_75t_SL _27577_ (.A(_05071_),
    .B(_05040_),
    .Y(_05179_));
 AOI21x1_ASAP7_75t_R _27579_ (.A1(_05062_),
    .A2(_05067_),
    .B(_05129_),
    .Y(_05181_));
 NOR2x1_ASAP7_75t_SL _27580_ (.A(_05090_),
    .B(_05181_),
    .Y(_05182_));
 OAI21x1_ASAP7_75t_R _27581_ (.A1(_05068_),
    .A2(_05179_),
    .B(_05182_),
    .Y(_05183_));
 NAND2x1_ASAP7_75t_R _27582_ (.A(_05090_),
    .B(_05162_),
    .Y(_05184_));
 NAND3x1_ASAP7_75t_R _27583_ (.A(_05183_),
    .B(_05184_),
    .C(_05103_),
    .Y(_05185_));
 AO21x1_ASAP7_75t_R _27585_ (.A1(_05162_),
    .A2(_05080_),
    .B(_05103_),
    .Y(_05187_));
 INVx1_ASAP7_75t_R _27586_ (.A(_05187_),
    .Y(_05188_));
 OAI21x1_ASAP7_75t_SL _27587_ (.A1(_05033_),
    .A2(_05028_),
    .B(_05038_),
    .Y(_05189_));
 OAI21x1_ASAP7_75t_SL _27588_ (.A1(_05037_),
    .A2(_05035_),
    .B(_00849_),
    .Y(_05190_));
 NAND2x2_ASAP7_75t_SL _27589_ (.A(_05190_),
    .B(_05189_),
    .Y(_01321_));
 NOR2x1_ASAP7_75t_R _27590_ (.A(_05051_),
    .B(_01321_),
    .Y(_05191_));
 OAI21x1_ASAP7_75t_R _27591_ (.A1(_05131_),
    .A2(_05132_),
    .B(_05172_),
    .Y(_05192_));
 NAND2x1_ASAP7_75t_R _27592_ (.A(_05090_),
    .B(_05192_),
    .Y(_05193_));
 AO21x1_ASAP7_75t_R _27593_ (.A1(_05074_),
    .A2(_05191_),
    .B(_05193_),
    .Y(_05194_));
 AOI21x1_ASAP7_75t_R _27594_ (.A1(_05188_),
    .A2(_05194_),
    .B(_05122_),
    .Y(_05195_));
 NAND2x1_ASAP7_75t_SL _27595_ (.A(_05185_),
    .B(_05195_),
    .Y(_05196_));
 XOR2x2_ASAP7_75t_R _27596_ (.A(_00581_),
    .B(_00582_),
    .Y(_05197_));
 XOR2x2_ASAP7_75t_R _27597_ (.A(_05197_),
    .B(_00677_),
    .Y(_05198_));
 XOR2x2_ASAP7_75t_SL _27598_ (.A(_05198_),
    .B(_10881_),
    .Y(_05199_));
 NOR2x1_ASAP7_75t_SL _27599_ (.A(_00574_),
    .B(_00565_),
    .Y(_05200_));
 AO21x1_ASAP7_75t_SL _27600_ (.A1(_05199_),
    .A2(_00574_),
    .B(_05200_),
    .Y(_05201_));
 XOR2x2_ASAP7_75t_SL _27601_ (.A(_05201_),
    .B(_00867_),
    .Y(_05202_));
 AOI21x1_ASAP7_75t_R _27603_ (.A1(_05178_),
    .A2(_05196_),
    .B(_05202_),
    .Y(_05204_));
 NAND2x1_ASAP7_75t_SL _27604_ (.A(_05158_),
    .B(_05204_),
    .Y(_05205_));
 AOI21x1_ASAP7_75t_SL _27605_ (.A1(_05072_),
    .A2(_05073_),
    .B(_01323_),
    .Y(_05206_));
 INVx2_ASAP7_75t_SL _27606_ (.A(_05206_),
    .Y(_05207_));
 AOI21x1_ASAP7_75t_R _27607_ (.A1(_05062_),
    .A2(_05067_),
    .B(_01331_),
    .Y(_05208_));
 INVx1_ASAP7_75t_R _27608_ (.A(_05208_),
    .Y(_05209_));
 AO21x1_ASAP7_75t_SL _27609_ (.A1(_05209_),
    .A2(_05207_),
    .B(_05090_),
    .Y(_05210_));
 AOI21x1_ASAP7_75t_SL _27610_ (.A1(_05074_),
    .A2(_05071_),
    .B(_05080_),
    .Y(_05211_));
 AOI21x1_ASAP7_75t_R _27611_ (.A1(_05179_),
    .A2(_05211_),
    .B(_05103_),
    .Y(_05212_));
 NAND2x1_ASAP7_75t_L _27612_ (.A(_05210_),
    .B(_05212_),
    .Y(_05213_));
 AOI21x1_ASAP7_75t_R _27614_ (.A1(_05068_),
    .A2(_05071_),
    .B(_05080_),
    .Y(_05215_));
 NOR2x1_ASAP7_75t_R _27615_ (.A(_05104_),
    .B(_05215_),
    .Y(_05216_));
 OAI21x1_ASAP7_75t_R _27616_ (.A1(_05074_),
    .A2(_05179_),
    .B(_05160_),
    .Y(_05217_));
 AOI21x1_ASAP7_75t_R _27617_ (.A1(_05216_),
    .A2(_05217_),
    .B(_05121_),
    .Y(_05218_));
 AOI21x1_ASAP7_75t_R _27618_ (.A1(_05213_),
    .A2(_05218_),
    .B(_05154_),
    .Y(_05219_));
 AO21x1_ASAP7_75t_R _27620_ (.A1(_05073_),
    .A2(_05072_),
    .B(_05172_),
    .Y(_05221_));
 AO21x1_ASAP7_75t_R _27621_ (.A1(_05164_),
    .A2(_05221_),
    .B(_05090_),
    .Y(_05222_));
 AOI21x1_ASAP7_75t_SL _27622_ (.A1(_05051_),
    .A2(_05040_),
    .B(_05074_),
    .Y(_05223_));
 OAI21x1_ASAP7_75t_R _27623_ (.A1(_05206_),
    .A2(_05223_),
    .B(_05090_),
    .Y(_05224_));
 NAND2x1_ASAP7_75t_R _27624_ (.A(_05222_),
    .B(_05224_),
    .Y(_05225_));
 NAND2x1_ASAP7_75t_SL _27625_ (.A(_05071_),
    .B(_01321_),
    .Y(_05226_));
 AOI21x1_ASAP7_75t_SL _27626_ (.A1(_05074_),
    .A2(_05051_),
    .B(_05080_),
    .Y(_05227_));
 NAND2x1_ASAP7_75t_SL _27627_ (.A(_05226_),
    .B(_05227_),
    .Y(_05228_));
 NAND2x1_ASAP7_75t_SL _27628_ (.A(_05068_),
    .B(_05051_),
    .Y(_05229_));
 AOI21x1_ASAP7_75t_R _27630_ (.A1(_05071_),
    .A2(_05040_),
    .B(_05090_),
    .Y(_05231_));
 AOI21x1_ASAP7_75t_R _27632_ (.A1(_05229_),
    .A2(_05231_),
    .B(_05103_),
    .Y(_05233_));
 AOI21x1_ASAP7_75t_SL _27633_ (.A1(_05228_),
    .A2(_05233_),
    .B(_05122_),
    .Y(_05234_));
 OAI21x1_ASAP7_75t_R _27634_ (.A1(_05104_),
    .A2(_05225_),
    .B(_05234_),
    .Y(_05235_));
 INVx1_ASAP7_75t_SL _27635_ (.A(_05202_),
    .Y(_05236_));
 AOI21x1_ASAP7_75t_R _27636_ (.A1(_05219_),
    .A2(_05235_),
    .B(_05236_),
    .Y(_05237_));
 AO21x1_ASAP7_75t_SL _27637_ (.A1(_05207_),
    .A2(_05164_),
    .B(_05090_),
    .Y(_05238_));
 INVx1_ASAP7_75t_R _27638_ (.A(_05173_),
    .Y(_05239_));
 NAND2x1_ASAP7_75t_R _27639_ (.A(_05090_),
    .B(_05239_),
    .Y(_05240_));
 NOR2x1_ASAP7_75t_SL _27640_ (.A(_05163_),
    .B(_05068_),
    .Y(_05241_));
 AOI21x1_ASAP7_75t_R _27642_ (.A1(_05090_),
    .A2(_05241_),
    .B(_05104_),
    .Y(_05243_));
 AND3x1_ASAP7_75t_R _27643_ (.A(_05238_),
    .B(_05240_),
    .C(_05243_),
    .Y(_05244_));
 NAND2x1_ASAP7_75t_L _27644_ (.A(_05068_),
    .B(_05040_),
    .Y(_05245_));
 NAND2x1p5_ASAP7_75t_L _27645_ (.A(_05245_),
    .B(_05207_),
    .Y(_05246_));
 AOI21x1_ASAP7_75t_SL _27646_ (.A1(_05062_),
    .A2(_05067_),
    .B(_05137_),
    .Y(_05247_));
 NOR2x1p5_ASAP7_75t_SL _27647_ (.A(_05247_),
    .B(_05090_),
    .Y(_05248_));
 INVx2_ASAP7_75t_SL _27648_ (.A(_05248_),
    .Y(_05249_));
 OAI21x1_ASAP7_75t_R _27649_ (.A1(_05080_),
    .A2(_05246_),
    .B(_05249_),
    .Y(_05250_));
 AO21x1_ASAP7_75t_SL _27650_ (.A1(_05250_),
    .A2(_05104_),
    .B(_05122_),
    .Y(_05251_));
 NAND2x2_ASAP7_75t_SL _27651_ (.A(_05068_),
    .B(_01321_),
    .Y(_05252_));
 NOR2x1_ASAP7_75t_R _27652_ (.A(_05080_),
    .B(_05252_),
    .Y(_05253_));
 AO21x1_ASAP7_75t_R _27653_ (.A1(_05073_),
    .A2(_05072_),
    .B(_01324_),
    .Y(_05254_));
 OAI21x1_ASAP7_75t_R _27655_ (.A1(_05080_),
    .A2(_05254_),
    .B(_05103_),
    .Y(_05256_));
 NOR2x1_ASAP7_75t_SL _27656_ (.A(_05253_),
    .B(_05256_),
    .Y(_05257_));
 NAND2x1_ASAP7_75t_R _27657_ (.A(_05144_),
    .B(_05257_),
    .Y(_05258_));
 INVx1_ASAP7_75t_R _27658_ (.A(_01331_),
    .Y(_05259_));
 AO21x2_ASAP7_75t_L _27659_ (.A1(_05073_),
    .A2(_05072_),
    .B(_05259_),
    .Y(_05260_));
 AOI21x1_ASAP7_75t_R _27660_ (.A1(_05260_),
    .A2(_05098_),
    .B(_05103_),
    .Y(_05261_));
 NAND2x1_ASAP7_75t_SL _27661_ (.A(_05074_),
    .B(_05040_),
    .Y(_05262_));
 INVx1_ASAP7_75t_R _27662_ (.A(_05262_),
    .Y(_05263_));
 AOI21x1_ASAP7_75t_R _27663_ (.A1(_05071_),
    .A2(_05040_),
    .B(_05074_),
    .Y(_05264_));
 OAI21x1_ASAP7_75t_R _27664_ (.A1(_05263_),
    .A2(_05264_),
    .B(_05090_),
    .Y(_05265_));
 AOI21x1_ASAP7_75t_R _27665_ (.A1(_05261_),
    .A2(_05265_),
    .B(_05121_),
    .Y(_05266_));
 AOI21x1_ASAP7_75t_SL _27666_ (.A1(_05258_),
    .A2(_05266_),
    .B(_05155_),
    .Y(_05267_));
 OAI21x1_ASAP7_75t_R _27667_ (.A1(_05244_),
    .A2(_05251_),
    .B(_05267_),
    .Y(_05268_));
 NAND2x1_ASAP7_75t_SL _27668_ (.A(_05237_),
    .B(_05268_),
    .Y(_05269_));
 NAND2x1_ASAP7_75t_SL _27669_ (.A(_05205_),
    .B(_05269_),
    .Y(_00128_));
 AND3x1_ASAP7_75t_L _27670_ (.A(_05143_),
    .B(_05074_),
    .C(_05090_),
    .Y(_05270_));
 NAND2x2_ASAP7_75t_SL _27671_ (.A(_05074_),
    .B(_01321_),
    .Y(_05271_));
 NOR2x1_ASAP7_75t_SL _27672_ (.A(_05259_),
    .B(_05074_),
    .Y(_05272_));
 NOR2x1_ASAP7_75t_R _27673_ (.A(_05090_),
    .B(_05272_),
    .Y(_05273_));
 AOI21x1_ASAP7_75t_R _27674_ (.A1(_05271_),
    .A2(_05273_),
    .B(_05103_),
    .Y(_05274_));
 INVx1_ASAP7_75t_R _27675_ (.A(_05274_),
    .Y(_05275_));
 AO21x1_ASAP7_75t_R _27676_ (.A1(_05073_),
    .A2(_05072_),
    .B(_01326_),
    .Y(_05276_));
 OA21x2_ASAP7_75t_R _27677_ (.A1(_05276_),
    .A2(_05080_),
    .B(_05103_),
    .Y(_05277_));
 OAI21x1_ASAP7_75t_SL _27679_ (.A1(_05138_),
    .A2(_05223_),
    .B(_05080_),
    .Y(_05279_));
 AOI21x1_ASAP7_75t_R _27680_ (.A1(_05277_),
    .A2(_05279_),
    .B(_05154_),
    .Y(_05280_));
 OAI21x1_ASAP7_75t_R _27681_ (.A1(_05270_),
    .A2(_05275_),
    .B(_05280_),
    .Y(_05281_));
 AO21x1_ASAP7_75t_SL _27682_ (.A1(_05073_),
    .A2(_05072_),
    .B(_05137_),
    .Y(_05282_));
 NAND2x1p5_ASAP7_75t_SL _27684_ (.A(_05282_),
    .B(_05080_),
    .Y(_05284_));
 NOR2x1_ASAP7_75t_L _27685_ (.A(_05086_),
    .B(_05284_),
    .Y(_05285_));
 AOI21x1_ASAP7_75t_R _27686_ (.A1(_05068_),
    .A2(_05051_),
    .B(_05080_),
    .Y(_05286_));
 INVx1_ASAP7_75t_R _27687_ (.A(_05241_),
    .Y(_05287_));
 AND2x2_ASAP7_75t_R _27688_ (.A(_05286_),
    .B(_05287_),
    .Y(_05288_));
 OAI21x1_ASAP7_75t_SL _27689_ (.A1(_05288_),
    .A2(_05285_),
    .B(_05104_),
    .Y(_05289_));
 AOI21x1_ASAP7_75t_R _27690_ (.A1(_05112_),
    .A2(_05211_),
    .B(_05104_),
    .Y(_05290_));
 NAND2x1_ASAP7_75t_L _27691_ (.A(_05074_),
    .B(_05071_),
    .Y(_05291_));
 AO21x1_ASAP7_75t_R _27692_ (.A1(_05143_),
    .A2(_05291_),
    .B(_05090_),
    .Y(_05292_));
 AOI21x1_ASAP7_75t_R _27694_ (.A1(_05290_),
    .A2(_05292_),
    .B(_05155_),
    .Y(_05294_));
 AOI21x1_ASAP7_75t_R _27695_ (.A1(_05289_),
    .A2(_05294_),
    .B(_05121_),
    .Y(_05295_));
 NAND2x1_ASAP7_75t_L _27696_ (.A(_05281_),
    .B(_05295_),
    .Y(_05296_));
 NAND2x1_ASAP7_75t_R _27697_ (.A(_05068_),
    .B(_05080_),
    .Y(_05297_));
 INVx1_ASAP7_75t_R _27698_ (.A(_05297_),
    .Y(_05298_));
 NAND2x1_ASAP7_75t_SL _27699_ (.A(_05179_),
    .B(_05298_),
    .Y(_05299_));
 NAND2x1_ASAP7_75t_R _27700_ (.A(_05226_),
    .B(_05169_),
    .Y(_05300_));
 AOI21x1_ASAP7_75t_R _27701_ (.A1(_05299_),
    .A2(_05300_),
    .B(_05104_),
    .Y(_05301_));
 INVx1_ASAP7_75t_R _27702_ (.A(_05159_),
    .Y(_05302_));
 NAND2x1_ASAP7_75t_R _27703_ (.A(_05302_),
    .B(_05286_),
    .Y(_05303_));
 NAND2x1_ASAP7_75t_R _27704_ (.A(_05282_),
    .B(_05098_),
    .Y(_05304_));
 AOI21x1_ASAP7_75t_R _27705_ (.A1(_05303_),
    .A2(_05304_),
    .B(_05103_),
    .Y(_05305_));
 OAI21x1_ASAP7_75t_R _27706_ (.A1(_05301_),
    .A2(_05305_),
    .B(_05155_),
    .Y(_05306_));
 AOI21x1_ASAP7_75t_SL _27707_ (.A1(_05260_),
    .A2(_05248_),
    .B(_05104_),
    .Y(_05307_));
 OAI21x1_ASAP7_75t_R _27708_ (.A1(_05080_),
    .A2(_05089_),
    .B(_05307_),
    .Y(_05308_));
 AO21x1_ASAP7_75t_R _27709_ (.A1(_05086_),
    .A2(_05090_),
    .B(_05103_),
    .Y(_05309_));
 INVx1_ASAP7_75t_R _27710_ (.A(_05309_),
    .Y(_05310_));
 INVx1_ASAP7_75t_R _27711_ (.A(_05271_),
    .Y(_05311_));
 AOI21x1_ASAP7_75t_R _27712_ (.A1(_05068_),
    .A2(_05040_),
    .B(_05090_),
    .Y(_05312_));
 NOR2x1_ASAP7_75t_SL _27713_ (.A(_05311_),
    .B(_05312_),
    .Y(_05313_));
 AOI21x1_ASAP7_75t_R _27715_ (.A1(_05310_),
    .A2(_05313_),
    .B(_05155_),
    .Y(_05315_));
 AOI21x1_ASAP7_75t_R _27717_ (.A1(_05308_),
    .A2(_05315_),
    .B(_05122_),
    .Y(_05317_));
 AOI21x1_ASAP7_75t_R _27718_ (.A1(_05306_),
    .A2(_05317_),
    .B(_05202_),
    .Y(_05318_));
 NAND2x1_ASAP7_75t_SL _27719_ (.A(_05296_),
    .B(_05318_),
    .Y(_05319_));
 AOI21x1_ASAP7_75t_R _27720_ (.A1(_05068_),
    .A2(_05040_),
    .B(_05080_),
    .Y(_05320_));
 NAND2x1_ASAP7_75t_R _27721_ (.A(_05171_),
    .B(_05320_),
    .Y(_05321_));
 NAND2x1_ASAP7_75t_L _27722_ (.A(_05252_),
    .B(_05160_),
    .Y(_05322_));
 AND3x1_ASAP7_75t_R _27724_ (.A(_05321_),
    .B(_05322_),
    .C(_05154_),
    .Y(_05324_));
 AO21x1_ASAP7_75t_R _27725_ (.A1(_05067_),
    .A2(_05062_),
    .B(_01322_),
    .Y(_05325_));
 AO21x1_ASAP7_75t_R _27726_ (.A1(_05211_),
    .A2(_05325_),
    .B(_05154_),
    .Y(_05326_));
 NAND2x1_ASAP7_75t_SL _27727_ (.A(_05291_),
    .B(_05271_),
    .Y(_05327_));
 OA21x2_ASAP7_75t_R _27729_ (.A1(_05327_),
    .A2(_05264_),
    .B(_05080_),
    .Y(_05329_));
 OAI21x1_ASAP7_75t_R _27730_ (.A1(_05326_),
    .A2(_05329_),
    .B(_05104_),
    .Y(_05330_));
 AOI21x1_ASAP7_75t_R _27732_ (.A1(_05172_),
    .A2(_05068_),
    .B(_05080_),
    .Y(_05332_));
 OAI21x1_ASAP7_75t_R _27733_ (.A1(_05068_),
    .A2(_05143_),
    .B(_05332_),
    .Y(_05333_));
 INVx1_ASAP7_75t_R _27734_ (.A(_01338_),
    .Y(_05334_));
 OR3x1_ASAP7_75t_R _27735_ (.A(_05155_),
    .B(_05334_),
    .C(_05090_),
    .Y(_05335_));
 NAND2x1_ASAP7_75t_R _27736_ (.A(_05333_),
    .B(_05335_),
    .Y(_05336_));
 AOI21x1_ASAP7_75t_R _27737_ (.A1(_05103_),
    .A2(_05336_),
    .B(_05122_),
    .Y(_05337_));
 OAI21x1_ASAP7_75t_R _27738_ (.A1(_05324_),
    .A2(_05330_),
    .B(_05337_),
    .Y(_05338_));
 AND2x2_ASAP7_75t_L _27739_ (.A(_05248_),
    .B(_05097_),
    .Y(_05339_));
 NOR2x1_ASAP7_75t_SL _27740_ (.A(_05074_),
    .B(_05071_),
    .Y(_05340_));
 AOI21x1_ASAP7_75t_R _27741_ (.A1(_05090_),
    .A2(_05340_),
    .B(_05103_),
    .Y(_05341_));
 NAND2x1_ASAP7_75t_SL _27742_ (.A(_05184_),
    .B(_05341_),
    .Y(_05342_));
 AOI21x1_ASAP7_75t_R _27743_ (.A1(_05325_),
    .A2(_05227_),
    .B(_05104_),
    .Y(_05343_));
 AOI21x1_ASAP7_75t_R _27744_ (.A1(_05322_),
    .A2(_05343_),
    .B(_05154_),
    .Y(_05344_));
 OAI21x1_ASAP7_75t_R _27745_ (.A1(_05339_),
    .A2(_05342_),
    .B(_05344_),
    .Y(_05345_));
 INVx1_ASAP7_75t_R _27746_ (.A(_01324_),
    .Y(_05346_));
 AO21x1_ASAP7_75t_R _27747_ (.A1(_05067_),
    .A2(_05062_),
    .B(_05346_),
    .Y(_05347_));
 AOI21x1_ASAP7_75t_R _27748_ (.A1(_01331_),
    .A2(_05074_),
    .B(_05080_),
    .Y(_05348_));
 AOI21x1_ASAP7_75t_R _27749_ (.A1(_05347_),
    .A2(_05348_),
    .B(_05103_),
    .Y(_05349_));
 NAND2x1_ASAP7_75t_R _27750_ (.A(_05349_),
    .B(_05279_),
    .Y(_05350_));
 OAI21x1_ASAP7_75t_R _27751_ (.A1(_05068_),
    .A2(_05143_),
    .B(_05215_),
    .Y(_05351_));
 NOR2x1_ASAP7_75t_L _27752_ (.A(_05104_),
    .B(_05139_),
    .Y(_05352_));
 AOI21x1_ASAP7_75t_SL _27753_ (.A1(_05351_),
    .A2(_05352_),
    .B(_05155_),
    .Y(_05353_));
 AOI21x1_ASAP7_75t_R _27754_ (.A1(_05350_),
    .A2(_05353_),
    .B(_05121_),
    .Y(_05354_));
 AOI21x1_ASAP7_75t_R _27755_ (.A1(_05345_),
    .A2(_05354_),
    .B(_05236_),
    .Y(_05355_));
 NAND2x1_ASAP7_75t_R _27756_ (.A(_05338_),
    .B(_05355_),
    .Y(_05356_));
 NAND2x1_ASAP7_75t_SL _27757_ (.A(_05319_),
    .B(_05356_),
    .Y(_00129_));
 NOR2x1_ASAP7_75t_R _27758_ (.A(_05071_),
    .B(_05262_),
    .Y(_05357_));
 OAI21x1_ASAP7_75t_SL _27760_ (.A1(_05193_),
    .A2(_05357_),
    .B(_05104_),
    .Y(_05359_));
 NAND2x1_ASAP7_75t_R _27761_ (.A(_01324_),
    .B(_01326_),
    .Y(_05360_));
 NAND2x1_ASAP7_75t_L _27762_ (.A(_05360_),
    .B(_05074_),
    .Y(_05361_));
 INVx1_ASAP7_75t_R _27763_ (.A(_05361_),
    .Y(_05362_));
 OA21x2_ASAP7_75t_SL _27764_ (.A1(_05223_),
    .A2(_05362_),
    .B(_05080_),
    .Y(_05363_));
 OAI21x1_ASAP7_75t_R _27765_ (.A1(_05086_),
    .A2(_05206_),
    .B(_05080_),
    .Y(_05364_));
 AOI21x1_ASAP7_75t_SL _27766_ (.A1(_05364_),
    .A2(_05243_),
    .B(_05154_),
    .Y(_05365_));
 OAI21x1_ASAP7_75t_SL _27767_ (.A1(_05359_),
    .A2(_05363_),
    .B(_05365_),
    .Y(_05366_));
 NAND2x1_ASAP7_75t_R _27768_ (.A(_01335_),
    .B(_05080_),
    .Y(_05367_));
 OAI21x1_ASAP7_75t_SL _27769_ (.A1(_05051_),
    .A2(_05245_),
    .B(_05090_),
    .Y(_05368_));
 NAND2x1_ASAP7_75t_SL _27770_ (.A(_05367_),
    .B(_05368_),
    .Y(_05369_));
 OA21x2_ASAP7_75t_R _27771_ (.A1(_05080_),
    .A2(_01340_),
    .B(_05104_),
    .Y(_05370_));
 AOI21x1_ASAP7_75t_SL _27772_ (.A1(_05074_),
    .A2(_05040_),
    .B(_05090_),
    .Y(_05371_));
 NAND2x1_ASAP7_75t_SL _27773_ (.A(_05179_),
    .B(_05371_),
    .Y(_05372_));
 AOI21x1_ASAP7_75t_SL _27774_ (.A1(_05370_),
    .A2(_05372_),
    .B(_05155_),
    .Y(_05373_));
 OAI21x1_ASAP7_75t_SL _27775_ (.A1(_05104_),
    .A2(_05369_),
    .B(_05373_),
    .Y(_05374_));
 AOI21x1_ASAP7_75t_SL _27776_ (.A1(_05366_),
    .A2(_05374_),
    .B(_05122_),
    .Y(_05375_));
 OA21x2_ASAP7_75t_R _27777_ (.A1(_05080_),
    .A2(_01336_),
    .B(_05103_),
    .Y(_05376_));
 OAI21x1_ASAP7_75t_R _27778_ (.A1(_05068_),
    .A2(_05179_),
    .B(_05248_),
    .Y(_05377_));
 AOI21x1_ASAP7_75t_SL _27779_ (.A1(_05376_),
    .A2(_05377_),
    .B(_05154_),
    .Y(_05378_));
 AOI21x1_ASAP7_75t_R _27780_ (.A1(_05112_),
    .A2(_05169_),
    .B(_05103_),
    .Y(_05379_));
 AO21x1_ASAP7_75t_R _27781_ (.A1(_05245_),
    .A2(_05171_),
    .B(_05090_),
    .Y(_05380_));
 NAND2x1_ASAP7_75t_SL _27782_ (.A(_05379_),
    .B(_05380_),
    .Y(_05381_));
 NAND2x1_ASAP7_75t_SL _27783_ (.A(_05378_),
    .B(_05381_),
    .Y(_05382_));
 INVx1_ASAP7_75t_R _27784_ (.A(_05112_),
    .Y(_05383_));
 NAND2x1_ASAP7_75t_R _27785_ (.A(_05080_),
    .B(_05221_),
    .Y(_05384_));
 NOR2x1_ASAP7_75t_R _27786_ (.A(_05383_),
    .B(_05384_),
    .Y(_05385_));
 AND2x2_ASAP7_75t_R _27787_ (.A(_05169_),
    .B(_05164_),
    .Y(_05386_));
 OAI21x1_ASAP7_75t_SL _27788_ (.A1(_05385_),
    .A2(_05386_),
    .B(_05104_),
    .Y(_05387_));
 NAND2x1_ASAP7_75t_R _27789_ (.A(_01338_),
    .B(_05090_),
    .Y(_05388_));
 AOI21x1_ASAP7_75t_SL _27790_ (.A1(_05226_),
    .A2(_05371_),
    .B(_05104_),
    .Y(_05389_));
 AOI21x1_ASAP7_75t_SL _27791_ (.A1(_05388_),
    .A2(_05389_),
    .B(_05155_),
    .Y(_05390_));
 NAND2x1_ASAP7_75t_SL _27792_ (.A(_05387_),
    .B(_05390_),
    .Y(_05391_));
 AOI21x1_ASAP7_75t_SL _27794_ (.A1(_05382_),
    .A2(_05391_),
    .B(_05121_),
    .Y(_05393_));
 OAI21x1_ASAP7_75t_SL _27795_ (.A1(_05375_),
    .A2(_05393_),
    .B(_05236_),
    .Y(_05394_));
 AO21x1_ASAP7_75t_SL _27796_ (.A1(_05067_),
    .A2(_05062_),
    .B(_05133_),
    .Y(_05395_));
 AOI21x1_ASAP7_75t_SL _27797_ (.A1(_05395_),
    .A2(_05291_),
    .B(_05090_),
    .Y(_05396_));
 NOR2x1_ASAP7_75t_SL _27798_ (.A(_05080_),
    .B(_05208_),
    .Y(_05397_));
 AND2x2_ASAP7_75t_SL _27799_ (.A(_05397_),
    .B(_05130_),
    .Y(_05398_));
 OAI21x1_ASAP7_75t_SL _27800_ (.A1(_05396_),
    .A2(_05398_),
    .B(_05104_),
    .Y(_05399_));
 AOI21x1_ASAP7_75t_R _27801_ (.A1(_01326_),
    .A2(_05068_),
    .B(_05090_),
    .Y(_05400_));
 NAND2x1_ASAP7_75t_SL _27802_ (.A(_05271_),
    .B(_05400_),
    .Y(_05401_));
 NAND2x1_ASAP7_75t_R _27803_ (.A(_05134_),
    .B(_05130_),
    .Y(_05402_));
 AOI21x1_ASAP7_75t_SL _27804_ (.A1(_05090_),
    .A2(_05402_),
    .B(_05104_),
    .Y(_05403_));
 AOI21x1_ASAP7_75t_SL _27805_ (.A1(_05401_),
    .A2(_05403_),
    .B(_05155_),
    .Y(_05404_));
 NAND2x1_ASAP7_75t_SL _27806_ (.A(_05399_),
    .B(_05404_),
    .Y(_05405_));
 OAI21x1_ASAP7_75t_SL _27807_ (.A1(_05247_),
    .A2(_05206_),
    .B(_05080_),
    .Y(_05406_));
 NOR2x1_ASAP7_75t_SL _27808_ (.A(_05080_),
    .B(_05181_),
    .Y(_05407_));
 NAND2x1_ASAP7_75t_SL _27809_ (.A(_05291_),
    .B(_05407_),
    .Y(_05408_));
 AOI21x1_ASAP7_75t_SL _27810_ (.A1(_05406_),
    .A2(_05408_),
    .B(_05104_),
    .Y(_05409_));
 AOI21x1_ASAP7_75t_R _27811_ (.A1(_05072_),
    .A2(_05073_),
    .B(_01329_),
    .Y(_05410_));
 AOI211x1_ASAP7_75t_SL _27812_ (.A1(_01321_),
    .A2(_05068_),
    .B(_05090_),
    .C(_05410_),
    .Y(_05411_));
 OAI21x1_ASAP7_75t_R _27813_ (.A1(_05068_),
    .A2(_05071_),
    .B(_05090_),
    .Y(_05412_));
 OAI21x1_ASAP7_75t_SL _27814_ (.A1(_05208_),
    .A2(_05412_),
    .B(_05104_),
    .Y(_05413_));
 NOR2x1_ASAP7_75t_SL _27815_ (.A(_05411_),
    .B(_05413_),
    .Y(_05414_));
 OAI21x1_ASAP7_75t_SL _27816_ (.A1(_05409_),
    .A2(_05414_),
    .B(_05155_),
    .Y(_05415_));
 AOI21x1_ASAP7_75t_SL _27817_ (.A1(_05405_),
    .A2(_05415_),
    .B(_05121_),
    .Y(_05416_));
 INVx1_ASAP7_75t_SL _27818_ (.A(_05170_),
    .Y(_05417_));
 NOR3x1_ASAP7_75t_SL _27819_ (.A(_05088_),
    .B(_05090_),
    .C(_05086_),
    .Y(_05418_));
 NOR2x1_ASAP7_75t_SL _27820_ (.A(_05417_),
    .B(_05418_),
    .Y(_05419_));
 NOR2x1_ASAP7_75t_L _27821_ (.A(_05080_),
    .B(_05159_),
    .Y(_05420_));
 NOR2x1_ASAP7_75t_R _27822_ (.A(_05103_),
    .B(_05272_),
    .Y(_05421_));
 AOI21x1_ASAP7_75t_SL _27823_ (.A1(_05420_),
    .A2(_05421_),
    .B(_05155_),
    .Y(_05422_));
 OAI21x1_ASAP7_75t_SL _27824_ (.A1(_05103_),
    .A2(_05372_),
    .B(_05422_),
    .Y(_05423_));
 NOR2x1_ASAP7_75t_SL _27825_ (.A(_05419_),
    .B(_05423_),
    .Y(_05424_));
 OAI21x1_ASAP7_75t_R _27826_ (.A1(_05068_),
    .A2(_05071_),
    .B(_05080_),
    .Y(_05425_));
 NOR2x1_ASAP7_75t_SL _27827_ (.A(_05093_),
    .B(_05425_),
    .Y(_05426_));
 OAI21x1_ASAP7_75t_R _27828_ (.A1(_05074_),
    .A2(_05040_),
    .B(_05090_),
    .Y(_05427_));
 OAI21x1_ASAP7_75t_SL _27829_ (.A1(_05206_),
    .A2(_05427_),
    .B(_05104_),
    .Y(_05428_));
 OAI21x1_ASAP7_75t_SL _27830_ (.A1(_05426_),
    .A2(_05428_),
    .B(_05155_),
    .Y(_05429_));
 NOR2x1_ASAP7_75t_R _27831_ (.A(_01331_),
    .B(_05068_),
    .Y(_05430_));
 OAI21x1_ASAP7_75t_SL _27832_ (.A1(_05430_),
    .A2(_05223_),
    .B(_05080_),
    .Y(_05431_));
 AOI21x1_ASAP7_75t_SL _27833_ (.A1(_05368_),
    .A2(_05431_),
    .B(_05104_),
    .Y(_05432_));
 OAI21x1_ASAP7_75t_SL _27834_ (.A1(_05429_),
    .A2(_05432_),
    .B(_05121_),
    .Y(_05433_));
 NOR2x1_ASAP7_75t_SL _27835_ (.A(_05424_),
    .B(_05433_),
    .Y(_05434_));
 OAI21x1_ASAP7_75t_SL _27836_ (.A1(_05416_),
    .A2(_05434_),
    .B(_05202_),
    .Y(_05435_));
 NAND2x1_ASAP7_75t_SL _27837_ (.A(_05394_),
    .B(_05435_),
    .Y(_00130_));
 AO21x1_ASAP7_75t_R _27838_ (.A1(_05080_),
    .A2(_05074_),
    .B(_05104_),
    .Y(_05436_));
 AO21x1_ASAP7_75t_R _27839_ (.A1(_05171_),
    .A2(_05179_),
    .B(_05436_),
    .Y(_05437_));
 NAND2x1p5_ASAP7_75t_L _27840_ (.A(_05207_),
    .B(_05407_),
    .Y(_05438_));
 NAND2x1_ASAP7_75t_R _27841_ (.A(_05438_),
    .B(_05274_),
    .Y(_05439_));
 AOI21x1_ASAP7_75t_R _27842_ (.A1(_05437_),
    .A2(_05439_),
    .B(_05155_),
    .Y(_05440_));
 OAI21x1_ASAP7_75t_R _27843_ (.A1(_05264_),
    .A2(_05384_),
    .B(_05103_),
    .Y(_05441_));
 NOR2x1_ASAP7_75t_SL _27844_ (.A(_05114_),
    .B(_05327_),
    .Y(_05442_));
 NOR2x1_ASAP7_75t_SL _27845_ (.A(_05441_),
    .B(_05442_),
    .Y(_05443_));
 AND3x1_ASAP7_75t_L _27846_ (.A(_05090_),
    .B(_05173_),
    .C(_05282_),
    .Y(_05444_));
 OAI21x1_ASAP7_75t_R _27847_ (.A1(_05051_),
    .A2(_01321_),
    .B(_05080_),
    .Y(_05445_));
 OAI21x1_ASAP7_75t_R _27848_ (.A1(_05340_),
    .A2(_05445_),
    .B(_05104_),
    .Y(_05446_));
 OAI21x1_ASAP7_75t_R _27849_ (.A1(_05444_),
    .A2(_05446_),
    .B(_05155_),
    .Y(_05447_));
 OAI21x1_ASAP7_75t_SL _27850_ (.A1(_05447_),
    .A2(_05443_),
    .B(_05236_),
    .Y(_05448_));
 NOR2x1_ASAP7_75t_L _27851_ (.A(_05440_),
    .B(_05448_),
    .Y(_05449_));
 NAND2x1_ASAP7_75t_SL _27852_ (.A(_05300_),
    .B(_05106_),
    .Y(_05450_));
 NAND2x1_ASAP7_75t_R _27853_ (.A(_05071_),
    .B(_05298_),
    .Y(_05451_));
 AOI21x1_ASAP7_75t_R _27854_ (.A1(_05080_),
    .A2(_05410_),
    .B(_05103_),
    .Y(_05452_));
 OAI21x1_ASAP7_75t_R _27855_ (.A1(_05206_),
    .A2(_05208_),
    .B(_05090_),
    .Y(_05453_));
 NAND3x1_ASAP7_75t_R _27856_ (.A(_05451_),
    .B(_05452_),
    .C(_05453_),
    .Y(_05454_));
 AOI21x1_ASAP7_75t_R _27857_ (.A1(_05450_),
    .A2(_05454_),
    .B(_05154_),
    .Y(_05455_));
 NAND2x1_ASAP7_75t_R _27858_ (.A(_05154_),
    .B(_05413_),
    .Y(_05456_));
 AO21x1_ASAP7_75t_R _27859_ (.A1(_05067_),
    .A2(_05062_),
    .B(_01329_),
    .Y(_05457_));
 AO21x1_ASAP7_75t_R _27860_ (.A1(_05361_),
    .A2(_05457_),
    .B(_05090_),
    .Y(_05458_));
 AOI21x1_ASAP7_75t_R _27861_ (.A1(_05458_),
    .A2(_05333_),
    .B(_05104_),
    .Y(_05459_));
 OAI21x1_ASAP7_75t_R _27862_ (.A1(_05456_),
    .A2(_05459_),
    .B(_05202_),
    .Y(_05460_));
 OAI21x1_ASAP7_75t_R _27863_ (.A1(_05455_),
    .A2(_05460_),
    .B(_05122_),
    .Y(_05461_));
 NOR2x1_ASAP7_75t_SL _27864_ (.A(_05449_),
    .B(_05461_),
    .Y(_05462_));
 NAND2x1_ASAP7_75t_R _27865_ (.A(_05262_),
    .B(_05332_),
    .Y(_05463_));
 INVx2_ASAP7_75t_SL _27866_ (.A(_05247_),
    .Y(_05464_));
 OA21x2_ASAP7_75t_SL _27867_ (.A1(_05464_),
    .A2(_05090_),
    .B(_05154_),
    .Y(_05465_));
 AOI21x1_ASAP7_75t_R _27868_ (.A1(_05090_),
    .A2(_05138_),
    .B(_05154_),
    .Y(_05466_));
 AOI21x1_ASAP7_75t_R _27869_ (.A1(_05463_),
    .A2(_05465_),
    .B(_05466_),
    .Y(_05467_));
 OAI21x1_ASAP7_75t_R _27870_ (.A1(_05187_),
    .A2(_05467_),
    .B(_05202_),
    .Y(_05468_));
 NAND2x1_ASAP7_75t_R _27871_ (.A(_05080_),
    .B(_05410_),
    .Y(_05469_));
 NAND3x1_ASAP7_75t_R _27872_ (.A(_05408_),
    .B(_05155_),
    .C(_05469_),
    .Y(_05470_));
 NAND2x1_ASAP7_75t_L _27873_ (.A(_05282_),
    .B(_05215_),
    .Y(_05471_));
 INVx2_ASAP7_75t_R _27874_ (.A(_05272_),
    .Y(_05472_));
 OA21x2_ASAP7_75t_R _27875_ (.A1(_05068_),
    .A2(_05360_),
    .B(_05080_),
    .Y(_05473_));
 AOI21x1_ASAP7_75t_R _27876_ (.A1(_05472_),
    .A2(_05473_),
    .B(_05155_),
    .Y(_05474_));
 NAND2x1_ASAP7_75t_SL _27877_ (.A(_05471_),
    .B(_05474_),
    .Y(_05475_));
 AOI21x1_ASAP7_75t_R _27878_ (.A1(_05470_),
    .A2(_05475_),
    .B(_05104_),
    .Y(_05476_));
 OAI21x1_ASAP7_75t_SL _27879_ (.A1(_05476_),
    .A2(_05468_),
    .B(_05121_),
    .Y(_05477_));
 AND2x2_ASAP7_75t_R _27880_ (.A(_05286_),
    .B(_05221_),
    .Y(_05478_));
 AO21x1_ASAP7_75t_SL _27881_ (.A1(_05287_),
    .A2(_05248_),
    .B(_05154_),
    .Y(_05479_));
 NOR2x1_ASAP7_75t_L _27882_ (.A(_05478_),
    .B(_05479_),
    .Y(_05480_));
 AO21x1_ASAP7_75t_SL _27883_ (.A1(_05465_),
    .A2(_05321_),
    .B(_05103_),
    .Y(_05481_));
 OAI21x1_ASAP7_75t_SL _27884_ (.A1(_05481_),
    .A2(_05480_),
    .B(_05236_),
    .Y(_05482_));
 NAND2x1_ASAP7_75t_SL _27885_ (.A(_05179_),
    .B(_05227_),
    .Y(_05483_));
 NAND2x1_ASAP7_75t_R _27886_ (.A(_05252_),
    .B(_05139_),
    .Y(_05484_));
 AOI21x1_ASAP7_75t_R _27887_ (.A1(_05483_),
    .A2(_05484_),
    .B(_05155_),
    .Y(_05485_));
 AOI21x1_ASAP7_75t_R _27888_ (.A1(_05068_),
    .A2(_01321_),
    .B(_05080_),
    .Y(_05486_));
 AOI22x1_ASAP7_75t_R _27889_ (.A1(_05486_),
    .A2(_05207_),
    .B1(_05400_),
    .B2(_05260_),
    .Y(_05487_));
 OAI21x1_ASAP7_75t_R _27890_ (.A1(_05154_),
    .A2(_05487_),
    .B(_05103_),
    .Y(_05488_));
 NOR2x1_ASAP7_75t_SL _27891_ (.A(_05485_),
    .B(_05488_),
    .Y(_05489_));
 NOR2x1_ASAP7_75t_SL _27892_ (.A(_05482_),
    .B(_05489_),
    .Y(_05490_));
 NOR2x1_ASAP7_75t_SL _27893_ (.A(_05477_),
    .B(_05490_),
    .Y(_05491_));
 NOR2x1_ASAP7_75t_SL _27894_ (.A(_05462_),
    .B(_05491_),
    .Y(_00131_));
 AO21x1_ASAP7_75t_SL _27895_ (.A1(_05389_),
    .A2(_05321_),
    .B(_05155_),
    .Y(_05492_));
 NAND2x1_ASAP7_75t_SL _27896_ (.A(_05179_),
    .B(_05486_),
    .Y(_05493_));
 NAND2x1_ASAP7_75t_R _27897_ (.A(_05164_),
    .B(_05371_),
    .Y(_05494_));
 AOI21x1_ASAP7_75t_R _27898_ (.A1(_05493_),
    .A2(_05494_),
    .B(_05103_),
    .Y(_05495_));
 AOI21x1_ASAP7_75t_R _27899_ (.A1(_05171_),
    .A2(_05252_),
    .B(_05090_),
    .Y(_05496_));
 AO21x1_ASAP7_75t_R _27900_ (.A1(_05211_),
    .A2(_05325_),
    .B(_05104_),
    .Y(_05497_));
 NAND2x1_ASAP7_75t_R _27901_ (.A(_05104_),
    .B(_05254_),
    .Y(_05498_));
 OA21x2_ASAP7_75t_R _27902_ (.A1(_05498_),
    .A2(_05182_),
    .B(_05155_),
    .Y(_05499_));
 OAI21x1_ASAP7_75t_R _27903_ (.A1(_05496_),
    .A2(_05497_),
    .B(_05499_),
    .Y(_05500_));
 OAI21x1_ASAP7_75t_R _27904_ (.A1(_05492_),
    .A2(_05495_),
    .B(_05500_),
    .Y(_05501_));
 NOR2x1_ASAP7_75t_R _27905_ (.A(_05121_),
    .B(_05501_),
    .Y(_05502_));
 AND2x2_ASAP7_75t_R _27906_ (.A(_05420_),
    .B(_05472_),
    .Y(_05503_));
 OAI21x1_ASAP7_75t_R _27907_ (.A1(_05051_),
    .A2(_01321_),
    .B(_05074_),
    .Y(_05504_));
 AOI21x1_ASAP7_75t_R _27909_ (.A1(_05245_),
    .A2(_05504_),
    .B(_05090_),
    .Y(_05506_));
 OAI21x1_ASAP7_75t_R _27910_ (.A1(_05503_),
    .A2(_05506_),
    .B(_05104_),
    .Y(_05507_));
 OAI21x1_ASAP7_75t_R _27911_ (.A1(_05080_),
    .A2(_05504_),
    .B(_05146_),
    .Y(_05508_));
 AND3x1_ASAP7_75t_R _27912_ (.A(_05252_),
    .B(_05080_),
    .C(_05097_),
    .Y(_05509_));
 OAI21x1_ASAP7_75t_R _27913_ (.A1(_05508_),
    .A2(_05509_),
    .B(_05103_),
    .Y(_05510_));
 AOI21x1_ASAP7_75t_R _27914_ (.A1(_05507_),
    .A2(_05510_),
    .B(_05155_),
    .Y(_05511_));
 NAND2x1_ASAP7_75t_R _27915_ (.A(_05464_),
    .B(_05348_),
    .Y(_05512_));
 AND3x1_ASAP7_75t_R _27916_ (.A(_05183_),
    .B(_05103_),
    .C(_05512_),
    .Y(_05513_));
 NOR2x1p5_ASAP7_75t_L _27917_ (.A(_05090_),
    .B(_05112_),
    .Y(_05514_));
 INVx1_ASAP7_75t_R _27918_ (.A(_05514_),
    .Y(_05515_));
 AO31x2_ASAP7_75t_R _27919_ (.A1(_05452_),
    .A2(_05515_),
    .A3(_05135_),
    .B(_05154_),
    .Y(_05516_));
 OAI21x1_ASAP7_75t_R _27920_ (.A1(_05513_),
    .A2(_05516_),
    .B(_05121_),
    .Y(_05517_));
 OAI21x1_ASAP7_75t_R _27921_ (.A1(_05511_),
    .A2(_05517_),
    .B(_05236_),
    .Y(_05518_));
 NAND2x1_ASAP7_75t_R _27922_ (.A(_05097_),
    .B(_05320_),
    .Y(_05519_));
 AOI21x1_ASAP7_75t_R _27923_ (.A1(_05252_),
    .A2(_05160_),
    .B(_05103_),
    .Y(_05520_));
 NAND2x1_ASAP7_75t_R _27924_ (.A(_05519_),
    .B(_05520_),
    .Y(_05521_));
 AND2x2_ASAP7_75t_R _27925_ (.A(_05297_),
    .B(_05103_),
    .Y(_05522_));
 NAND2x1_ASAP7_75t_R _27926_ (.A(_05472_),
    .B(_05227_),
    .Y(_05523_));
 AOI21x1_ASAP7_75t_SL _27927_ (.A1(_05522_),
    .A2(_05523_),
    .B(_05121_),
    .Y(_05524_));
 AOI21x1_ASAP7_75t_R _27928_ (.A1(_05521_),
    .A2(_05524_),
    .B(_05155_),
    .Y(_05525_));
 NAND2x1_ASAP7_75t_R _27929_ (.A(_05171_),
    .B(_05182_),
    .Y(_05526_));
 AOI21x1_ASAP7_75t_R _27930_ (.A1(_05526_),
    .A2(_05493_),
    .B(_05103_),
    .Y(_05527_));
 NAND2x1_ASAP7_75t_R _27931_ (.A(_05229_),
    .B(_05231_),
    .Y(_05528_));
 AOI21x1_ASAP7_75t_R _27932_ (.A1(_05167_),
    .A2(_05528_),
    .B(_05104_),
    .Y(_05529_));
 OAI21x1_ASAP7_75t_R _27933_ (.A1(_05527_),
    .A2(_05529_),
    .B(_05121_),
    .Y(_05530_));
 NAND2x1_ASAP7_75t_SL _27934_ (.A(_05525_),
    .B(_05530_),
    .Y(_05531_));
 AOI21x1_ASAP7_75t_R _27935_ (.A1(_05112_),
    .A2(_05420_),
    .B(_05104_),
    .Y(_05532_));
 NAND2x1_ASAP7_75t_R _27936_ (.A(_05532_),
    .B(_05144_),
    .Y(_05533_));
 AOI21x1_ASAP7_75t_R _27937_ (.A1(_05090_),
    .A2(_05347_),
    .B(_05103_),
    .Y(_05534_));
 OAI21x1_ASAP7_75t_R _27938_ (.A1(_05071_),
    .A2(_05245_),
    .B(_05080_),
    .Y(_05535_));
 AOI21x1_ASAP7_75t_R _27939_ (.A1(_05534_),
    .A2(_05535_),
    .B(_05121_),
    .Y(_05536_));
 AOI21x1_ASAP7_75t_R _27940_ (.A1(_05533_),
    .A2(_05536_),
    .B(_05154_),
    .Y(_05537_));
 INVx1_ASAP7_75t_R _27941_ (.A(_01330_),
    .Y(_05538_));
 AOI211x1_ASAP7_75t_R _27942_ (.A1(_05538_),
    .A2(_05090_),
    .B(_05514_),
    .C(_05104_),
    .Y(_05539_));
 NAND2x1_ASAP7_75t_L _27943_ (.A(_05271_),
    .B(_05182_),
    .Y(_05540_));
 NAND2x1_ASAP7_75t_R _27944_ (.A(_05090_),
    .B(_05088_),
    .Y(_05541_));
 AOI21x1_ASAP7_75t_R _27945_ (.A1(_05540_),
    .A2(_05541_),
    .B(_05103_),
    .Y(_05542_));
 OAI21x1_ASAP7_75t_R _27946_ (.A1(_05539_),
    .A2(_05542_),
    .B(_05121_),
    .Y(_05543_));
 AOI21x1_ASAP7_75t_R _27947_ (.A1(_05537_),
    .A2(_05543_),
    .B(_05236_),
    .Y(_05544_));
 NAND2x1_ASAP7_75t_SL _27948_ (.A(_05531_),
    .B(_05544_),
    .Y(_05545_));
 OAI21x1_ASAP7_75t_SL _27949_ (.A1(_05502_),
    .A2(_05518_),
    .B(_05545_),
    .Y(_00132_));
 OR2x2_ASAP7_75t_SL _27950_ (.A(_05473_),
    .B(_05104_),
    .Y(_05546_));
 NOR2x1_ASAP7_75t_SL _27951_ (.A(_05357_),
    .B(_05368_),
    .Y(_05547_));
 OA21x2_ASAP7_75t_SL _27952_ (.A1(_05309_),
    .A2(_05273_),
    .B(_05155_),
    .Y(_05548_));
 OAI21x1_ASAP7_75t_SL _27953_ (.A1(_05546_),
    .A2(_05547_),
    .B(_05548_),
    .Y(_05549_));
 OA21x2_ASAP7_75t_SL _27954_ (.A1(_05090_),
    .A2(_05172_),
    .B(_05103_),
    .Y(_05550_));
 NOR2x1_ASAP7_75t_SL _27955_ (.A(_05080_),
    .B(_05051_),
    .Y(_05551_));
 NOR2x1_ASAP7_75t_SL _27956_ (.A(_05551_),
    .B(_05169_),
    .Y(_05552_));
 AOI21x1_ASAP7_75t_SL _27957_ (.A1(_05550_),
    .A2(_05552_),
    .B(_05155_),
    .Y(_05553_));
 AO21x1_ASAP7_75t_SL _27958_ (.A1(_05282_),
    .A2(_05209_),
    .B(_05080_),
    .Y(_05554_));
 AO21x1_ASAP7_75t_SL _27959_ (.A1(_05207_),
    .A2(_05173_),
    .B(_05090_),
    .Y(_05555_));
 NAND3x1_ASAP7_75t_SL _27960_ (.A(_05554_),
    .B(_05555_),
    .C(_05104_),
    .Y(_05556_));
 AOI21x1_ASAP7_75t_SL _27961_ (.A1(_05553_),
    .A2(_05556_),
    .B(_05122_),
    .Y(_05557_));
 NAND2x1_ASAP7_75t_SL _27962_ (.A(_05549_),
    .B(_05557_),
    .Y(_05558_));
 OA21x2_ASAP7_75t_SL _27963_ (.A1(_05071_),
    .A2(_05090_),
    .B(_05103_),
    .Y(_05559_));
 AOI21x1_ASAP7_75t_SL _27964_ (.A1(_05559_),
    .A2(_05228_),
    .B(_05154_),
    .Y(_05560_));
 NOR2x1_ASAP7_75t_SL _27965_ (.A(_05051_),
    .B(_05245_),
    .Y(_05561_));
 AOI21x1_ASAP7_75t_SL _27966_ (.A1(_05271_),
    .A2(_05407_),
    .B(_05103_),
    .Y(_05562_));
 OAI21x1_ASAP7_75t_SL _27967_ (.A1(_05284_),
    .A2(_05561_),
    .B(_05562_),
    .Y(_05563_));
 AOI21x1_ASAP7_75t_SL _27968_ (.A1(_05560_),
    .A2(_05563_),
    .B(_05121_),
    .Y(_05564_));
 NAND2x1_ASAP7_75t_SL _27969_ (.A(_05103_),
    .B(_05144_),
    .Y(_05565_));
 AND2x2_ASAP7_75t_SL _27970_ (.A(_05211_),
    .B(_05395_),
    .Y(_05566_));
 OA21x2_ASAP7_75t_SL _27971_ (.A1(_05173_),
    .A2(_05090_),
    .B(_05104_),
    .Y(_05567_));
 OAI21x1_ASAP7_75t_SL _27972_ (.A1(_05551_),
    .A2(_05169_),
    .B(_05472_),
    .Y(_05568_));
 AOI21x1_ASAP7_75t_SL _27973_ (.A1(_05567_),
    .A2(_05568_),
    .B(_05155_),
    .Y(_05569_));
 OAI21x1_ASAP7_75t_SL _27974_ (.A1(_05565_),
    .A2(_05566_),
    .B(_05569_),
    .Y(_05570_));
 AOI21x1_ASAP7_75t_SL _27975_ (.A1(_05564_),
    .A2(_05570_),
    .B(_05236_),
    .Y(_05571_));
 NAND2x1_ASAP7_75t_SL _27976_ (.A(_05558_),
    .B(_05571_),
    .Y(_05572_));
 NOR2x1_ASAP7_75t_SL _27977_ (.A(_05103_),
    .B(_05420_),
    .Y(_05573_));
 AOI21x1_ASAP7_75t_SL _27978_ (.A1(_05573_),
    .A2(_05299_),
    .B(_05155_),
    .Y(_05574_));
 NOR2x1_ASAP7_75t_R _27979_ (.A(_05074_),
    .B(_05051_),
    .Y(_05575_));
 OAI21x1_ASAP7_75t_SL _27980_ (.A1(_05410_),
    .A2(_05575_),
    .B(_05080_),
    .Y(_05576_));
 AO21x1_ASAP7_75t_SL _27981_ (.A1(_05090_),
    .A2(_05282_),
    .B(_05104_),
    .Y(_05577_));
 INVx1_ASAP7_75t_SL _27982_ (.A(_05577_),
    .Y(_05578_));
 NAND2x1_ASAP7_75t_SL _27983_ (.A(_05576_),
    .B(_05578_),
    .Y(_05579_));
 AOI21x1_ASAP7_75t_SL _27984_ (.A1(_05574_),
    .A2(_05579_),
    .B(_05121_),
    .Y(_05580_));
 NOR2x1_ASAP7_75t_R _27985_ (.A(_01326_),
    .B(_05090_),
    .Y(_05581_));
 AOI211x1_ASAP7_75t_SL _27986_ (.A1(_05162_),
    .A2(_05080_),
    .B(_05103_),
    .C(_05581_),
    .Y(_05582_));
 AO21x1_ASAP7_75t_SL _27987_ (.A1(_05504_),
    .A2(_05457_),
    .B(_05080_),
    .Y(_05583_));
 NAND2x1_ASAP7_75t_SL _27988_ (.A(_05582_),
    .B(_05583_),
    .Y(_05584_));
 AO21x1_ASAP7_75t_SL _27989_ (.A1(_05276_),
    .A2(_05209_),
    .B(_05090_),
    .Y(_05585_));
 AOI21x1_ASAP7_75t_SL _27990_ (.A1(_05585_),
    .A2(_05257_),
    .B(_05154_),
    .Y(_05586_));
 NAND2x1_ASAP7_75t_SL _27991_ (.A(_05584_),
    .B(_05586_),
    .Y(_05587_));
 AOI21x1_ASAP7_75t_SL _27992_ (.A1(_05580_),
    .A2(_05587_),
    .B(_05202_),
    .Y(_05588_));
 AOI211x1_ASAP7_75t_SL _27993_ (.A1(_05139_),
    .A2(_05164_),
    .B(_05397_),
    .C(_05155_),
    .Y(_05589_));
 OA21x2_ASAP7_75t_SL _27994_ (.A1(_05040_),
    .A2(_05090_),
    .B(_05155_),
    .Y(_05590_));
 AO21x1_ASAP7_75t_SL _27995_ (.A1(_05590_),
    .A2(_05493_),
    .B(_05104_),
    .Y(_05591_));
 NOR2x1_ASAP7_75t_SL _27996_ (.A(_05589_),
    .B(_05591_),
    .Y(_05592_));
 OA21x2_ASAP7_75t_SL _27997_ (.A1(_05074_),
    .A2(_05346_),
    .B(_05090_),
    .Y(_05593_));
 AOI21x1_ASAP7_75t_SL _27998_ (.A1(_05262_),
    .A2(_05593_),
    .B(_05514_),
    .Y(_05594_));
 OAI21x1_ASAP7_75t_SL _27999_ (.A1(_05155_),
    .A2(_05594_),
    .B(_05104_),
    .Y(_05595_));
 NAND2x1_ASAP7_75t_SL _28000_ (.A(_05080_),
    .B(_05173_),
    .Y(_05596_));
 AOI21x1_ASAP7_75t_SL _28001_ (.A1(_05143_),
    .A2(_05215_),
    .B(_05154_),
    .Y(_05597_));
 OA21x2_ASAP7_75t_SL _28002_ (.A1(_05327_),
    .A2(_05596_),
    .B(_05597_),
    .Y(_05598_));
 NOR2x1_ASAP7_75t_SL _28003_ (.A(_05595_),
    .B(_05598_),
    .Y(_05599_));
 OAI21x1_ASAP7_75t_SL _28004_ (.A1(_05592_),
    .A2(_05599_),
    .B(_05121_),
    .Y(_05600_));
 NAND2x1_ASAP7_75t_SL _28005_ (.A(_05588_),
    .B(_05600_),
    .Y(_05601_));
 NAND2x1_ASAP7_75t_SL _28006_ (.A(_05572_),
    .B(_05601_),
    .Y(_00133_));
 OA21x2_ASAP7_75t_R _28007_ (.A1(_05282_),
    .A2(_05080_),
    .B(_05104_),
    .Y(_05602_));
 AOI21x1_ASAP7_75t_R _28008_ (.A1(_05602_),
    .A2(_05369_),
    .B(_05154_),
    .Y(_05603_));
 OA21x2_ASAP7_75t_R _28009_ (.A1(_05264_),
    .A2(_05263_),
    .B(_05080_),
    .Y(_05604_));
 AOI21x1_ASAP7_75t_R _28010_ (.A1(_05090_),
    .A2(_05206_),
    .B(_05104_),
    .Y(_05605_));
 OAI21x1_ASAP7_75t_R _28011_ (.A1(_05593_),
    .A2(_05604_),
    .B(_05605_),
    .Y(_05606_));
 NAND2x1_ASAP7_75t_SL _28012_ (.A(_05603_),
    .B(_05606_),
    .Y(_05607_));
 OAI21x1_ASAP7_75t_R _28013_ (.A1(_05051_),
    .A2(_05297_),
    .B(_05103_),
    .Y(_05608_));
 AOI21x1_ASAP7_75t_R _28014_ (.A1(_05464_),
    .A2(_05361_),
    .B(_05080_),
    .Y(_05609_));
 AOI211x1_ASAP7_75t_R _28015_ (.A1(_05229_),
    .A2(_05231_),
    .B(_05608_),
    .C(_05609_),
    .Y(_05610_));
 NAND2x1_ASAP7_75t_R _28016_ (.A(_05179_),
    .B(_05312_),
    .Y(_05611_));
 AND3x1_ASAP7_75t_R _28017_ (.A(_05611_),
    .B(_05104_),
    .C(_05240_),
    .Y(_05612_));
 OAI21x1_ASAP7_75t_R _28018_ (.A1(_05610_),
    .A2(_05612_),
    .B(_05154_),
    .Y(_05613_));
 AOI21x1_ASAP7_75t_R _28019_ (.A1(_05607_),
    .A2(_05613_),
    .B(_05122_),
    .Y(_05614_));
 NAND2x1_ASAP7_75t_R _28020_ (.A(_05090_),
    .B(_05241_),
    .Y(_05615_));
 AO21x1_ASAP7_75t_R _28021_ (.A1(_05615_),
    .A2(_05469_),
    .B(_05154_),
    .Y(_05616_));
 NAND2x1_ASAP7_75t_R _28022_ (.A(_05154_),
    .B(_05171_),
    .Y(_05617_));
 NAND2x1_ASAP7_75t_R _28023_ (.A(_05080_),
    .B(_05093_),
    .Y(_05618_));
 OAI21x1_ASAP7_75t_R _28024_ (.A1(_05114_),
    .A2(_05617_),
    .B(_05618_),
    .Y(_05619_));
 AND3x1_ASAP7_75t_SL _28025_ (.A(_05402_),
    .B(_05080_),
    .C(_05154_),
    .Y(_05620_));
 NOR2x1_ASAP7_75t_R _28026_ (.A(_05619_),
    .B(_05620_),
    .Y(_05621_));
 AOI21x1_ASAP7_75t_R _28027_ (.A1(_05616_),
    .A2(_05621_),
    .B(_05103_),
    .Y(_05622_));
 NAND2x1_ASAP7_75t_R _28028_ (.A(_01339_),
    .B(_01333_),
    .Y(_05623_));
 AO21x1_ASAP7_75t_R _28029_ (.A1(_05090_),
    .A2(_05623_),
    .B(_05154_),
    .Y(_05624_));
 AND3x1_ASAP7_75t_SL _28030_ (.A(_05179_),
    .B(_05080_),
    .C(_05252_),
    .Y(_05625_));
 OAI21x1_ASAP7_75t_R _28031_ (.A1(_05624_),
    .A2(_05625_),
    .B(_05103_),
    .Y(_05626_));
 AO21x1_ASAP7_75t_R _28032_ (.A1(_05162_),
    .A2(_05080_),
    .B(_05155_),
    .Y(_05627_));
 AND2x2_ASAP7_75t_R _28033_ (.A(_05407_),
    .B(_05260_),
    .Y(_05628_));
 AOI211x1_ASAP7_75t_R _28034_ (.A1(_05143_),
    .A2(_05298_),
    .B(_05627_),
    .C(_05628_),
    .Y(_05629_));
 OAI21x1_ASAP7_75t_R _28035_ (.A1(_05626_),
    .A2(_05629_),
    .B(_05122_),
    .Y(_05630_));
 OAI21x1_ASAP7_75t_R _28036_ (.A1(_05622_),
    .A2(_05630_),
    .B(_05236_),
    .Y(_05631_));
 AOI21x1_ASAP7_75t_R _28037_ (.A1(_01334_),
    .A2(_05080_),
    .B(_05104_),
    .Y(_05632_));
 NAND2x1_ASAP7_75t_R _28038_ (.A(_05271_),
    .B(_05407_),
    .Y(_05633_));
 AOI21x1_ASAP7_75t_R _28039_ (.A1(_05632_),
    .A2(_05633_),
    .B(_05154_),
    .Y(_05634_));
 AO21x1_ASAP7_75t_R _28040_ (.A1(_05282_),
    .A2(_05209_),
    .B(_05090_),
    .Y(_05635_));
 NAND2x1_ASAP7_75t_R _28041_ (.A(_05341_),
    .B(_05635_),
    .Y(_05636_));
 NAND2x1_ASAP7_75t_SL _28042_ (.A(_05634_),
    .B(_05636_),
    .Y(_05637_));
 NAND2x1_ASAP7_75t_R _28043_ (.A(_05271_),
    .B(_05396_),
    .Y(_05638_));
 AOI21x1_ASAP7_75t_R _28044_ (.A1(_05090_),
    .A2(_05192_),
    .B(_05103_),
    .Y(_05639_));
 AOI21x1_ASAP7_75t_R _28045_ (.A1(_05639_),
    .A2(_05540_),
    .B(_05155_),
    .Y(_05640_));
 OAI21x1_ASAP7_75t_R _28046_ (.A1(_05104_),
    .A2(_05638_),
    .B(_05640_),
    .Y(_05641_));
 AOI21x1_ASAP7_75t_R _28047_ (.A1(_05637_),
    .A2(_05641_),
    .B(_05122_),
    .Y(_05642_));
 AND2x2_ASAP7_75t_R _28048_ (.A(_05286_),
    .B(_05260_),
    .Y(_05643_));
 NAND2x1_ASAP7_75t_R _28049_ (.A(_05229_),
    .B(_05226_),
    .Y(_05644_));
 OAI21x1_ASAP7_75t_R _28050_ (.A1(_05090_),
    .A2(_05644_),
    .B(_05104_),
    .Y(_05645_));
 AO21x1_ASAP7_75t_R _28051_ (.A1(_05051_),
    .A2(_05080_),
    .B(_05040_),
    .Y(_05646_));
 NOR2x1_ASAP7_75t_R _28052_ (.A(_05104_),
    .B(_05340_),
    .Y(_05647_));
 AOI21x1_ASAP7_75t_R _28053_ (.A1(_05646_),
    .A2(_05647_),
    .B(_05154_),
    .Y(_05648_));
 OAI21x1_ASAP7_75t_R _28054_ (.A1(_05643_),
    .A2(_05645_),
    .B(_05648_),
    .Y(_05649_));
 OAI21x1_ASAP7_75t_R _28055_ (.A1(_05074_),
    .A2(_01321_),
    .B(_05080_),
    .Y(_05650_));
 NAND2x1_ASAP7_75t_R _28056_ (.A(_05650_),
    .B(_05212_),
    .Y(_05651_));
 AOI21x1_ASAP7_75t_R _28057_ (.A1(_05605_),
    .A2(_05576_),
    .B(_05155_),
    .Y(_05652_));
 NAND2x1_ASAP7_75t_SL _28058_ (.A(_05651_),
    .B(_05652_),
    .Y(_05653_));
 AOI21x1_ASAP7_75t_R _28059_ (.A1(_05649_),
    .A2(_05653_),
    .B(_05121_),
    .Y(_05654_));
 OAI21x1_ASAP7_75t_SL _28060_ (.A1(_05642_),
    .A2(_05654_),
    .B(_05202_),
    .Y(_05655_));
 OAI21x1_ASAP7_75t_SL _28061_ (.A1(_05614_),
    .A2(_05631_),
    .B(_05655_),
    .Y(_00134_));
 NOR2x1_ASAP7_75t_R _28062_ (.A(_01326_),
    .B(_05080_),
    .Y(_05656_));
 OAI21x1_ASAP7_75t_R _28063_ (.A1(_05656_),
    .A2(_05625_),
    .B(_05104_),
    .Y(_05657_));
 NOR2x1_ASAP7_75t_R _28064_ (.A(_05312_),
    .B(_05593_),
    .Y(_05658_));
 NAND2x1_ASAP7_75t_R _28065_ (.A(_05103_),
    .B(_05097_),
    .Y(_05659_));
 OA21x2_ASAP7_75t_R _28066_ (.A1(_05658_),
    .A2(_05659_),
    .B(_05154_),
    .Y(_05660_));
 NAND2x1_ASAP7_75t_R _28067_ (.A(_05657_),
    .B(_05660_),
    .Y(_05661_));
 NAND2x1_ASAP7_75t_R _28068_ (.A(_05143_),
    .B(_05169_),
    .Y(_05662_));
 AO21x1_ASAP7_75t_L _28069_ (.A1(_05458_),
    .A2(_05662_),
    .B(_05103_),
    .Y(_05663_));
 NOR2x1_ASAP7_75t_SL _28070_ (.A(_05241_),
    .B(_05223_),
    .Y(_05664_));
 NAND2x1_ASAP7_75t_R _28071_ (.A(_05090_),
    .B(_05664_),
    .Y(_05665_));
 OA21x2_ASAP7_75t_SL _28072_ (.A1(_05239_),
    .A2(_05284_),
    .B(_05103_),
    .Y(_05666_));
 AOI21x1_ASAP7_75t_R _28073_ (.A1(_05665_),
    .A2(_05666_),
    .B(_05154_),
    .Y(_05667_));
 NAND2x1_ASAP7_75t_L _28074_ (.A(_05663_),
    .B(_05667_),
    .Y(_05668_));
 AOI21x1_ASAP7_75t_R _28075_ (.A1(_05661_),
    .A2(_05668_),
    .B(_05202_),
    .Y(_05669_));
 NOR2x1_ASAP7_75t_R _28076_ (.A(_05104_),
    .B(_05348_),
    .Y(_05670_));
 AO21x1_ASAP7_75t_R _28077_ (.A1(_05670_),
    .A2(_05540_),
    .B(_05154_),
    .Y(_05671_));
 NAND2x1_ASAP7_75t_SL _28078_ (.A(_05341_),
    .B(_05541_),
    .Y(_05672_));
 NOR2x1_ASAP7_75t_R _28079_ (.A(_05090_),
    .B(_05664_),
    .Y(_05673_));
 NOR2x1_ASAP7_75t_R _28080_ (.A(_05672_),
    .B(_05673_),
    .Y(_05674_));
 OAI21x1_ASAP7_75t_SL _28081_ (.A1(_05671_),
    .A2(_05674_),
    .B(_05202_),
    .Y(_05675_));
 NAND2x1_ASAP7_75t_R _28082_ (.A(_05260_),
    .B(_05248_),
    .Y(_05676_));
 AO21x1_ASAP7_75t_SL _28083_ (.A1(_05676_),
    .A2(_05471_),
    .B(_05103_),
    .Y(_05677_));
 INVx1_ASAP7_75t_R _28084_ (.A(_05380_),
    .Y(_05678_));
 OAI21x1_ASAP7_75t_R _28085_ (.A1(_05628_),
    .A2(_05678_),
    .B(_05103_),
    .Y(_05679_));
 AOI21x1_ASAP7_75t_R _28086_ (.A1(_05677_),
    .A2(_05679_),
    .B(_05155_),
    .Y(_05680_));
 OAI21x1_ASAP7_75t_R _28087_ (.A1(_05675_),
    .A2(_05680_),
    .B(_05122_),
    .Y(_05681_));
 AND3x1_ASAP7_75t_L _28088_ (.A(_05464_),
    .B(_05207_),
    .C(_05080_),
    .Y(_05682_));
 AO21x1_ASAP7_75t_R _28089_ (.A1(_05215_),
    .A2(_05271_),
    .B(_05103_),
    .Y(_05683_));
 OAI21x1_ASAP7_75t_R _28090_ (.A1(_05410_),
    .A2(_05247_),
    .B(_05090_),
    .Y(_05684_));
 OA21x2_ASAP7_75t_R _28091_ (.A1(_05090_),
    .A2(_01339_),
    .B(_05103_),
    .Y(_05685_));
 AOI21x1_ASAP7_75t_R _28092_ (.A1(_05684_),
    .A2(_05685_),
    .B(_05155_),
    .Y(_05686_));
 OAI21x1_ASAP7_75t_R _28093_ (.A1(_05682_),
    .A2(_05683_),
    .B(_05686_),
    .Y(_05687_));
 OA21x2_ASAP7_75t_R _28094_ (.A1(_05090_),
    .A2(_05538_),
    .B(_05103_),
    .Y(_05688_));
 AOI21x1_ASAP7_75t_SL _28095_ (.A1(_05094_),
    .A2(_05688_),
    .B(_05154_),
    .Y(_05689_));
 NAND2x1_ASAP7_75t_R _28096_ (.A(_05179_),
    .B(_05320_),
    .Y(_05690_));
 NAND2x1_ASAP7_75t_R _28097_ (.A(_05690_),
    .B(_05520_),
    .Y(_05691_));
 AOI21x1_ASAP7_75t_R _28098_ (.A1(_05689_),
    .A2(_05691_),
    .B(_05202_),
    .Y(_05692_));
 AOI21x1_ASAP7_75t_R _28099_ (.A1(_05687_),
    .A2(_05692_),
    .B(_05122_),
    .Y(_05693_));
 OAI21x1_ASAP7_75t_R _28100_ (.A1(_05051_),
    .A2(_05262_),
    .B(_05080_),
    .Y(_05694_));
 NOR2x1_ASAP7_75t_R _28101_ (.A(_05551_),
    .B(_05320_),
    .Y(_05695_));
 AO21x1_ASAP7_75t_R _28102_ (.A1(_05206_),
    .A2(_05090_),
    .B(_05103_),
    .Y(_05696_));
 AOI21x1_ASAP7_75t_R _28103_ (.A1(_05694_),
    .A2(_05695_),
    .B(_05696_),
    .Y(_05697_));
 AOI21x1_ASAP7_75t_R _28104_ (.A1(_05074_),
    .A2(_05143_),
    .B(_05090_),
    .Y(_05698_));
 OAI21x1_ASAP7_75t_R _28105_ (.A1(_05698_),
    .A2(_05577_),
    .B(_05154_),
    .Y(_05699_));
 NOR2x1_ASAP7_75t_L _28106_ (.A(_05697_),
    .B(_05699_),
    .Y(_05700_));
 OAI21x1_ASAP7_75t_R _28107_ (.A1(_05551_),
    .A2(_05320_),
    .B(_05271_),
    .Y(_05701_));
 NAND2x1_ASAP7_75t_R _28108_ (.A(_05701_),
    .B(_05389_),
    .Y(_05702_));
 OAI21x1_ASAP7_75t_R _28109_ (.A1(_05551_),
    .A2(_05496_),
    .B(_05104_),
    .Y(_05703_));
 AOI21x1_ASAP7_75t_R _28110_ (.A1(_05702_),
    .A2(_05703_),
    .B(_05154_),
    .Y(_05704_));
 OAI21x1_ASAP7_75t_R _28111_ (.A1(_05700_),
    .A2(_05704_),
    .B(_05202_),
    .Y(_05705_));
 NAND2x1_ASAP7_75t_SL _28112_ (.A(_05693_),
    .B(_05705_),
    .Y(_05706_));
 OAI21x1_ASAP7_75t_SL _28113_ (.A1(_05669_),
    .A2(_05681_),
    .B(_05706_),
    .Y(_00135_));
 NOR2x1_ASAP7_75t_L _28114_ (.A(_00574_),
    .B(_00483_),
    .Y(_05707_));
 XOR2x2_ASAP7_75t_L _28115_ (.A(_11388_),
    .B(_00648_),
    .Y(_05708_));
 XOR2x2_ASAP7_75t_L _28116_ (.A(_11426_),
    .B(_02992_),
    .Y(_05709_));
 NAND2x1_ASAP7_75t_SL _28117_ (.A(_05708_),
    .B(_05709_),
    .Y(_05710_));
 XNOR2x2_ASAP7_75t_SL _28118_ (.A(_11388_),
    .B(_00648_),
    .Y(_05711_));
 XOR2x2_ASAP7_75t_SL _28119_ (.A(_02992_),
    .B(_11434_),
    .Y(_05712_));
 NAND2x1p5_ASAP7_75t_SL _28120_ (.A(_05712_),
    .B(_05711_),
    .Y(_05713_));
 AOI21x1_ASAP7_75t_SL _28121_ (.A1(_05713_),
    .A2(_05710_),
    .B(_10675_),
    .Y(_05714_));
 OAI21x1_ASAP7_75t_SL _28122_ (.A1(_05707_),
    .A2(_05714_),
    .B(_00881_),
    .Y(_05715_));
 AND2x2_ASAP7_75t_R _28123_ (.A(_10675_),
    .B(_00483_),
    .Y(_05716_));
 NAND2x1_ASAP7_75t_R _28124_ (.A(_05708_),
    .B(_05712_),
    .Y(_05717_));
 NAND2x1p5_ASAP7_75t_L _28125_ (.A(_05711_),
    .B(_05709_),
    .Y(_05718_));
 AOI21x1_ASAP7_75t_SL _28126_ (.A1(_05718_),
    .A2(_05717_),
    .B(_10675_),
    .Y(_05719_));
 INVx1_ASAP7_75t_R _28127_ (.A(_00881_),
    .Y(_05720_));
 OAI21x1_ASAP7_75t_SL _28128_ (.A1(_05716_),
    .A2(_05719_),
    .B(_05720_),
    .Y(_05721_));
 NAND2x2_ASAP7_75t_SL _28129_ (.A(_05715_),
    .B(_05721_),
    .Y(_05722_));
 NAND2x1_ASAP7_75t_L _28131_ (.A(_00484_),
    .B(_10675_),
    .Y(_05723_));
 XOR2x2_ASAP7_75t_SL _28132_ (.A(_11589_),
    .B(_11417_),
    .Y(_05724_));
 NAND2x1p5_ASAP7_75t_SL _28133_ (.A(_05724_),
    .B(_11394_),
    .Y(_05725_));
 NOR2x1_ASAP7_75t_R _28134_ (.A(_11589_),
    .B(_11417_),
    .Y(_05726_));
 NOR2x1_ASAP7_75t_L _28135_ (.A(_00686_),
    .B(_11413_),
    .Y(_05727_));
 OAI21x1_ASAP7_75t_SL _28136_ (.A1(_05727_),
    .A2(_05726_),
    .B(_11388_),
    .Y(_05728_));
 NAND3x1_ASAP7_75t_SL _28137_ (.A(_05725_),
    .B(_05728_),
    .C(_00574_),
    .Y(_05729_));
 INVx1_ASAP7_75t_R _28138_ (.A(_00870_),
    .Y(_05730_));
 AOI21x1_ASAP7_75t_R _28139_ (.A1(_05723_),
    .A2(_05729_),
    .B(_05730_),
    .Y(_05731_));
 OR2x2_ASAP7_75t_R _28140_ (.A(_00574_),
    .B(_00484_),
    .Y(_05732_));
 INVx1_ASAP7_75t_SL _28141_ (.A(_05728_),
    .Y(_05733_));
 INVx2_ASAP7_75t_SL _28142_ (.A(_05725_),
    .Y(_05734_));
 OAI21x1_ASAP7_75t_SL _28143_ (.A1(_05734_),
    .A2(_05733_),
    .B(_00574_),
    .Y(_05735_));
 AOI21x1_ASAP7_75t_SL _28144_ (.A1(_05732_),
    .A2(_05735_),
    .B(_00870_),
    .Y(_05736_));
 NOR2x2_ASAP7_75t_SL _28145_ (.A(_05731_),
    .B(_05736_),
    .Y(_05737_));
 NOR2x1_ASAP7_75t_R _28147_ (.A(_00574_),
    .B(_00485_),
    .Y(_05738_));
 XOR2x1_ASAP7_75t_SL _28148_ (.A(_00649_),
    .Y(_05739_),
    .B(_00680_));
 NOR2x1_ASAP7_75t_R _28149_ (.A(_00584_),
    .B(_05739_),
    .Y(_05740_));
 AND2x2_ASAP7_75t_SL _28150_ (.A(_05739_),
    .B(_00584_),
    .Y(_05741_));
 OAI21x1_ASAP7_75t_SL _28151_ (.A1(_05740_),
    .A2(_05741_),
    .B(_03026_),
    .Y(_05742_));
 XOR2x1_ASAP7_75t_SL _28152_ (.A(_05739_),
    .Y(_05743_),
    .B(_00584_));
 NAND2x1_ASAP7_75t_SL _28153_ (.A(_03025_),
    .B(_05743_),
    .Y(_05744_));
 AOI21x1_ASAP7_75t_SL _28154_ (.A1(_05742_),
    .A2(_05744_),
    .B(_10675_),
    .Y(_05745_));
 INVx1_ASAP7_75t_SL _28155_ (.A(_00892_),
    .Y(_05746_));
 OAI21x1_ASAP7_75t_SL _28156_ (.A1(_05738_),
    .A2(_05745_),
    .B(_05746_),
    .Y(_05747_));
 XOR2x1_ASAP7_75t_SL _28157_ (.A(_00584_),
    .Y(_05748_),
    .B(_00649_));
 NAND2x1_ASAP7_75t_R _28158_ (.A(_11392_),
    .B(_05748_),
    .Y(_05749_));
 INVx1_ASAP7_75t_R _28159_ (.A(_05748_),
    .Y(_05750_));
 NAND2x1_ASAP7_75t_R _28160_ (.A(_00680_),
    .B(_05750_),
    .Y(_05751_));
 AOI21x1_ASAP7_75t_SL _28161_ (.A1(_05749_),
    .A2(_05751_),
    .B(_03026_),
    .Y(_05752_));
 NOR2x1_ASAP7_75t_SL _28162_ (.A(_03025_),
    .B(_05743_),
    .Y(_05753_));
 OAI21x1_ASAP7_75t_SL _28163_ (.A1(_05752_),
    .A2(_05753_),
    .B(_00574_),
    .Y(_05754_));
 INVx1_ASAP7_75t_SL _28164_ (.A(_05738_),
    .Y(_05755_));
 NAND3x2_ASAP7_75t_SL _28165_ (.B(_00892_),
    .C(_05755_),
    .Y(_05756_),
    .A(_05754_));
 NAND2x1_ASAP7_75t_SL _28166_ (.A(_05747_),
    .B(_05756_),
    .Y(_05757_));
 AOI21x1_ASAP7_75t_SL _28169_ (.A1(_05723_),
    .A2(_05729_),
    .B(_00870_),
    .Y(_05759_));
 AOI21x1_ASAP7_75t_SL _28170_ (.A1(_05735_),
    .A2(_05732_),
    .B(_05730_),
    .Y(_05760_));
 NOR2x2_ASAP7_75t_SL _28171_ (.A(_05760_),
    .B(_05759_),
    .Y(_05761_));
 OAI21x1_ASAP7_75t_SL _28173_ (.A1(_05738_),
    .A2(_05745_),
    .B(_00892_),
    .Y(_05762_));
 NAND3x2_ASAP7_75t_SL _28174_ (.B(_05746_),
    .C(_05755_),
    .Y(_05763_),
    .A(_05754_));
 NAND2x2_ASAP7_75t_SL _28175_ (.A(_05762_),
    .B(_05763_),
    .Y(_05764_));
 OAI21x1_ASAP7_75t_SL _28177_ (.A1(_05714_),
    .A2(_05707_),
    .B(_05720_),
    .Y(_05765_));
 OAI21x1_ASAP7_75t_SL _28178_ (.A1(_05716_),
    .A2(_05719_),
    .B(_00881_),
    .Y(_05766_));
 NAND2x2_ASAP7_75t_SL _28179_ (.A(_05766_),
    .B(_05765_),
    .Y(_01342_));
 NAND2x2_ASAP7_75t_SL _28180_ (.A(_01342_),
    .B(_05764_),
    .Y(_05767_));
 INVx1_ASAP7_75t_SL _28181_ (.A(_05767_),
    .Y(_05768_));
 NAND2x1_ASAP7_75t_SL _28182_ (.A(_05722_),
    .B(_05757_),
    .Y(_05769_));
 XNOR2x2_ASAP7_75t_L _28183_ (.A(_03056_),
    .B(_03055_),
    .Y(_05770_));
 XOR2x2_ASAP7_75t_R _28184_ (.A(_11457_),
    .B(_00650_),
    .Y(_05771_));
 AND2x2_ASAP7_75t_SL _28185_ (.A(_05770_),
    .B(_05771_),
    .Y(_05772_));
 OAI21x1_ASAP7_75t_SL _28186_ (.A1(_05771_),
    .A2(_05770_),
    .B(_00574_),
    .Y(_05773_));
 NAND2x1_ASAP7_75t_SL _28187_ (.A(_00511_),
    .B(_10675_),
    .Y(_05774_));
 OAI21x1_ASAP7_75t_SL _28188_ (.A1(_05772_),
    .A2(_05773_),
    .B(_05774_),
    .Y(_05775_));
 XNOR2x2_ASAP7_75t_SL _28189_ (.A(_00895_),
    .B(_05775_),
    .Y(_05776_));
 OAI21x1_ASAP7_75t_SL _28191_ (.A1(_05737_),
    .A2(_05769_),
    .B(_05776_),
    .Y(_05778_));
 NOR2x1_ASAP7_75t_SL _28192_ (.A(_05768_),
    .B(_05778_),
    .Y(_05779_));
 AOI21x1_ASAP7_75t_SL _28195_ (.A1(_05757_),
    .A2(_05761_),
    .B(_05776_),
    .Y(_05782_));
 INVx1_ASAP7_75t_SL _28196_ (.A(_01352_),
    .Y(_05783_));
 AO21x1_ASAP7_75t_SL _28197_ (.A1(_05763_),
    .A2(_05762_),
    .B(_05783_),
    .Y(_05784_));
 XOR2x2_ASAP7_75t_R _28198_ (.A(_11484_),
    .B(_00651_),
    .Y(_05785_));
 XOR2x2_ASAP7_75t_SL _28199_ (.A(_03076_),
    .B(_05785_),
    .Y(_05786_));
 NOR2x1_ASAP7_75t_R _28200_ (.A(_00574_),
    .B(_00510_),
    .Y(_05787_));
 AOI21x1_ASAP7_75t_SL _28201_ (.A1(_00574_),
    .A2(_05786_),
    .B(_05787_),
    .Y(_05788_));
 XNOR2x2_ASAP7_75t_SL _28202_ (.A(_00896_),
    .B(_05788_),
    .Y(_05789_));
 AO21x1_ASAP7_75t_SL _28204_ (.A1(_05782_),
    .A2(_05784_),
    .B(_05789_),
    .Y(_05791_));
 NOR2x1_ASAP7_75t_R _28205_ (.A(_00574_),
    .B(_00509_),
    .Y(_05792_));
 INVx1_ASAP7_75t_R _28206_ (.A(_05792_),
    .Y(_05793_));
 XOR2x2_ASAP7_75t_SL _28207_ (.A(_00587_),
    .B(_00588_),
    .Y(_05794_));
 XOR2x2_ASAP7_75t_R _28208_ (.A(_05794_),
    .B(_14268_),
    .Y(_05795_));
 XOR2x2_ASAP7_75t_SL _28209_ (.A(_05795_),
    .B(_11543_),
    .Y(_05796_));
 NAND2x1_ASAP7_75t_R _28210_ (.A(_00574_),
    .B(_05796_),
    .Y(_05797_));
 INVx1_ASAP7_75t_R _28211_ (.A(_00897_),
    .Y(_05798_));
 AOI21x1_ASAP7_75t_R _28212_ (.A1(_05793_),
    .A2(_05797_),
    .B(_05798_),
    .Y(_05799_));
 AND3x1_ASAP7_75t_SL _28213_ (.A(_05797_),
    .B(_05798_),
    .C(_05793_),
    .Y(_05800_));
 NOR2x1_ASAP7_75t_SL _28214_ (.A(_05799_),
    .B(_05800_),
    .Y(_05801_));
 OAI21x1_ASAP7_75t_SL _28217_ (.A1(_05779_),
    .A2(_05791_),
    .B(_05801_),
    .Y(_05804_));
 NOR2x2_ASAP7_75t_SL _28218_ (.A(_01342_),
    .B(_05757_),
    .Y(_05805_));
 NAND2x2_ASAP7_75t_SL _28219_ (.A(_05737_),
    .B(_05805_),
    .Y(_05806_));
 NAND2x1_ASAP7_75t_SL _28220_ (.A(_05782_),
    .B(_05806_),
    .Y(_05807_));
 NAND2x1_ASAP7_75t_SL _28223_ (.A(_01342_),
    .B(_05757_),
    .Y(_05810_));
 AOI21x1_ASAP7_75t_SL _28224_ (.A1(_05762_),
    .A2(_05763_),
    .B(_01345_),
    .Y(_05811_));
 INVx1_ASAP7_75t_SL _28225_ (.A(_05811_),
    .Y(_05812_));
 XOR2x2_ASAP7_75t_SL _28226_ (.A(_05775_),
    .B(_00895_),
    .Y(_05813_));
 AO21x1_ASAP7_75t_SL _28229_ (.A1(_05810_),
    .A2(_05812_),
    .B(_05813_),
    .Y(_05816_));
 AND3x1_ASAP7_75t_SL _28230_ (.A(_05807_),
    .B(_05789_),
    .C(_05816_),
    .Y(_05817_));
 NOR2x1_ASAP7_75t_SL _28231_ (.A(_05804_),
    .B(_05817_),
    .Y(_05818_));
 NAND2x1_ASAP7_75t_SL _28232_ (.A(_05722_),
    .B(_05761_),
    .Y(_05819_));
 AOI21x1_ASAP7_75t_SL _28236_ (.A1(_05764_),
    .A2(_05761_),
    .B(_05813_),
    .Y(_05823_));
 AOI21x1_ASAP7_75t_SL _28238_ (.A1(_05819_),
    .A2(_05823_),
    .B(_05789_),
    .Y(_05825_));
 AOI21x1_ASAP7_75t_R _28239_ (.A1(_05755_),
    .A2(_05754_),
    .B(_05746_),
    .Y(_05826_));
 NAND2x1_ASAP7_75t_R _28240_ (.A(_00485_),
    .B(_10675_),
    .Y(_05827_));
 NAND3x1_ASAP7_75t_SL _28241_ (.A(_05744_),
    .B(_05742_),
    .C(_00574_),
    .Y(_05828_));
 AOI21x1_ASAP7_75t_R _28242_ (.A1(_05827_),
    .A2(_05828_),
    .B(_00892_),
    .Y(_05829_));
 INVx2_ASAP7_75t_SL _28243_ (.A(_01344_),
    .Y(_05830_));
 OAI21x1_ASAP7_75t_SL _28244_ (.A1(_05826_),
    .A2(_05829_),
    .B(_05830_),
    .Y(_05831_));
 AOI21x1_ASAP7_75t_SL _28245_ (.A1(_05755_),
    .A2(_05754_),
    .B(_00892_),
    .Y(_05832_));
 AOI21x1_ASAP7_75t_SL _28246_ (.A1(_05827_),
    .A2(_05828_),
    .B(_05746_),
    .Y(_05833_));
 OAI21x1_ASAP7_75t_SL _28247_ (.A1(_05832_),
    .A2(_05833_),
    .B(_05783_),
    .Y(_05834_));
 AO21x1_ASAP7_75t_SL _28249_ (.A1(_05831_),
    .A2(_05834_),
    .B(_05776_),
    .Y(_05836_));
 AND2x2_ASAP7_75t_SL _28250_ (.A(_05825_),
    .B(_05836_),
    .Y(_05837_));
 AOI21x1_ASAP7_75t_SL _28253_ (.A1(_01347_),
    .A2(_05764_),
    .B(_05776_),
    .Y(_05840_));
 NOR2x1_ASAP7_75t_SL _28254_ (.A(_01342_),
    .B(_05764_),
    .Y(_05841_));
 NAND2x1_ASAP7_75t_SL _28255_ (.A(_05761_),
    .B(_05841_),
    .Y(_05842_));
 NAND2x1_ASAP7_75t_SL _28256_ (.A(_05840_),
    .B(_05842_),
    .Y(_05843_));
 INVx2_ASAP7_75t_SL _28257_ (.A(_05789_),
    .Y(_05844_));
 AOI21x1_ASAP7_75t_SL _28259_ (.A1(_05757_),
    .A2(_05761_),
    .B(_05813_),
    .Y(_05846_));
 NOR2x1_ASAP7_75t_SL _28260_ (.A(_05844_),
    .B(_05846_),
    .Y(_05847_));
 AO21x1_ASAP7_75t_SL _28262_ (.A1(_05843_),
    .A2(_05847_),
    .B(_05801_),
    .Y(_05849_));
 XOR2x2_ASAP7_75t_R _28263_ (.A(_00588_),
    .B(_00589_),
    .Y(_05850_));
 XOR2x2_ASAP7_75t_R _28264_ (.A(_05850_),
    .B(_14295_),
    .Y(_05851_));
 XOR2x2_ASAP7_75t_R _28265_ (.A(_05851_),
    .B(_11504_),
    .Y(_05852_));
 NOR2x1_ASAP7_75t_SL _28266_ (.A(_00574_),
    .B(_00507_),
    .Y(_05853_));
 AO21x1_ASAP7_75t_SL _28267_ (.A1(_05852_),
    .A2(_00574_),
    .B(_05853_),
    .Y(_05854_));
 XOR2x2_ASAP7_75t_SL _28268_ (.A(_05854_),
    .B(_00898_),
    .Y(_05855_));
 INVx1_ASAP7_75t_SL _28269_ (.A(_05855_),
    .Y(_05856_));
 OAI21x1_ASAP7_75t_SL _28271_ (.A1(_05837_),
    .A2(_05849_),
    .B(_05856_),
    .Y(_05858_));
 XOR2x2_ASAP7_75t_R _28272_ (.A(_00589_),
    .B(_00590_),
    .Y(_05859_));
 XOR2x2_ASAP7_75t_R _28273_ (.A(_05859_),
    .B(_00685_),
    .Y(_05860_));
 XOR2x2_ASAP7_75t_SL _28274_ (.A(_05860_),
    .B(_11591_),
    .Y(_05861_));
 NOR2x1_ASAP7_75t_SL _28275_ (.A(_00574_),
    .B(_00506_),
    .Y(_05862_));
 AO21x1_ASAP7_75t_SL _28276_ (.A1(_05861_),
    .A2(_00574_),
    .B(_05862_),
    .Y(_05863_));
 XOR2x2_ASAP7_75t_SL _28277_ (.A(_05863_),
    .B(_00899_),
    .Y(_05864_));
 OAI21x1_ASAP7_75t_SL _28279_ (.A1(_05818_),
    .A2(_05858_),
    .B(_05864_),
    .Y(_05866_));
 NAND2x1_ASAP7_75t_SL _28280_ (.A(_05757_),
    .B(_05737_),
    .Y(_05867_));
 INVx1_ASAP7_75t_SL _28281_ (.A(_05867_),
    .Y(_05868_));
 OAI21x1_ASAP7_75t_SL _28283_ (.A1(_01342_),
    .A2(_05737_),
    .B(_05813_),
    .Y(_05870_));
 OAI21x1_ASAP7_75t_SL _28285_ (.A1(_05868_),
    .A2(_05870_),
    .B(_05844_),
    .Y(_05872_));
 NOR2x1_ASAP7_75t_SL _28286_ (.A(_05722_),
    .B(_05737_),
    .Y(_05873_));
 OAI21x1_ASAP7_75t_R _28287_ (.A1(_05757_),
    .A2(_05761_),
    .B(_05776_),
    .Y(_05874_));
 NOR2x1_ASAP7_75t_SL _28288_ (.A(_05873_),
    .B(_05874_),
    .Y(_05875_));
 INVx1_ASAP7_75t_SL _28289_ (.A(_05801_),
    .Y(_05876_));
 OA21x2_ASAP7_75t_SL _28292_ (.A1(_05872_),
    .A2(_05875_),
    .B(_05876_),
    .Y(_05879_));
 INVx1_ASAP7_75t_SL _28293_ (.A(_01349_),
    .Y(_05880_));
 AO21x1_ASAP7_75t_SL _28294_ (.A1(_05763_),
    .A2(_05762_),
    .B(_05880_),
    .Y(_05881_));
 INVx1_ASAP7_75t_SL _28295_ (.A(_01343_),
    .Y(_05882_));
 AOI21x1_ASAP7_75t_SL _28296_ (.A1(_05747_),
    .A2(_05756_),
    .B(_05882_),
    .Y(_05883_));
 INVx2_ASAP7_75t_SL _28297_ (.A(_05883_),
    .Y(_05884_));
 AO21x1_ASAP7_75t_SL _28299_ (.A1(_05881_),
    .A2(_05884_),
    .B(_05776_),
    .Y(_05886_));
 NAND2x1_ASAP7_75t_SL _28300_ (.A(_05722_),
    .B(_05737_),
    .Y(_05887_));
 AOI21x1_ASAP7_75t_SL _28301_ (.A1(_05762_),
    .A2(_05763_),
    .B(_05830_),
    .Y(_05888_));
 NOR2x1p5_ASAP7_75t_SL _28302_ (.A(_05888_),
    .B(_05813_),
    .Y(_05889_));
 OAI21x1_ASAP7_75t_SL _28303_ (.A1(_05764_),
    .A2(_05887_),
    .B(_05889_),
    .Y(_05890_));
 NAND3x1_ASAP7_75t_SL _28304_ (.A(_05886_),
    .B(_05890_),
    .C(_05789_),
    .Y(_05891_));
 AOI21x1_ASAP7_75t_SL _28305_ (.A1(_05762_),
    .A2(_05763_),
    .B(_01344_),
    .Y(_05892_));
 OA21x2_ASAP7_75t_SL _28307_ (.A1(_05883_),
    .A2(_05892_),
    .B(_05813_),
    .Y(_05894_));
 NOR2x1_ASAP7_75t_SL _28308_ (.A(_01343_),
    .B(_05757_),
    .Y(_05895_));
 INVx2_ASAP7_75t_SL _28309_ (.A(_05895_),
    .Y(_05896_));
 AOI21x1_ASAP7_75t_SL _28310_ (.A1(_05880_),
    .A2(_05757_),
    .B(_05813_),
    .Y(_05897_));
 AND2x2_ASAP7_75t_SL _28311_ (.A(_05896_),
    .B(_05897_),
    .Y(_05898_));
 OAI21x1_ASAP7_75t_SL _28312_ (.A1(_05894_),
    .A2(_05898_),
    .B(_05789_),
    .Y(_05899_));
 AOI21x1_ASAP7_75t_SL _28313_ (.A1(_05747_),
    .A2(_05756_),
    .B(_05830_),
    .Y(_05900_));
 NAND2x1_ASAP7_75t_SL _28314_ (.A(_05813_),
    .B(_05900_),
    .Y(_05901_));
 OAI21x1_ASAP7_75t_R _28315_ (.A1(_05722_),
    .A2(_05764_),
    .B(_05776_),
    .Y(_05902_));
 AO21x1_ASAP7_75t_SL _28316_ (.A1(_05776_),
    .A2(_05888_),
    .B(_05789_),
    .Y(_05903_));
 AO21x1_ASAP7_75t_SL _28317_ (.A1(_05901_),
    .A2(_05902_),
    .B(_05903_),
    .Y(_05904_));
 AOI21x1_ASAP7_75t_SL _28318_ (.A1(_05899_),
    .A2(_05904_),
    .B(_05876_),
    .Y(_05905_));
 AOI211x1_ASAP7_75t_SL _28319_ (.A1(_05879_),
    .A2(_05891_),
    .B(_05856_),
    .C(_05905_),
    .Y(_05906_));
 AOI21x1_ASAP7_75t_SL _28320_ (.A1(_05747_),
    .A2(_05756_),
    .B(_01347_),
    .Y(_05907_));
 AOI21x1_ASAP7_75t_SL _28321_ (.A1(_05722_),
    .A2(_05761_),
    .B(_05757_),
    .Y(_05908_));
 OAI21x1_ASAP7_75t_SL _28322_ (.A1(_05907_),
    .A2(_05908_),
    .B(_05776_),
    .Y(_05909_));
 INVx1_ASAP7_75t_SL _28323_ (.A(_05782_),
    .Y(_05910_));
 NOR2x1_ASAP7_75t_R _28326_ (.A(_01345_),
    .B(_05764_),
    .Y(_05913_));
 AOI21x1_ASAP7_75t_SL _28327_ (.A1(_05776_),
    .A2(_05913_),
    .B(_05844_),
    .Y(_05914_));
 OA21x2_ASAP7_75t_SL _28328_ (.A1(_05895_),
    .A2(_05910_),
    .B(_05914_),
    .Y(_05915_));
 AOI21x1_ASAP7_75t_SL _28329_ (.A1(_05747_),
    .A2(_05756_),
    .B(_01344_),
    .Y(_05916_));
 NOR2x1p5_ASAP7_75t_SL _28330_ (.A(_05813_),
    .B(_05916_),
    .Y(_05917_));
 AOI21x1_ASAP7_75t_SL _28331_ (.A1(_01357_),
    .A2(_05813_),
    .B(_05917_),
    .Y(_05918_));
 OAI21x1_ASAP7_75t_SL _28332_ (.A1(_05789_),
    .A2(_05918_),
    .B(_05801_),
    .Y(_05919_));
 AOI21x1_ASAP7_75t_SL _28333_ (.A1(_05909_),
    .A2(_05915_),
    .B(_05919_),
    .Y(_05920_));
 AO21x1_ASAP7_75t_SL _28334_ (.A1(_05811_),
    .A2(_05813_),
    .B(_05789_),
    .Y(_05921_));
 INVx1_ASAP7_75t_SL _28335_ (.A(_05897_),
    .Y(_05922_));
 NAND2x1_ASAP7_75t_SL _28336_ (.A(_05722_),
    .B(_05764_),
    .Y(_05923_));
 NOR2x1_ASAP7_75t_SL _28337_ (.A(_05737_),
    .B(_05923_),
    .Y(_05924_));
 NOR2x1_ASAP7_75t_SL _28338_ (.A(_05922_),
    .B(_05924_),
    .Y(_05925_));
 OAI21x1_ASAP7_75t_SL _28339_ (.A1(_05921_),
    .A2(_05925_),
    .B(_05876_),
    .Y(_05926_));
 INVx1_ASAP7_75t_SL _28340_ (.A(_05924_),
    .Y(_05927_));
 AOI21x1_ASAP7_75t_SL _28341_ (.A1(_01350_),
    .A2(_05757_),
    .B(_05776_),
    .Y(_05928_));
 AND2x2_ASAP7_75t_SL _28343_ (.A(_05811_),
    .B(_05776_),
    .Y(_05930_));
 AOI211x1_ASAP7_75t_SL _28344_ (.A1(_05927_),
    .A2(_05928_),
    .B(_05844_),
    .C(_05930_),
    .Y(_05931_));
 OAI21x1_ASAP7_75t_SL _28346_ (.A1(_05926_),
    .A2(_05931_),
    .B(_05855_),
    .Y(_05933_));
 AO21x2_ASAP7_75t_SL _28347_ (.A1(_05756_),
    .A2(_05747_),
    .B(_05880_),
    .Y(_05934_));
 NAND2x1_ASAP7_75t_L _28348_ (.A(_05764_),
    .B(_05737_),
    .Y(_05935_));
 AOI21x1_ASAP7_75t_SL _28349_ (.A1(_05934_),
    .A2(_05935_),
    .B(_05776_),
    .Y(_05936_));
 AOI21x1_ASAP7_75t_SL _28350_ (.A1(_05722_),
    .A2(_05764_),
    .B(_05813_),
    .Y(_05937_));
 INVx2_ASAP7_75t_SL _28351_ (.A(_05916_),
    .Y(_05938_));
 AO21x1_ASAP7_75t_SL _28352_ (.A1(_05937_),
    .A2(_05938_),
    .B(_05844_),
    .Y(_05939_));
 OAI21x1_ASAP7_75t_SL _28353_ (.A1(_05883_),
    .A2(_05811_),
    .B(_05776_),
    .Y(_05940_));
 NOR2x1_ASAP7_75t_SL _28354_ (.A(_05789_),
    .B(_05840_),
    .Y(_05941_));
 AOI21x1_ASAP7_75t_SL _28355_ (.A1(_05940_),
    .A2(_05941_),
    .B(_05801_),
    .Y(_05942_));
 OAI21x1_ASAP7_75t_SL _28356_ (.A1(_05936_),
    .A2(_05939_),
    .B(_05942_),
    .Y(_05943_));
 INVx1_ASAP7_75t_SL _28357_ (.A(_05806_),
    .Y(_05944_));
 INVx2_ASAP7_75t_SL _28358_ (.A(_01347_),
    .Y(_05945_));
 OAI21x1_ASAP7_75t_SL _28359_ (.A1(_05832_),
    .A2(_05833_),
    .B(_05945_),
    .Y(_05946_));
 OA21x2_ASAP7_75t_SL _28360_ (.A1(_05946_),
    .A2(_05813_),
    .B(_05789_),
    .Y(_05947_));
 OAI21x1_ASAP7_75t_SL _28361_ (.A1(_05910_),
    .A2(_05944_),
    .B(_05947_),
    .Y(_05948_));
 AOI21x1_ASAP7_75t_SL _28362_ (.A1(_05762_),
    .A2(_05763_),
    .B(_01350_),
    .Y(_05949_));
 OAI21x1_ASAP7_75t_R _28363_ (.A1(_05907_),
    .A2(_05949_),
    .B(_05776_),
    .Y(_05950_));
 NOR2x2_ASAP7_75t_SL _28364_ (.A(_05888_),
    .B(_05776_),
    .Y(_05951_));
 NOR2x1p5_ASAP7_75t_SL _28365_ (.A(_05951_),
    .B(_05789_),
    .Y(_05952_));
 AOI21x1_ASAP7_75t_SL _28367_ (.A1(_05950_),
    .A2(_05952_),
    .B(_05876_),
    .Y(_05954_));
 AOI21x1_ASAP7_75t_SL _28368_ (.A1(_05954_),
    .A2(_05948_),
    .B(_05855_),
    .Y(_05955_));
 AOI21x1_ASAP7_75t_SL _28369_ (.A1(_05955_),
    .A2(_05943_),
    .B(_05864_),
    .Y(_05956_));
 OAI21x1_ASAP7_75t_SL _28370_ (.A1(_05920_),
    .A2(_05933_),
    .B(_05956_),
    .Y(_05957_));
 OAI21x1_ASAP7_75t_SL _28371_ (.A1(_05866_),
    .A2(_05906_),
    .B(_05957_),
    .Y(_00136_));
 AOI21x1_ASAP7_75t_SL _28372_ (.A1(_05722_),
    .A2(_05737_),
    .B(_05757_),
    .Y(_05958_));
 INVx1_ASAP7_75t_SL _28373_ (.A(_05958_),
    .Y(_05959_));
 AOI21x1_ASAP7_75t_SL _28374_ (.A1(_01352_),
    .A2(_05757_),
    .B(_05776_),
    .Y(_05960_));
 AOI21x1_ASAP7_75t_SL _28375_ (.A1(_05767_),
    .A2(_05960_),
    .B(_05789_),
    .Y(_05961_));
 OA21x2_ASAP7_75t_SL _28376_ (.A1(_05813_),
    .A2(_05959_),
    .B(_05961_),
    .Y(_05962_));
 AOI21x1_ASAP7_75t_SL _28377_ (.A1(_05722_),
    .A2(_05737_),
    .B(_05764_),
    .Y(_05963_));
 OAI21x1_ASAP7_75t_SL _28379_ (.A1(_05888_),
    .A2(_05963_),
    .B(_05813_),
    .Y(_05965_));
 OAI21x1_ASAP7_75t_SL _28380_ (.A1(_05826_),
    .A2(_05829_),
    .B(_05945_),
    .Y(_05966_));
 OA21x2_ASAP7_75t_SL _28381_ (.A1(_05966_),
    .A2(_05813_),
    .B(_05789_),
    .Y(_05967_));
 AO21x1_ASAP7_75t_SL _28382_ (.A1(_05965_),
    .A2(_05967_),
    .B(_05801_),
    .Y(_05968_));
 OAI21x1_ASAP7_75t_SL _28383_ (.A1(_05962_),
    .A2(_05968_),
    .B(_05856_),
    .Y(_05969_));
 AO21x1_ASAP7_75t_SL _28384_ (.A1(_05763_),
    .A2(_05762_),
    .B(_05882_),
    .Y(_05970_));
 AO32x1_ASAP7_75t_SL _28385_ (.A1(_05776_),
    .A2(_05867_),
    .A3(_05970_),
    .B1(_05951_),
    .B2(_05946_),
    .Y(_05971_));
 NAND2x1_ASAP7_75t_SL _28386_ (.A(_05764_),
    .B(_05761_),
    .Y(_05972_));
 AO21x1_ASAP7_75t_SL _28387_ (.A1(_05972_),
    .A2(_05887_),
    .B(_05776_),
    .Y(_05973_));
 AOI21x1_ASAP7_75t_SL _28388_ (.A1(_05972_),
    .A2(_05917_),
    .B(_05844_),
    .Y(_05974_));
 AO21x1_ASAP7_75t_SL _28389_ (.A1(_05973_),
    .A2(_05974_),
    .B(_05876_),
    .Y(_05975_));
 AOI21x1_ASAP7_75t_SL _28390_ (.A1(_05844_),
    .A2(_05971_),
    .B(_05975_),
    .Y(_05976_));
 NOR2x1_ASAP7_75t_SL _28391_ (.A(_05776_),
    .B(_05764_),
    .Y(_05977_));
 NAND2x1_ASAP7_75t_SL _28392_ (.A(_05977_),
    .B(_05819_),
    .Y(_05978_));
 NAND2x1_ASAP7_75t_SL _28393_ (.A(_01342_),
    .B(_05761_),
    .Y(_05979_));
 NAND2x1_ASAP7_75t_SL _28394_ (.A(_05979_),
    .B(_05937_),
    .Y(_05980_));
 AOI21x1_ASAP7_75t_SL _28397_ (.A1(_05978_),
    .A2(_05980_),
    .B(_05844_),
    .Y(_05983_));
 INVx2_ASAP7_75t_SL _28398_ (.A(_05888_),
    .Y(_05984_));
 NAND2x1_ASAP7_75t_SL _28399_ (.A(_05984_),
    .B(_05782_),
    .Y(_05985_));
 AO21x1_ASAP7_75t_R _28400_ (.A1(_05763_),
    .A2(_05762_),
    .B(_05945_),
    .Y(_05986_));
 AOI21x1_ASAP7_75t_SL _28401_ (.A1(_05757_),
    .A2(_05737_),
    .B(_05813_),
    .Y(_05987_));
 NAND2x1_ASAP7_75t_SL _28402_ (.A(_05986_),
    .B(_05987_),
    .Y(_05988_));
 AOI21x1_ASAP7_75t_SL _28404_ (.A1(_05985_),
    .A2(_05988_),
    .B(_05789_),
    .Y(_05990_));
 OAI21x1_ASAP7_75t_SL _28405_ (.A1(_05983_),
    .A2(_05990_),
    .B(_05876_),
    .Y(_05991_));
 NOR2x1p5_ASAP7_75t_SL _28406_ (.A(_05900_),
    .B(_05776_),
    .Y(_05992_));
 AOI21x1_ASAP7_75t_SL _28407_ (.A1(_05784_),
    .A2(_05992_),
    .B(_05844_),
    .Y(_05993_));
 NAND2x1_ASAP7_75t_SL _28408_ (.A(_05993_),
    .B(_05909_),
    .Y(_05994_));
 OA21x2_ASAP7_75t_SL _28409_ (.A1(_05946_),
    .A2(_05813_),
    .B(_05844_),
    .Y(_05995_));
 AOI21x1_ASAP7_75t_SL _28410_ (.A1(_05722_),
    .A2(_05757_),
    .B(_05776_),
    .Y(_05996_));
 NOR2x1_ASAP7_75t_SL _28411_ (.A(_05768_),
    .B(_05996_),
    .Y(_05997_));
 AOI21x1_ASAP7_75t_SL _28412_ (.A1(_05995_),
    .A2(_05997_),
    .B(_05876_),
    .Y(_05998_));
 AOI21x1_ASAP7_75t_SL _28413_ (.A1(_05994_),
    .A2(_05998_),
    .B(_05856_),
    .Y(_05999_));
 AOI21x1_ASAP7_75t_SL _28414_ (.A1(_05991_),
    .A2(_05999_),
    .B(_05864_),
    .Y(_06000_));
 OAI21x1_ASAP7_75t_SL _28415_ (.A1(_05976_),
    .A2(_05969_),
    .B(_06000_),
    .Y(_06001_));
 NAND2x1_ASAP7_75t_R _28416_ (.A(_05810_),
    .B(_05840_),
    .Y(_06002_));
 AOI21x1_ASAP7_75t_SL _28417_ (.A1(_05764_),
    .A2(_05737_),
    .B(_05813_),
    .Y(_06003_));
 NAND2x1_ASAP7_75t_R _28418_ (.A(_05769_),
    .B(_06003_),
    .Y(_06004_));
 NAND2x1_ASAP7_75t_SL _28419_ (.A(_06002_),
    .B(_06004_),
    .Y(_06005_));
 AO21x1_ASAP7_75t_R _28420_ (.A1(_05756_),
    .A2(_05747_),
    .B(_01343_),
    .Y(_06006_));
 AOI21x1_ASAP7_75t_R _28421_ (.A1(_06006_),
    .A2(_05823_),
    .B(_05801_),
    .Y(_06007_));
 AOI21x1_ASAP7_75t_SL _28422_ (.A1(_05722_),
    .A2(_05761_),
    .B(_05764_),
    .Y(_06008_));
 OAI21x1_ASAP7_75t_R _28423_ (.A1(_05958_),
    .A2(_06008_),
    .B(_05813_),
    .Y(_06009_));
 NAND2x1_ASAP7_75t_SL _28424_ (.A(_06007_),
    .B(_06009_),
    .Y(_06010_));
 OAI21x1_ASAP7_75t_SL _28425_ (.A1(_05876_),
    .A2(_06005_),
    .B(_06010_),
    .Y(_06011_));
 NAND2x1_ASAP7_75t_R _28427_ (.A(_01359_),
    .B(_05813_),
    .Y(_06013_));
 OA21x2_ASAP7_75t_SL _28428_ (.A1(_05876_),
    .A2(_06013_),
    .B(_05789_),
    .Y(_06014_));
 NAND2x1_ASAP7_75t_SL _28429_ (.A(_05897_),
    .B(_05806_),
    .Y(_06015_));
 AO21x1_ASAP7_75t_SL _28430_ (.A1(_06014_),
    .A2(_06015_),
    .B(_05856_),
    .Y(_06016_));
 AOI21x1_ASAP7_75t_SL _28431_ (.A1(_05844_),
    .A2(_06011_),
    .B(_06016_),
    .Y(_06017_));
 NAND2x1_ASAP7_75t_R _28432_ (.A(_01345_),
    .B(_05757_),
    .Y(_06018_));
 AOI21x1_ASAP7_75t_R _28433_ (.A1(_01352_),
    .A2(_05764_),
    .B(_05813_),
    .Y(_06019_));
 AOI21x1_ASAP7_75t_SL _28434_ (.A1(_06018_),
    .A2(_06019_),
    .B(_05789_),
    .Y(_06020_));
 NAND2x1_ASAP7_75t_SL _28435_ (.A(_06020_),
    .B(_05965_),
    .Y(_06021_));
 NOR2x1p5_ASAP7_75t_SL _28436_ (.A(_05951_),
    .B(_05844_),
    .Y(_06022_));
 NAND2x1_ASAP7_75t_SL _28437_ (.A(_05846_),
    .B(_05806_),
    .Y(_06023_));
 AOI21x1_ASAP7_75t_SL _28438_ (.A1(_06022_),
    .A2(_06023_),
    .B(_05876_),
    .Y(_06024_));
 NAND2x1_ASAP7_75t_SL _28439_ (.A(_06021_),
    .B(_06024_),
    .Y(_06025_));
 AOI21x1_ASAP7_75t_SL _28440_ (.A1(_05776_),
    .A2(_05868_),
    .B(_05789_),
    .Y(_06026_));
 INVx1_ASAP7_75t_SL _28441_ (.A(_06026_),
    .Y(_06027_));
 AO21x1_ASAP7_75t_SL _28442_ (.A1(_05896_),
    .A2(_05992_),
    .B(_05930_),
    .Y(_06028_));
 NAND2x1_ASAP7_75t_SL _28443_ (.A(_06006_),
    .B(_06003_),
    .Y(_06029_));
 AOI21x1_ASAP7_75t_SL _28444_ (.A1(_05810_),
    .A2(_05840_),
    .B(_05844_),
    .Y(_06030_));
 AOI21x1_ASAP7_75t_SL _28445_ (.A1(_06029_),
    .A2(_06030_),
    .B(_05801_),
    .Y(_06031_));
 OAI21x1_ASAP7_75t_SL _28446_ (.A1(_06027_),
    .A2(_06028_),
    .B(_06031_),
    .Y(_06032_));
 AOI21x1_ASAP7_75t_SL _28447_ (.A1(_06025_),
    .A2(_06032_),
    .B(_05855_),
    .Y(_06033_));
 OAI21x1_ASAP7_75t_SL _28448_ (.A1(_06017_),
    .A2(_06033_),
    .B(_05864_),
    .Y(_06034_));
 NAND2x1_ASAP7_75t_SL _28449_ (.A(_06034_),
    .B(_06001_),
    .Y(_00137_));
 AOI21x1_ASAP7_75t_SL _28450_ (.A1(_01342_),
    .A2(_05757_),
    .B(_05776_),
    .Y(_06035_));
 NAND2x1_ASAP7_75t_SL _28451_ (.A(_05972_),
    .B(_06035_),
    .Y(_06036_));
 AOI21x1_ASAP7_75t_SL _28452_ (.A1(_05938_),
    .A2(_05937_),
    .B(_05789_),
    .Y(_06037_));
 NAND2x1_ASAP7_75t_SL _28453_ (.A(_06036_),
    .B(_06037_),
    .Y(_06038_));
 OA21x2_ASAP7_75t_SL _28454_ (.A1(_01357_),
    .A2(_05813_),
    .B(_05789_),
    .Y(_06039_));
 OAI21x1_ASAP7_75t_SL _28455_ (.A1(_05757_),
    .A2(_05819_),
    .B(_05992_),
    .Y(_06040_));
 AOI21x1_ASAP7_75t_SL _28456_ (.A1(_06039_),
    .A2(_06040_),
    .B(_05801_),
    .Y(_06041_));
 NAND2x1_ASAP7_75t_SL _28457_ (.A(_06038_),
    .B(_06041_),
    .Y(_06042_));
 NAND2x1_ASAP7_75t_SL _28458_ (.A(_01359_),
    .B(_05776_),
    .Y(_06043_));
 AOI21x1_ASAP7_75t_SL _28459_ (.A1(_05722_),
    .A2(_05764_),
    .B(_05776_),
    .Y(_06044_));
 AOI21x1_ASAP7_75t_SL _28460_ (.A1(_05979_),
    .A2(_06044_),
    .B(_05844_),
    .Y(_06045_));
 AOI21x1_ASAP7_75t_SL _28461_ (.A1(_06043_),
    .A2(_06045_),
    .B(_05876_),
    .Y(_06046_));
 AND2x2_ASAP7_75t_SL _28462_ (.A(_05937_),
    .B(_05884_),
    .Y(_06047_));
 NAND2x1_ASAP7_75t_SL _28463_ (.A(_05813_),
    .B(_05881_),
    .Y(_06048_));
 NOR2x1_ASAP7_75t_SL _28464_ (.A(_05916_),
    .B(_06048_),
    .Y(_06049_));
 OAI21x1_ASAP7_75t_SL _28465_ (.A1(_06047_),
    .A2(_06049_),
    .B(_05844_),
    .Y(_06050_));
 NAND2x1_ASAP7_75t_SL _28466_ (.A(_06046_),
    .B(_06050_),
    .Y(_06051_));
 AOI21x1_ASAP7_75t_SL _28467_ (.A1(_06042_),
    .A2(_06051_),
    .B(_05855_),
    .Y(_06052_));
 NAND2x1_ASAP7_75t_SL _28468_ (.A(_01356_),
    .B(_05813_),
    .Y(_06053_));
 AOI21x1_ASAP7_75t_SL _28469_ (.A1(_06053_),
    .A2(_05778_),
    .B(_05844_),
    .Y(_06054_));
 OAI21x1_ASAP7_75t_SL _28470_ (.A1(_05764_),
    .A2(_05761_),
    .B(_05722_),
    .Y(_06055_));
 NOR2x1_ASAP7_75t_SL _28471_ (.A(_01361_),
    .B(_05813_),
    .Y(_06056_));
 AOI21x1_ASAP7_75t_SL _28472_ (.A1(_05813_),
    .A2(_06055_),
    .B(_06056_),
    .Y(_06057_));
 NOR2x1_ASAP7_75t_SL _28473_ (.A(_05789_),
    .B(_06057_),
    .Y(_06058_));
 OAI21x1_ASAP7_75t_SL _28474_ (.A1(_06054_),
    .A2(_06058_),
    .B(_05801_),
    .Y(_06059_));
 AND2x2_ASAP7_75t_R _28475_ (.A(_01345_),
    .B(_01347_),
    .Y(_06060_));
 NOR2x1_ASAP7_75t_SL _28476_ (.A(_06060_),
    .B(_05757_),
    .Y(_06061_));
 OAI21x1_ASAP7_75t_SL _28477_ (.A1(_06061_),
    .A2(_05963_),
    .B(_05813_),
    .Y(_06062_));
 AOI21x1_ASAP7_75t_SL _28478_ (.A1(_05897_),
    .A2(_05806_),
    .B(_05789_),
    .Y(_06063_));
 NAND2x1_ASAP7_75t_SL _28479_ (.A(_06062_),
    .B(_06063_),
    .Y(_06064_));
 AOI21x1_ASAP7_75t_SL _28480_ (.A1(_05831_),
    .A2(_05946_),
    .B(_05776_),
    .Y(_06065_));
 NOR2x1_ASAP7_75t_SL _28481_ (.A(_05813_),
    .B(_05970_),
    .Y(_06066_));
 NOR2x1_ASAP7_75t_SL _28482_ (.A(_06065_),
    .B(_06066_),
    .Y(_06067_));
 AOI21x1_ASAP7_75t_SL _28483_ (.A1(_05789_),
    .A2(_06067_),
    .B(_05801_),
    .Y(_06068_));
 NAND2x1_ASAP7_75t_SL _28484_ (.A(_06064_),
    .B(_06068_),
    .Y(_06069_));
 AOI21x1_ASAP7_75t_SL _28485_ (.A1(_06059_),
    .A2(_06069_),
    .B(_05856_),
    .Y(_06070_));
 INVx2_ASAP7_75t_SL _28486_ (.A(_05864_),
    .Y(_06071_));
 OAI21x1_ASAP7_75t_SL _28487_ (.A1(_06052_),
    .A2(_06070_),
    .B(_06071_),
    .Y(_06072_));
 AO21x1_ASAP7_75t_SL _28488_ (.A1(_05923_),
    .A2(_05946_),
    .B(_05776_),
    .Y(_06073_));
 AND2x2_ASAP7_75t_SL _28489_ (.A(_05950_),
    .B(_05789_),
    .Y(_06074_));
 NAND2x1_ASAP7_75t_SL _28490_ (.A(_06073_),
    .B(_06074_),
    .Y(_06075_));
 INVx1_ASAP7_75t_SL _28491_ (.A(_05949_),
    .Y(_06076_));
 OA21x2_ASAP7_75t_SL _28492_ (.A1(_06076_),
    .A2(_05813_),
    .B(_05844_),
    .Y(_06077_));
 OAI21x1_ASAP7_75t_SL _28493_ (.A1(_05757_),
    .A2(_05761_),
    .B(_05813_),
    .Y(_06078_));
 NAND2x1_ASAP7_75t_SL _28494_ (.A(_05776_),
    .B(_05834_),
    .Y(_06079_));
 OAI21x1_ASAP7_75t_SL _28495_ (.A1(_05907_),
    .A2(_06078_),
    .B(_06079_),
    .Y(_06080_));
 AOI21x1_ASAP7_75t_SL _28496_ (.A1(_06077_),
    .A2(_06080_),
    .B(_05876_),
    .Y(_06081_));
 NAND2x1_ASAP7_75t_SL _28497_ (.A(_06075_),
    .B(_06081_),
    .Y(_06082_));
 AOI21x1_ASAP7_75t_SL _28498_ (.A1(_01350_),
    .A2(_05757_),
    .B(_05813_),
    .Y(_06083_));
 NAND2x1_ASAP7_75t_SL _28499_ (.A(_05972_),
    .B(_06083_),
    .Y(_06084_));
 NAND2x1p5_ASAP7_75t_SL _28500_ (.A(_05951_),
    .B(_05938_),
    .Y(_06085_));
 AOI21x1_ASAP7_75t_SL _28501_ (.A1(_06084_),
    .A2(_06085_),
    .B(_05844_),
    .Y(_06086_));
 AND2x2_ASAP7_75t_SL _28502_ (.A(_06035_),
    .B(_06076_),
    .Y(_06087_));
 INVx1_ASAP7_75t_SL _28503_ (.A(_05834_),
    .Y(_06088_));
 OAI21x1_ASAP7_75t_SL _28504_ (.A1(_06088_),
    .A2(_05874_),
    .B(_05844_),
    .Y(_06089_));
 NOR2x1_ASAP7_75t_SL _28505_ (.A(_06087_),
    .B(_06089_),
    .Y(_06090_));
 OAI21x1_ASAP7_75t_SL _28506_ (.A1(_06090_),
    .A2(_06086_),
    .B(_05876_),
    .Y(_06091_));
 AOI21x1_ASAP7_75t_SL _28507_ (.A1(_06091_),
    .A2(_06082_),
    .B(_05855_),
    .Y(_06092_));
 NOR2x1_ASAP7_75t_SL _28508_ (.A(_05913_),
    .B(_06078_),
    .Y(_06093_));
 OAI21x1_ASAP7_75t_SL _28509_ (.A1(_05892_),
    .A2(_05902_),
    .B(_05844_),
    .Y(_06094_));
 OAI21x1_ASAP7_75t_SL _28510_ (.A1(_06093_),
    .A2(_06094_),
    .B(_05876_),
    .Y(_06095_));
 AO21x1_ASAP7_75t_SL _28511_ (.A1(_05763_),
    .A2(_05762_),
    .B(_01352_),
    .Y(_06096_));
 INVx1_ASAP7_75t_R _28512_ (.A(_06096_),
    .Y(_06097_));
 OAI21x1_ASAP7_75t_SL _28513_ (.A1(_06097_),
    .A2(_05963_),
    .B(_05813_),
    .Y(_06098_));
 AOI21x1_ASAP7_75t_SL _28514_ (.A1(_05778_),
    .A2(_06098_),
    .B(_05844_),
    .Y(_06099_));
 OAI21x1_ASAP7_75t_SL _28515_ (.A1(_06095_),
    .A2(_06099_),
    .B(_05855_),
    .Y(_06100_));
 NOR2x1_ASAP7_75t_SL _28516_ (.A(_05907_),
    .B(_05908_),
    .Y(_06101_));
 AOI21x1_ASAP7_75t_SL _28517_ (.A1(_05813_),
    .A2(_06101_),
    .B(_05939_),
    .Y(_06102_));
 AOI21x1_ASAP7_75t_SL _28518_ (.A1(_01347_),
    .A2(_05764_),
    .B(_05813_),
    .Y(_06103_));
 AO21x1_ASAP7_75t_R _28519_ (.A1(_05756_),
    .A2(_05747_),
    .B(_05783_),
    .Y(_06104_));
 AOI22x1_ASAP7_75t_SL _28520_ (.A1(_06103_),
    .A2(_06104_),
    .B1(_06055_),
    .B2(_05813_),
    .Y(_06105_));
 OAI21x1_ASAP7_75t_SL _28521_ (.A1(_05789_),
    .A2(_06105_),
    .B(_05801_),
    .Y(_06106_));
 NOR2x1_ASAP7_75t_SL _28522_ (.A(_06102_),
    .B(_06106_),
    .Y(_06107_));
 NOR2x1_ASAP7_75t_SL _28523_ (.A(_06100_),
    .B(_06107_),
    .Y(_06108_));
 OAI21x1_ASAP7_75t_SL _28524_ (.A1(_06108_),
    .A2(_06092_),
    .B(_05864_),
    .Y(_06109_));
 NAND2x1_ASAP7_75t_SL _28525_ (.A(_06109_),
    .B(_06072_),
    .Y(_00138_));
 OAI21x1_ASAP7_75t_SL _28526_ (.A1(_06088_),
    .A2(_06061_),
    .B(_05813_),
    .Y(_06110_));
 AOI21x1_ASAP7_75t_SL _28527_ (.A1(_05846_),
    .A2(_05984_),
    .B(_05876_),
    .Y(_06111_));
 NAND2x1_ASAP7_75t_SL _28528_ (.A(_06110_),
    .B(_06111_),
    .Y(_06112_));
 NAND2x1_ASAP7_75t_SL _28529_ (.A(_05813_),
    .B(_05949_),
    .Y(_06113_));
 NAND3x1_ASAP7_75t_SL _28530_ (.A(_06084_),
    .B(_05876_),
    .C(_06113_),
    .Y(_06114_));
 AOI21x1_ASAP7_75t_SL _28531_ (.A1(_06112_),
    .A2(_06114_),
    .B(_05844_),
    .Y(_06115_));
 NAND2x1_ASAP7_75t_SL _28532_ (.A(_05923_),
    .B(_05897_),
    .Y(_06116_));
 AOI21x1_ASAP7_75t_SL _28533_ (.A1(_05901_),
    .A2(_06116_),
    .B(_05876_),
    .Y(_06117_));
 AND2x2_ASAP7_75t_SL _28534_ (.A(_05776_),
    .B(_05888_),
    .Y(_06118_));
 AO21x1_ASAP7_75t_SL _28535_ (.A1(_05876_),
    .A2(_06118_),
    .B(_05921_),
    .Y(_06119_));
 OAI21x1_ASAP7_75t_SL _28536_ (.A1(_06117_),
    .A2(_06119_),
    .B(_05864_),
    .Y(_06120_));
 OAI21x1_ASAP7_75t_SL _28537_ (.A1(_06120_),
    .A2(_06115_),
    .B(_05855_),
    .Y(_06121_));
 AOI21x1_ASAP7_75t_SL _28538_ (.A1(_05946_),
    .A2(_06096_),
    .B(_05776_),
    .Y(_06122_));
 NOR2x1_ASAP7_75t_SL _28539_ (.A(_05892_),
    .B(_05902_),
    .Y(_06123_));
 NOR2x1_ASAP7_75t_SL _28540_ (.A(_06122_),
    .B(_06123_),
    .Y(_06124_));
 OAI21x1_ASAP7_75t_SL _28541_ (.A1(_05801_),
    .A2(_06124_),
    .B(_05789_),
    .Y(_06125_));
 AND2x2_ASAP7_75t_SL _28542_ (.A(_06003_),
    .B(_05819_),
    .Y(_06126_));
 AND2x2_ASAP7_75t_SL _28543_ (.A(_05984_),
    .B(_06035_),
    .Y(_06127_));
 OA21x2_ASAP7_75t_SL _28544_ (.A1(_06126_),
    .A2(_06127_),
    .B(_05801_),
    .Y(_06128_));
 NOR2x1p5_ASAP7_75t_SL _28545_ (.A(_06125_),
    .B(_06128_),
    .Y(_06129_));
 AND3x1_ASAP7_75t_SL _28546_ (.A(_06004_),
    .B(_05801_),
    .C(_05901_),
    .Y(_06130_));
 AND2x2_ASAP7_75t_SL _28547_ (.A(_05987_),
    .B(_05881_),
    .Y(_06131_));
 AO21x1_ASAP7_75t_SL _28548_ (.A1(_05970_),
    .A2(_05992_),
    .B(_05801_),
    .Y(_06132_));
 OAI21x1_ASAP7_75t_SL _28549_ (.A1(_06131_),
    .A2(_06132_),
    .B(_05844_),
    .Y(_06133_));
 OAI21x1_ASAP7_75t_SL _28550_ (.A1(_06130_),
    .A2(_06133_),
    .B(_06071_),
    .Y(_06134_));
 NOR2x1_ASAP7_75t_SL _28551_ (.A(_06134_),
    .B(_06129_),
    .Y(_06135_));
 NOR2x1_ASAP7_75t_SL _28552_ (.A(_06121_),
    .B(_06135_),
    .Y(_06136_));
 AOI21x1_ASAP7_75t_SL _28553_ (.A1(_06104_),
    .A2(_05889_),
    .B(_05789_),
    .Y(_06137_));
 NAND2x1_ASAP7_75t_SL _28554_ (.A(_05757_),
    .B(_05761_),
    .Y(_06138_));
 AOI21x1_ASAP7_75t_SL _28555_ (.A1(_06076_),
    .A2(_06138_),
    .B(_05776_),
    .Y(_06139_));
 INVx1_ASAP7_75t_SL _28556_ (.A(_06139_),
    .Y(_06140_));
 NAND2x1_ASAP7_75t_SL _28557_ (.A(_06140_),
    .B(_06137_),
    .Y(_06141_));
 AOI21x1_ASAP7_75t_SL _28558_ (.A1(_05896_),
    .A2(_05782_),
    .B(_05844_),
    .Y(_06142_));
 AOI21x1_ASAP7_75t_SL _28559_ (.A1(_05980_),
    .A2(_06142_),
    .B(_05801_),
    .Y(_06143_));
 AOI21x1_ASAP7_75t_SL _28560_ (.A1(_06141_),
    .A2(_06143_),
    .B(_06071_),
    .Y(_06144_));
 INVx1_ASAP7_75t_SL _28561_ (.A(_06089_),
    .Y(_06145_));
 NOR2x1_ASAP7_75t_SL _28562_ (.A(_01350_),
    .B(_05764_),
    .Y(_06146_));
 OAI21x1_ASAP7_75t_SL _28563_ (.A1(_06146_),
    .A2(_06061_),
    .B(_05813_),
    .Y(_06147_));
 AOI21x1_ASAP7_75t_SL _28564_ (.A1(_06147_),
    .A2(_06015_),
    .B(_05844_),
    .Y(_06148_));
 OAI21x1_ASAP7_75t_SL _28565_ (.A1(_06145_),
    .A2(_06148_),
    .B(_05801_),
    .Y(_06149_));
 NAND2x1_ASAP7_75t_SL _28566_ (.A(_06144_),
    .B(_06149_),
    .Y(_06150_));
 NOR2x1_ASAP7_75t_SL _28567_ (.A(_05776_),
    .B(_05757_),
    .Y(_06151_));
 AOI21x1_ASAP7_75t_SL _28568_ (.A1(_05819_),
    .A2(_05935_),
    .B(_06151_),
    .Y(_06152_));
 NAND2x1_ASAP7_75t_SL _28569_ (.A(_05789_),
    .B(_06152_),
    .Y(_06153_));
 NAND2x1_ASAP7_75t_SL _28570_ (.A(_05831_),
    .B(_06083_),
    .Y(_06154_));
 NAND2x1_ASAP7_75t_SL _28571_ (.A(_06154_),
    .B(_05961_),
    .Y(_06155_));
 AOI21x1_ASAP7_75t_SL _28572_ (.A1(_06153_),
    .A2(_06155_),
    .B(_05876_),
    .Y(_06156_));
 AND2x2_ASAP7_75t_SL _28573_ (.A(_05934_),
    .B(_05889_),
    .Y(_06157_));
 OAI21x1_ASAP7_75t_SL _28574_ (.A1(_05872_),
    .A2(_06157_),
    .B(_05876_),
    .Y(_06158_));
 AND2x2_ASAP7_75t_SL _28575_ (.A(_05959_),
    .B(_05917_),
    .Y(_06159_));
 OAI21x1_ASAP7_75t_SL _28576_ (.A1(_06008_),
    .A2(_06048_),
    .B(_05789_),
    .Y(_06160_));
 NOR2x1_ASAP7_75t_SL _28577_ (.A(_06159_),
    .B(_06160_),
    .Y(_06161_));
 NOR2x1_ASAP7_75t_SL _28578_ (.A(_06161_),
    .B(_06158_),
    .Y(_06162_));
 OAI21x1_ASAP7_75t_SL _28579_ (.A1(_06156_),
    .A2(_06162_),
    .B(_06071_),
    .Y(_06163_));
 AOI21x1_ASAP7_75t_SL _28580_ (.A1(_06150_),
    .A2(_06163_),
    .B(_05855_),
    .Y(_06164_));
 NOR2x1_ASAP7_75t_SL _28581_ (.A(_06136_),
    .B(_06164_),
    .Y(_00139_));
 NOR2x1_ASAP7_75t_R _28582_ (.A(_05757_),
    .B(_05761_),
    .Y(_06165_));
 OAI21x1_ASAP7_75t_R _28583_ (.A1(_05873_),
    .A2(_06165_),
    .B(_05813_),
    .Y(_06166_));
 AO21x1_ASAP7_75t_R _28584_ (.A1(_06166_),
    .A2(_05940_),
    .B(_05844_),
    .Y(_06167_));
 NAND2x1_ASAP7_75t_R _28585_ (.A(_05935_),
    .B(_05928_),
    .Y(_06168_));
 AOI21x1_ASAP7_75t_SL _28586_ (.A1(_05767_),
    .A2(_05887_),
    .B(_05813_),
    .Y(_06169_));
 INVx1_ASAP7_75t_SL _28587_ (.A(_06169_),
    .Y(_06170_));
 NAND2x1_ASAP7_75t_SL _28588_ (.A(_06168_),
    .B(_06170_),
    .Y(_06171_));
 AOI21x1_ASAP7_75t_R _28589_ (.A1(_05844_),
    .A2(_06171_),
    .B(_05876_),
    .Y(_06172_));
 NAND2x1_ASAP7_75t_SL _28590_ (.A(_05767_),
    .B(_05928_),
    .Y(_06173_));
 NAND2x1_ASAP7_75t_SL _28591_ (.A(_05776_),
    .B(_05908_),
    .Y(_06174_));
 NAND2x1_ASAP7_75t_R _28592_ (.A(_06173_),
    .B(_06174_),
    .Y(_06175_));
 NOR2x1_ASAP7_75t_R _28593_ (.A(_01351_),
    .B(_05813_),
    .Y(_06176_));
 AO21x1_ASAP7_75t_SL _28594_ (.A1(_05813_),
    .A2(_05916_),
    .B(_05844_),
    .Y(_06177_));
 OAI21x1_ASAP7_75t_R _28595_ (.A1(_06176_),
    .A2(_06177_),
    .B(_05876_),
    .Y(_06178_));
 AOI21x1_ASAP7_75t_R _28596_ (.A1(_05844_),
    .A2(_06175_),
    .B(_06178_),
    .Y(_06179_));
 AOI21x1_ASAP7_75t_R _28597_ (.A1(_06167_),
    .A2(_06172_),
    .B(_06179_),
    .Y(_06180_));
 AOI21x1_ASAP7_75t_R _28598_ (.A1(_05810_),
    .A2(_05840_),
    .B(_05789_),
    .Y(_06181_));
 AO21x1_ASAP7_75t_SL _28599_ (.A1(_05810_),
    .A2(_05970_),
    .B(_05813_),
    .Y(_06182_));
 NAND2x1_ASAP7_75t_SL _28600_ (.A(_06181_),
    .B(_06182_),
    .Y(_06183_));
 AOI21x1_ASAP7_75t_R _28601_ (.A1(_06104_),
    .A2(_06003_),
    .B(_05977_),
    .Y(_06184_));
 AOI21x1_ASAP7_75t_R _28602_ (.A1(_05789_),
    .A2(_06184_),
    .B(_05876_),
    .Y(_06185_));
 NAND2x1_ASAP7_75t_SL _28603_ (.A(_06183_),
    .B(_06185_),
    .Y(_06186_));
 OAI21x1_ASAP7_75t_R _28604_ (.A1(_05761_),
    .A2(_05769_),
    .B(_05813_),
    .Y(_06187_));
 AOI21x1_ASAP7_75t_SL _28605_ (.A1(_01345_),
    .A2(_05757_),
    .B(_05813_),
    .Y(_06188_));
 NOR2x1_ASAP7_75t_R _28606_ (.A(_05789_),
    .B(_06188_),
    .Y(_06189_));
 AOI21x1_ASAP7_75t_R _28607_ (.A1(_06187_),
    .A2(_06189_),
    .B(_05801_),
    .Y(_06190_));
 AOI21x1_ASAP7_75t_R _28608_ (.A1(_06103_),
    .A2(_05938_),
    .B(_05844_),
    .Y(_06191_));
 NAND2x1_ASAP7_75t_SL _28609_ (.A(_06191_),
    .B(_05807_),
    .Y(_06192_));
 AOI21x1_ASAP7_75t_SL _28610_ (.A1(_06190_),
    .A2(_06192_),
    .B(_05855_),
    .Y(_06193_));
 AOI21x1_ASAP7_75t_SL _28611_ (.A1(_06193_),
    .A2(_06186_),
    .B(_06071_),
    .Y(_06194_));
 OAI21x1_ASAP7_75t_SL _28612_ (.A1(_05856_),
    .A2(_06180_),
    .B(_06194_),
    .Y(_06195_));
 NAND2x1_ASAP7_75t_R _28613_ (.A(_06004_),
    .B(_06045_),
    .Y(_06196_));
 AND2x2_ASAP7_75t_R _28614_ (.A(_06044_),
    .B(_05884_),
    .Y(_06197_));
 OAI21x1_ASAP7_75t_R _28615_ (.A1(_06169_),
    .A2(_06197_),
    .B(_05844_),
    .Y(_06198_));
 AOI21x1_ASAP7_75t_R _28616_ (.A1(_06196_),
    .A2(_06198_),
    .B(_05876_),
    .Y(_06199_));
 AO22x1_ASAP7_75t_L _28617_ (.A1(_05823_),
    .A2(_06006_),
    .B1(_05996_),
    .B2(_05972_),
    .Y(_06200_));
 OAI21x1_ASAP7_75t_R _28618_ (.A1(_05811_),
    .A2(_05928_),
    .B(_05844_),
    .Y(_06201_));
 NAND2x1_ASAP7_75t_R _28619_ (.A(_05876_),
    .B(_06201_),
    .Y(_06202_));
 AOI21x1_ASAP7_75t_R _28620_ (.A1(_05789_),
    .A2(_06200_),
    .B(_06202_),
    .Y(_06203_));
 OAI21x1_ASAP7_75t_R _28621_ (.A1(_06199_),
    .A2(_06203_),
    .B(_05856_),
    .Y(_06204_));
 NAND2x1_ASAP7_75t_L _28622_ (.A(_06035_),
    .B(_05896_),
    .Y(_06205_));
 AOI21x1_ASAP7_75t_SL _28623_ (.A1(_06205_),
    .A2(_05909_),
    .B(_05844_),
    .Y(_06206_));
 AO21x1_ASAP7_75t_R _28624_ (.A1(_05834_),
    .A2(_05966_),
    .B(_05813_),
    .Y(_06207_));
 OAI21x1_ASAP7_75t_R _28625_ (.A1(_05841_),
    .A2(_05908_),
    .B(_05813_),
    .Y(_06208_));
 AOI21x1_ASAP7_75t_R _28626_ (.A1(_06207_),
    .A2(_06208_),
    .B(_05789_),
    .Y(_06209_));
 OAI21x1_ASAP7_75t_R _28627_ (.A1(_06206_),
    .A2(_06209_),
    .B(_05801_),
    .Y(_06210_));
 AO21x1_ASAP7_75t_SL _28628_ (.A1(_05907_),
    .A2(_05776_),
    .B(_05789_),
    .Y(_06211_));
 AO21x1_ASAP7_75t_SL _28629_ (.A1(_05813_),
    .A2(_05916_),
    .B(_05949_),
    .Y(_06212_));
 OA21x2_ASAP7_75t_R _28630_ (.A1(_06211_),
    .A2(_06212_),
    .B(_05876_),
    .Y(_06213_));
 OAI21x1_ASAP7_75t_R _28631_ (.A1(_05757_),
    .A2(_05819_),
    .B(_05928_),
    .Y(_06214_));
 INVx1_ASAP7_75t_SL _28632_ (.A(_05900_),
    .Y(_06215_));
 NAND2x1_ASAP7_75t_SL _28633_ (.A(_06019_),
    .B(_06215_),
    .Y(_06216_));
 NAND3x1_ASAP7_75t_SL _28634_ (.A(_06216_),
    .B(_05789_),
    .C(_06214_),
    .Y(_06217_));
 AOI21x1_ASAP7_75t_SL _28635_ (.A1(_06217_),
    .A2(_06213_),
    .B(_05856_),
    .Y(_06218_));
 AOI21x1_ASAP7_75t_SL _28636_ (.A1(_06218_),
    .A2(_06210_),
    .B(_05864_),
    .Y(_06219_));
 NAND2x1_ASAP7_75t_SL _28637_ (.A(_06204_),
    .B(_06219_),
    .Y(_06220_));
 NAND2x1_ASAP7_75t_SL _28638_ (.A(_06195_),
    .B(_06220_),
    .Y(_00140_));
 NOR2x1_ASAP7_75t_SL _28639_ (.A(_05880_),
    .B(_05776_),
    .Y(_06221_));
 AO21x1_ASAP7_75t_SL _28640_ (.A1(_06221_),
    .A2(_05757_),
    .B(_05789_),
    .Y(_06222_));
 NOR2x1_ASAP7_75t_R _28641_ (.A(_05813_),
    .B(_05737_),
    .Y(_06223_));
 OA21x2_ASAP7_75t_SL _28642_ (.A1(_05937_),
    .A2(_06223_),
    .B(_06104_),
    .Y(_06224_));
 OAI21x1_ASAP7_75t_SL _28643_ (.A1(_06222_),
    .A2(_06224_),
    .B(_05801_),
    .Y(_06225_));
 AO21x1_ASAP7_75t_SL _28644_ (.A1(_05935_),
    .A2(_05946_),
    .B(_05813_),
    .Y(_06226_));
 AND3x1_ASAP7_75t_SL _28645_ (.A(_06226_),
    .B(_05807_),
    .C(_05789_),
    .Y(_06227_));
 NOR2x1_ASAP7_75t_SL _28646_ (.A(_06225_),
    .B(_06227_),
    .Y(_06228_));
 AOI211x1_ASAP7_75t_SL _28647_ (.A1(_05737_),
    .A2(_05813_),
    .B(_05875_),
    .C(_05844_),
    .Y(_06229_));
 AO21x1_ASAP7_75t_SL _28648_ (.A1(_06083_),
    .A2(_05767_),
    .B(_05789_),
    .Y(_06230_));
 AND2x2_ASAP7_75t_SL _28649_ (.A(_05951_),
    .B(_05842_),
    .Y(_06231_));
 OAI21x1_ASAP7_75t_SL _28650_ (.A1(_06231_),
    .A2(_06230_),
    .B(_05876_),
    .Y(_06232_));
 OAI21x1_ASAP7_75t_SL _28651_ (.A1(_06232_),
    .A2(_06229_),
    .B(_05856_),
    .Y(_06233_));
 NOR2x1_ASAP7_75t_SL _28652_ (.A(_06228_),
    .B(_06233_),
    .Y(_06234_));
 OAI21x1_ASAP7_75t_SL _28653_ (.A1(_05960_),
    .A2(_06211_),
    .B(_05876_),
    .Y(_06235_));
 AOI21x1_ASAP7_75t_SL _28654_ (.A1(_05737_),
    .A2(_05805_),
    .B(_05813_),
    .Y(_06236_));
 AND3x1_ASAP7_75t_R _28655_ (.A(_05756_),
    .B(_05747_),
    .C(_06060_),
    .Y(_06237_));
 OAI21x1_ASAP7_75t_SL _28656_ (.A1(_05776_),
    .A2(_06237_),
    .B(_05789_),
    .Y(_06238_));
 AOI21x1_ASAP7_75t_SL _28657_ (.A1(_05842_),
    .A2(_06236_),
    .B(_06238_),
    .Y(_06239_));
 OAI21x1_ASAP7_75t_SL _28658_ (.A1(_06235_),
    .A2(_06239_),
    .B(_05855_),
    .Y(_06240_));
 OAI21x1_ASAP7_75t_SL _28659_ (.A1(_06221_),
    .A2(_06236_),
    .B(_05789_),
    .Y(_06241_));
 AOI21x1_ASAP7_75t_SL _28660_ (.A1(_05831_),
    .A2(_05934_),
    .B(_05776_),
    .Y(_06242_));
 OA21x2_ASAP7_75t_SL _28661_ (.A1(_05888_),
    .A2(_06088_),
    .B(_05776_),
    .Y(_06243_));
 OAI21x1_ASAP7_75t_SL _28662_ (.A1(_06242_),
    .A2(_06243_),
    .B(_05844_),
    .Y(_06244_));
 AOI21x1_ASAP7_75t_SL _28663_ (.A1(_06241_),
    .A2(_06244_),
    .B(_05876_),
    .Y(_06245_));
 OAI21x1_ASAP7_75t_SL _28664_ (.A1(_06240_),
    .A2(_06245_),
    .B(_05864_),
    .Y(_06246_));
 AOI211x1_ASAP7_75t_SL _28665_ (.A1(_05819_),
    .A2(_05977_),
    .B(_05789_),
    .C(_06103_),
    .Y(_06247_));
 AO21x1_ASAP7_75t_SL _28666_ (.A1(_05776_),
    .A2(_05984_),
    .B(_05844_),
    .Y(_06248_));
 OAI21x1_ASAP7_75t_SL _28667_ (.A1(_06139_),
    .A2(_06248_),
    .B(_05801_),
    .Y(_06249_));
 OAI21x1_ASAP7_75t_SL _28668_ (.A1(_06249_),
    .A2(_06247_),
    .B(_05856_),
    .Y(_06250_));
 NOR2x1_ASAP7_75t_SL _28669_ (.A(_01347_),
    .B(_05776_),
    .Y(_06251_));
 AOI211x1_ASAP7_75t_SL _28670_ (.A1(_05927_),
    .A2(_06083_),
    .B(_05921_),
    .C(_06251_),
    .Y(_06252_));
 AOI21x1_ASAP7_75t_SL _28671_ (.A1(_01342_),
    .A2(_05757_),
    .B(_05811_),
    .Y(_06253_));
 AO21x1_ASAP7_75t_SL _28672_ (.A1(_05834_),
    .A2(_05966_),
    .B(_05776_),
    .Y(_06254_));
 OAI21x1_ASAP7_75t_SL _28673_ (.A1(_05813_),
    .A2(_06253_),
    .B(_06254_),
    .Y(_06255_));
 OAI21x1_ASAP7_75t_SL _28674_ (.A1(_05844_),
    .A2(_06255_),
    .B(_05876_),
    .Y(_06256_));
 NOR2x1_ASAP7_75t_SL _28675_ (.A(_06252_),
    .B(_06256_),
    .Y(_06257_));
 NOR2x1_ASAP7_75t_SL _28676_ (.A(_06257_),
    .B(_06250_),
    .Y(_06258_));
 NAND2x1p5_ASAP7_75t_SL _28677_ (.A(_05951_),
    .B(_05884_),
    .Y(_06259_));
 AOI21x1_ASAP7_75t_SL _28678_ (.A1(_06079_),
    .A2(_06259_),
    .B(_05844_),
    .Y(_06260_));
 AO21x1_ASAP7_75t_SL _28679_ (.A1(_05916_),
    .A2(_05813_),
    .B(_05789_),
    .Y(_06261_));
 AND2x2_ASAP7_75t_SL _28680_ (.A(_06188_),
    .B(_05923_),
    .Y(_06262_));
 OAI21x1_ASAP7_75t_SL _28681_ (.A1(_06261_),
    .A2(_06262_),
    .B(_05801_),
    .Y(_06263_));
 OAI21x1_ASAP7_75t_SL _28682_ (.A1(_06263_),
    .A2(_06260_),
    .B(_05855_),
    .Y(_06264_));
 OA21x2_ASAP7_75t_SL _28683_ (.A1(_05722_),
    .A2(_05776_),
    .B(_05789_),
    .Y(_06265_));
 NAND2x1_ASAP7_75t_SL _28684_ (.A(_06265_),
    .B(_06170_),
    .Y(_06266_));
 NAND2x1_ASAP7_75t_SL _28685_ (.A(_05934_),
    .B(_05959_),
    .Y(_06267_));
 AOI21x1_ASAP7_75t_SL _28686_ (.A1(_05887_),
    .A2(_05846_),
    .B(_05789_),
    .Y(_06268_));
 OAI21x1_ASAP7_75t_SL _28687_ (.A1(_05776_),
    .A2(_06267_),
    .B(_06268_),
    .Y(_06269_));
 AOI21x1_ASAP7_75t_SL _28688_ (.A1(_06266_),
    .A2(_06269_),
    .B(_05801_),
    .Y(_06270_));
 OAI21x1_ASAP7_75t_SL _28689_ (.A1(_06270_),
    .A2(_06264_),
    .B(_06071_),
    .Y(_06271_));
 OAI22x1_ASAP7_75t_SL _28690_ (.A1(_06234_),
    .A2(_06246_),
    .B1(_06271_),
    .B2(_06258_),
    .Y(_00141_));
 NOR2x1_ASAP7_75t_R _28691_ (.A(_05789_),
    .B(_05897_),
    .Y(_06272_));
 AOI21x1_ASAP7_75t_SL _28692_ (.A1(_06173_),
    .A2(_06272_),
    .B(_05876_),
    .Y(_06273_));
 OR4x1_ASAP7_75t_L _28693_ (.A(_05908_),
    .B(_05776_),
    .C(_05844_),
    .D(_05907_),
    .Y(_06274_));
 AOI21x1_ASAP7_75t_R _28694_ (.A1(_06273_),
    .A2(_06274_),
    .B(_06071_),
    .Y(_06275_));
 AND2x2_ASAP7_75t_SL _28695_ (.A(_06083_),
    .B(_05767_),
    .Y(_06276_));
 AO21x1_ASAP7_75t_R _28696_ (.A1(_01355_),
    .A2(_05813_),
    .B(_05844_),
    .Y(_06277_));
 OA21x2_ASAP7_75t_R _28697_ (.A1(_06276_),
    .A2(_06277_),
    .B(_05876_),
    .Y(_06278_));
 AO21x1_ASAP7_75t_R _28698_ (.A1(_05831_),
    .A2(_05960_),
    .B(_06027_),
    .Y(_06279_));
 NAND2x1_ASAP7_75t_R _28699_ (.A(_06278_),
    .B(_06279_),
    .Y(_06280_));
 NAND2x1_ASAP7_75t_SL _28700_ (.A(_06275_),
    .B(_06280_),
    .Y(_06281_));
 AOI21x1_ASAP7_75t_SL _28701_ (.A1(_06053_),
    .A2(_05778_),
    .B(_05903_),
    .Y(_06282_));
 INVx1_ASAP7_75t_R _28702_ (.A(_06188_),
    .Y(_06283_));
 OAI21x1_ASAP7_75t_R _28703_ (.A1(_05805_),
    .A2(_06008_),
    .B(_05813_),
    .Y(_06284_));
 AO21x1_ASAP7_75t_R _28704_ (.A1(_05892_),
    .A2(_05776_),
    .B(_05844_),
    .Y(_06285_));
 AOI21x1_ASAP7_75t_R _28705_ (.A1(_06283_),
    .A2(_06284_),
    .B(_06285_),
    .Y(_06286_));
 OAI21x1_ASAP7_75t_SL _28706_ (.A1(_06286_),
    .A2(_06282_),
    .B(_05876_),
    .Y(_06287_));
 NAND2x1_ASAP7_75t_SL _28707_ (.A(_05819_),
    .B(_05996_),
    .Y(_06288_));
 OA21x2_ASAP7_75t_R _28708_ (.A1(_05934_),
    .A2(_05813_),
    .B(_05844_),
    .Y(_06289_));
 AOI21x1_ASAP7_75t_R _28709_ (.A1(_06288_),
    .A2(_06289_),
    .B(_05876_),
    .Y(_06290_));
 AOI21x1_ASAP7_75t_R _28710_ (.A1(_05761_),
    .A2(_05977_),
    .B(_05844_),
    .Y(_06291_));
 OAI21x1_ASAP7_75t_R _28711_ (.A1(_05900_),
    .A2(_06061_),
    .B(_05776_),
    .Y(_06292_));
 NAND3x1_ASAP7_75t_SL _28712_ (.A(_06166_),
    .B(_06291_),
    .C(_06292_),
    .Y(_06293_));
 AOI21x1_ASAP7_75t_R _28713_ (.A1(_06290_),
    .A2(_06293_),
    .B(_05864_),
    .Y(_06294_));
 AOI21x1_ASAP7_75t_SL _28714_ (.A1(_06294_),
    .A2(_06287_),
    .B(_05856_),
    .Y(_06295_));
 NAND2x1_ASAP7_75t_SL _28715_ (.A(_06295_),
    .B(_06281_),
    .Y(_06296_));
 AOI21x1_ASAP7_75t_R _28716_ (.A1(_05784_),
    .A2(_06083_),
    .B(_05876_),
    .Y(_06297_));
 OAI21x1_ASAP7_75t_R _28717_ (.A1(_05811_),
    .A2(_05963_),
    .B(_05813_),
    .Y(_06298_));
 NAND2x1_ASAP7_75t_SL _28718_ (.A(_06297_),
    .B(_06298_),
    .Y(_06299_));
 NAND2x1_ASAP7_75t_SL _28719_ (.A(_05819_),
    .B(_06035_),
    .Y(_06300_));
 AO21x1_ASAP7_75t_R _28720_ (.A1(_01354_),
    .A2(_01360_),
    .B(_05813_),
    .Y(_06301_));
 NAND3x1_ASAP7_75t_R _28721_ (.A(_06300_),
    .B(_05876_),
    .C(_06301_),
    .Y(_06302_));
 AOI21x1_ASAP7_75t_SL _28722_ (.A1(_06299_),
    .A2(_06302_),
    .B(_05844_),
    .Y(_06303_));
 NOR2x1_ASAP7_75t_R _28723_ (.A(_05801_),
    .B(_06066_),
    .Y(_06304_));
 NAND2x1_ASAP7_75t_R _28724_ (.A(_06113_),
    .B(_06304_),
    .Y(_06305_));
 AND2x2_ASAP7_75t_R _28725_ (.A(_06113_),
    .B(_05801_),
    .Y(_06306_));
 NAND2x1_ASAP7_75t_SL _28726_ (.A(_05935_),
    .B(_05917_),
    .Y(_06307_));
 NAND2x1_ASAP7_75t_R _28727_ (.A(_05813_),
    .B(_05907_),
    .Y(_06308_));
 NAND3x1_ASAP7_75t_R _28728_ (.A(_06306_),
    .B(_06307_),
    .C(_06308_),
    .Y(_06309_));
 AO21x1_ASAP7_75t_R _28729_ (.A1(_05913_),
    .A2(_05813_),
    .B(_05789_),
    .Y(_06310_));
 AOI21x1_ASAP7_75t_SL _28730_ (.A1(_06305_),
    .A2(_06309_),
    .B(_06310_),
    .Y(_06311_));
 OAI21x1_ASAP7_75t_R _28731_ (.A1(_06303_),
    .A2(_06311_),
    .B(_06071_),
    .Y(_06312_));
 OAI21x1_ASAP7_75t_R _28732_ (.A1(_05776_),
    .A2(_05841_),
    .B(_05825_),
    .Y(_06313_));
 OA21x2_ASAP7_75t_R _28733_ (.A1(_06139_),
    .A2(_06285_),
    .B(_05801_),
    .Y(_06314_));
 AOI21x1_ASAP7_75t_R _28734_ (.A1(_06313_),
    .A2(_06314_),
    .B(_06071_),
    .Y(_06315_));
 NAND2x1_ASAP7_75t_R _28735_ (.A(_05867_),
    .B(_06019_),
    .Y(_06316_));
 AO21x1_ASAP7_75t_R _28736_ (.A1(_05935_),
    .A2(_05819_),
    .B(_05776_),
    .Y(_06317_));
 AOI21x1_ASAP7_75t_R _28737_ (.A1(_06316_),
    .A2(_06317_),
    .B(_05789_),
    .Y(_06318_));
 NAND2x1_ASAP7_75t_R _28738_ (.A(_05776_),
    .B(_06055_),
    .Y(_06319_));
 AO21x1_ASAP7_75t_R _28739_ (.A1(_05867_),
    .A2(_05979_),
    .B(_05776_),
    .Y(_06320_));
 AOI21x1_ASAP7_75t_R _28740_ (.A1(_06319_),
    .A2(_06320_),
    .B(_05844_),
    .Y(_06321_));
 OAI21x1_ASAP7_75t_R _28741_ (.A1(_06318_),
    .A2(_06321_),
    .B(_05876_),
    .Y(_06322_));
 AOI21x1_ASAP7_75t_R _28742_ (.A1(_06315_),
    .A2(_06322_),
    .B(_05855_),
    .Y(_06323_));
 NAND2x1_ASAP7_75t_SL _28743_ (.A(_06312_),
    .B(_06323_),
    .Y(_06324_));
 NAND2x1_ASAP7_75t_SL _28744_ (.A(_06324_),
    .B(_06296_),
    .Y(_00142_));
 OAI21x1_ASAP7_75t_R _28745_ (.A1(_05761_),
    .A2(_05769_),
    .B(_05896_),
    .Y(_06325_));
 NOR2x1_ASAP7_75t_R _28746_ (.A(_05776_),
    .B(_06325_),
    .Y(_06326_));
 NAND2x1_ASAP7_75t_R _28747_ (.A(_06174_),
    .B(_06026_),
    .Y(_06327_));
 NOR2x1_ASAP7_75t_R _28748_ (.A(_05844_),
    .B(_06019_),
    .Y(_06328_));
 AOI21x1_ASAP7_75t_R _28749_ (.A1(_06173_),
    .A2(_06328_),
    .B(_05801_),
    .Y(_06329_));
 OAI21x1_ASAP7_75t_R _28750_ (.A1(_06326_),
    .A2(_06327_),
    .B(_06329_),
    .Y(_06330_));
 NAND2x1_ASAP7_75t_R _28751_ (.A(_05784_),
    .B(_06083_),
    .Y(_06331_));
 AOI21x1_ASAP7_75t_R _28752_ (.A1(_06036_),
    .A2(_06331_),
    .B(_05844_),
    .Y(_06332_));
 NAND2x1_ASAP7_75t_R _28753_ (.A(_05784_),
    .B(_05992_),
    .Y(_06333_));
 NAND2x1_ASAP7_75t_L _28754_ (.A(_05984_),
    .B(_05846_),
    .Y(_06334_));
 AOI21x1_ASAP7_75t_SL _28755_ (.A1(_06333_),
    .A2(_06334_),
    .B(_05789_),
    .Y(_06335_));
 OAI21x1_ASAP7_75t_SL _28756_ (.A1(_06335_),
    .A2(_06332_),
    .B(_05801_),
    .Y(_06336_));
 AOI21x1_ASAP7_75t_SL _28757_ (.A1(_06336_),
    .A2(_06330_),
    .B(_05855_),
    .Y(_06337_));
 AO21x1_ASAP7_75t_SL _28758_ (.A1(_05996_),
    .A2(_05972_),
    .B(_06223_),
    .Y(_06338_));
 NAND2x1_ASAP7_75t_R _28759_ (.A(_05844_),
    .B(_06338_),
    .Y(_06339_));
 OAI21x1_ASAP7_75t_R _28760_ (.A1(_05805_),
    .A2(_05963_),
    .B(_05776_),
    .Y(_06340_));
 AOI21x1_ASAP7_75t_R _28761_ (.A1(_06045_),
    .A2(_06340_),
    .B(_05801_),
    .Y(_06341_));
 NAND2x1_ASAP7_75t_SL _28762_ (.A(_06339_),
    .B(_06341_),
    .Y(_06342_));
 OAI21x1_ASAP7_75t_R _28763_ (.A1(_05888_),
    .A2(_05963_),
    .B(_05776_),
    .Y(_06343_));
 AO21x1_ASAP7_75t_R _28764_ (.A1(_05805_),
    .A2(_05761_),
    .B(_05776_),
    .Y(_06344_));
 NAND2x1_ASAP7_75t_SL _28765_ (.A(_06343_),
    .B(_06344_),
    .Y(_06345_));
 NAND2x1_ASAP7_75t_R _28766_ (.A(_06151_),
    .B(_05887_),
    .Y(_06346_));
 AOI21x1_ASAP7_75t_SL _28767_ (.A1(_05888_),
    .A2(_05776_),
    .B(_05844_),
    .Y(_06347_));
 AOI21x1_ASAP7_75t_SL _28768_ (.A1(_06347_),
    .A2(_06346_),
    .B(_05876_),
    .Y(_06348_));
 OAI21x1_ASAP7_75t_R _28769_ (.A1(_05789_),
    .A2(_06345_),
    .B(_06348_),
    .Y(_06349_));
 AOI21x1_ASAP7_75t_R _28770_ (.A1(_06342_),
    .A2(_06349_),
    .B(_05856_),
    .Y(_06350_));
 OAI21x1_ASAP7_75t_SL _28771_ (.A1(_06337_),
    .A2(_06350_),
    .B(_05864_),
    .Y(_06351_));
 AND2x2_ASAP7_75t_SL _28772_ (.A(_05846_),
    .B(_05767_),
    .Y(_06352_));
 AO21x1_ASAP7_75t_R _28773_ (.A1(_05992_),
    .A2(_05831_),
    .B(_05789_),
    .Y(_06353_));
 NAND2x1_ASAP7_75t_R _28774_ (.A(_01360_),
    .B(_05813_),
    .Y(_06354_));
 OAI21x1_ASAP7_75t_R _28775_ (.A1(_05813_),
    .A2(_05900_),
    .B(_06354_),
    .Y(_06355_));
 AOI21x1_ASAP7_75t_R _28776_ (.A1(_05776_),
    .A2(_05949_),
    .B(_05844_),
    .Y(_06356_));
 AOI21x1_ASAP7_75t_R _28777_ (.A1(_06355_),
    .A2(_06356_),
    .B(_05876_),
    .Y(_06357_));
 OAI21x1_ASAP7_75t_R _28778_ (.A1(_06352_),
    .A2(_06353_),
    .B(_06357_),
    .Y(_06358_));
 INVx1_ASAP7_75t_R _28779_ (.A(_06181_),
    .Y(_06359_));
 AND3x1_ASAP7_75t_R _28780_ (.A(_05819_),
    .B(_05776_),
    .C(_05769_),
    .Y(_06360_));
 NAND2x1_ASAP7_75t_R _28781_ (.A(_01351_),
    .B(_05813_),
    .Y(_06361_));
 AOI21x1_ASAP7_75t_R _28782_ (.A1(_06361_),
    .A2(_05914_),
    .B(_05801_),
    .Y(_06362_));
 OAI21x1_ASAP7_75t_R _28783_ (.A1(_06359_),
    .A2(_06360_),
    .B(_06362_),
    .Y(_06363_));
 AOI21x1_ASAP7_75t_R _28784_ (.A1(_06358_),
    .A2(_06363_),
    .B(_05856_),
    .Y(_06364_));
 NAND2x1p5_ASAP7_75t_SL _28785_ (.A(_05951_),
    .B(_05934_),
    .Y(_06365_));
 AOI21x1_ASAP7_75t_R _28786_ (.A1(_05776_),
    .A2(_06325_),
    .B(_05844_),
    .Y(_06366_));
 NAND2x1_ASAP7_75t_R _28787_ (.A(_05887_),
    .B(_05937_),
    .Y(_06367_));
 AOI21x1_ASAP7_75t_R _28788_ (.A1(_06367_),
    .A2(_06147_),
    .B(_05789_),
    .Y(_06368_));
 AOI21x1_ASAP7_75t_SL _28789_ (.A1(_06366_),
    .A2(_06365_),
    .B(_06368_),
    .Y(_06369_));
 NAND2x1_ASAP7_75t_R _28790_ (.A(_05945_),
    .B(_05776_),
    .Y(_06370_));
 AOI21x1_ASAP7_75t_R _28791_ (.A1(_06370_),
    .A2(_06300_),
    .B(_05789_),
    .Y(_06371_));
 NAND2x1_ASAP7_75t_R _28792_ (.A(_05789_),
    .B(_05896_),
    .Y(_06372_));
 NOR2x1_ASAP7_75t_SL _28793_ (.A(_05996_),
    .B(_06188_),
    .Y(_06373_));
 OAI21x1_ASAP7_75t_SL _28794_ (.A1(_06372_),
    .A2(_06373_),
    .B(_05801_),
    .Y(_06374_));
 OAI21x1_ASAP7_75t_R _28795_ (.A1(_06371_),
    .A2(_06374_),
    .B(_05856_),
    .Y(_06375_));
 AOI21x1_ASAP7_75t_SL _28796_ (.A1(_05876_),
    .A2(_06369_),
    .B(_06375_),
    .Y(_06376_));
 OAI21x1_ASAP7_75t_SL _28797_ (.A1(_06364_),
    .A2(_06376_),
    .B(_06071_),
    .Y(_06377_));
 NAND2x1_ASAP7_75t_SL _28798_ (.A(_06351_),
    .B(_06377_),
    .Y(_00143_));
 NOR2x1_ASAP7_75t_L _28799_ (.A(_00574_),
    .B(_00405_),
    .Y(_06378_));
 XOR2x2_ASAP7_75t_SL _28800_ (.A(_03677_),
    .B(_12118_),
    .Y(_06379_));
 XOR2x2_ASAP7_75t_SL _28801_ (.A(_12078_),
    .B(_00656_),
    .Y(_06380_));
 INVx1_ASAP7_75t_R _28802_ (.A(_06380_),
    .Y(_06381_));
 NAND2x1_ASAP7_75t_L _28803_ (.A(_06379_),
    .B(_06381_),
    .Y(_06382_));
 INVx2_ASAP7_75t_SL _28804_ (.A(_06379_),
    .Y(_06383_));
 NAND2x1p5_ASAP7_75t_SL _28805_ (.A(_06383_),
    .B(_06380_),
    .Y(_06384_));
 AOI21x1_ASAP7_75t_SL _28806_ (.A1(_06384_),
    .A2(_06382_),
    .B(_10675_),
    .Y(_06385_));
 OAI21x1_ASAP7_75t_R _28807_ (.A1(_06378_),
    .A2(_06385_),
    .B(_00913_),
    .Y(_06386_));
 AND2x2_ASAP7_75t_R _28808_ (.A(_10675_),
    .B(_00405_),
    .Y(_06387_));
 XOR2x1_ASAP7_75t_SL _28809_ (.A(_06380_),
    .Y(_06388_),
    .B(_06379_));
 NOR2x1p5_ASAP7_75t_SL _28810_ (.A(_10675_),
    .B(_06388_),
    .Y(_06389_));
 INVx1_ASAP7_75t_R _28811_ (.A(_00913_),
    .Y(_06390_));
 OAI21x1_ASAP7_75t_R _28812_ (.A1(_06387_),
    .A2(_06389_),
    .B(_06390_),
    .Y(_06391_));
 NAND2x1_ASAP7_75t_SL _28813_ (.A(_06386_),
    .B(_06391_),
    .Y(_06392_));
 OR2x2_ASAP7_75t_R _28816_ (.A(_00574_),
    .B(_00406_),
    .Y(_06394_));
 XOR2x2_ASAP7_75t_SL _28817_ (.A(_12102_),
    .B(_12268_),
    .Y(_06395_));
 NOR2x1_ASAP7_75t_R _28818_ (.A(_12084_),
    .B(_06395_),
    .Y(_06396_));
 AND2x2_ASAP7_75t_R _28819_ (.A(_06395_),
    .B(_12084_),
    .Y(_06397_));
 OAI21x1_ASAP7_75t_SL _28820_ (.A1(_06396_),
    .A2(_06397_),
    .B(_00574_),
    .Y(_06398_));
 AOI21x1_ASAP7_75t_R _28821_ (.A1(_06394_),
    .A2(_06398_),
    .B(_00902_),
    .Y(_06399_));
 NAND2x1_ASAP7_75t_L _28822_ (.A(_00406_),
    .B(_10675_),
    .Y(_06400_));
 XOR2x2_ASAP7_75t_SL _28823_ (.A(_06395_),
    .B(_12084_),
    .Y(_06401_));
 NAND2x1p5_ASAP7_75t_L _28824_ (.A(_00574_),
    .B(_06401_),
    .Y(_06402_));
 INVx1_ASAP7_75t_R _28825_ (.A(_00902_),
    .Y(_06403_));
 AOI21x1_ASAP7_75t_R _28826_ (.A1(_06400_),
    .A2(_06402_),
    .B(_06403_),
    .Y(_06404_));
 NOR2x2_ASAP7_75t_SL _28827_ (.A(_06399_),
    .B(_06404_),
    .Y(_06405_));
 NOR2x1_ASAP7_75t_R _28829_ (.A(_00574_),
    .B(_00407_),
    .Y(_06406_));
 XOR2x2_ASAP7_75t_SL _28830_ (.A(_00592_),
    .B(_00657_),
    .Y(_06407_));
 NAND2x1_ASAP7_75t_L _28831_ (.A(_12082_),
    .B(_06407_),
    .Y(_06408_));
 XNOR2x2_ASAP7_75t_L _28832_ (.A(_00592_),
    .B(_00657_),
    .Y(_06409_));
 NAND2x1_ASAP7_75t_R _28833_ (.A(_00688_),
    .B(_06409_),
    .Y(_06410_));
 AOI21x1_ASAP7_75t_SL _28834_ (.A1(_06408_),
    .A2(_06410_),
    .B(_03707_),
    .Y(_06411_));
 INVx1_ASAP7_75t_SL _28835_ (.A(_06411_),
    .Y(_06412_));
 NAND3x1_ASAP7_75t_L _28836_ (.A(_06410_),
    .B(_06408_),
    .C(_03707_),
    .Y(_06413_));
 AOI21x1_ASAP7_75t_SL _28837_ (.A1(_06412_),
    .A2(_06413_),
    .B(_10675_),
    .Y(_06414_));
 OAI21x1_ASAP7_75t_SL _28838_ (.A1(_06406_),
    .A2(_06414_),
    .B(_08790_),
    .Y(_06415_));
 XOR2x2_ASAP7_75t_SL _28839_ (.A(_06407_),
    .B(_00688_),
    .Y(_06416_));
 NOR2x1_ASAP7_75t_R _28840_ (.A(_03706_),
    .B(_06416_),
    .Y(_06417_));
 OAI21x1_ASAP7_75t_L _28841_ (.A1(_06411_),
    .A2(_06417_),
    .B(_00574_),
    .Y(_06418_));
 INVx1_ASAP7_75t_R _28842_ (.A(_06406_),
    .Y(_06419_));
 NAND3x1_ASAP7_75t_SL _28843_ (.A(_06418_),
    .B(_00924_),
    .C(_06419_),
    .Y(_06420_));
 NAND2x2_ASAP7_75t_SL _28844_ (.A(_06415_),
    .B(_06420_),
    .Y(_06421_));
 AOI21x1_ASAP7_75t_SL _28846_ (.A1(_06394_),
    .A2(_06398_),
    .B(_06403_),
    .Y(_06422_));
 AOI21x1_ASAP7_75t_R _28847_ (.A1(_06400_),
    .A2(_06402_),
    .B(_00902_),
    .Y(_06423_));
 NOR2x1_ASAP7_75t_SL _28848_ (.A(_06422_),
    .B(_06423_),
    .Y(_06424_));
 OAI21x1_ASAP7_75t_SL _28851_ (.A1(_06406_),
    .A2(_06414_),
    .B(_00924_),
    .Y(_06426_));
 NAND3x1_ASAP7_75t_SL _28852_ (.A(_06418_),
    .B(_08790_),
    .C(_06419_),
    .Y(_06427_));
 NAND2x2_ASAP7_75t_SL _28853_ (.A(_06426_),
    .B(_06427_),
    .Y(_06428_));
 XOR2x2_ASAP7_75t_L _28855_ (.A(_12161_),
    .B(_00659_),
    .Y(_06429_));
 XOR2x2_ASAP7_75t_SL _28856_ (.A(_03758_),
    .B(_06429_),
    .Y(_06430_));
 NOR2x1_ASAP7_75t_R _28857_ (.A(_00574_),
    .B(_00533_),
    .Y(_06431_));
 AOI21x1_ASAP7_75t_SL _28858_ (.A1(_00574_),
    .A2(_06430_),
    .B(_06431_),
    .Y(_06432_));
 XNOR2x2_ASAP7_75t_SL _28859_ (.A(_00928_),
    .B(_06432_),
    .Y(_06433_));
 OAI21x1_ASAP7_75t_SL _28863_ (.A1(_06385_),
    .A2(_06378_),
    .B(_06390_),
    .Y(_06437_));
 OAI21x1_ASAP7_75t_SL _28864_ (.A1(_06389_),
    .A2(_06387_),
    .B(_00913_),
    .Y(_06438_));
 NAND2x2_ASAP7_75t_SL _28865_ (.A(_06438_),
    .B(_06437_),
    .Y(_06439_));
 NAND2x1_ASAP7_75t_SL _28867_ (.A(_06421_),
    .B(_06405_),
    .Y(_06440_));
 NOR2x1_ASAP7_75t_SL _28868_ (.A(_06439_),
    .B(_06440_),
    .Y(_06441_));
 XNOR2x2_ASAP7_75t_L _28869_ (.A(_03741_),
    .B(_03740_),
    .Y(_06442_));
 XOR2x2_ASAP7_75t_SL _28870_ (.A(_12148_),
    .B(_00658_),
    .Y(_06443_));
 AND2x2_ASAP7_75t_SL _28871_ (.A(_06442_),
    .B(_06443_),
    .Y(_06444_));
 OAI21x1_ASAP7_75t_R _28872_ (.A1(_06443_),
    .A2(_06442_),
    .B(_00574_),
    .Y(_06445_));
 NAND2x1_ASAP7_75t_R _28873_ (.A(_00534_),
    .B(_10675_),
    .Y(_06446_));
 OAI21x1_ASAP7_75t_SL _28874_ (.A1(_06444_),
    .A2(_06445_),
    .B(_06446_),
    .Y(_06447_));
 XNOR2x2_ASAP7_75t_SL _28875_ (.A(_00927_),
    .B(_06447_),
    .Y(_06448_));
 INVx2_ASAP7_75t_SL _28877_ (.A(_01365_),
    .Y(_06450_));
 AOI21x1_ASAP7_75t_SL _28878_ (.A1(_06426_),
    .A2(_06427_),
    .B(_06450_),
    .Y(_06451_));
 INVx2_ASAP7_75t_SL _28879_ (.A(_06451_),
    .Y(_06452_));
 NAND2x1p5_ASAP7_75t_SL _28880_ (.A(_06452_),
    .B(_06448_),
    .Y(_06453_));
 INVx1_ASAP7_75t_R _28881_ (.A(_01370_),
    .Y(_06454_));
 AO21x1_ASAP7_75t_SL _28882_ (.A1(_06427_),
    .A2(_06426_),
    .B(_06454_),
    .Y(_06455_));
 INVx2_ASAP7_75t_SL _28883_ (.A(_01364_),
    .Y(_06456_));
 AOI21x1_ASAP7_75t_SL _28884_ (.A1(_06415_),
    .A2(_06420_),
    .B(_06456_),
    .Y(_06457_));
 INVx1_ASAP7_75t_SL _28885_ (.A(_06457_),
    .Y(_06458_));
 AO21x1_ASAP7_75t_SL _28887_ (.A1(_06455_),
    .A2(_06458_),
    .B(_06448_),
    .Y(_06460_));
 OA21x2_ASAP7_75t_SL _28888_ (.A1(_06441_),
    .A2(_06453_),
    .B(_06460_),
    .Y(_06461_));
 NOR2x1_ASAP7_75t_R _28889_ (.A(_06405_),
    .B(_06392_),
    .Y(_06462_));
 OAI21x1_ASAP7_75t_SL _28892_ (.A1(_06421_),
    .A2(_06424_),
    .B(_06448_),
    .Y(_06465_));
 NOR2x1_ASAP7_75t_SL _28893_ (.A(_06462_),
    .B(_06465_),
    .Y(_06466_));
 NOR2x1_ASAP7_75t_SL _28894_ (.A(_06428_),
    .B(_06424_),
    .Y(_06467_));
 AO21x1_ASAP7_75t_SL _28895_ (.A1(_06392_),
    .A2(_06424_),
    .B(_06448_),
    .Y(_06468_));
 INVx2_ASAP7_75t_SL _28896_ (.A(_06433_),
    .Y(_06469_));
 OAI21x1_ASAP7_75t_SL _28898_ (.A1(_06467_),
    .A2(_06468_),
    .B(_06469_),
    .Y(_06471_));
 XOR2x1_ASAP7_75t_SL _28899_ (.A(_00595_),
    .Y(_06472_),
    .B(_00596_));
 XOR2x2_ASAP7_75t_R _28900_ (.A(_06472_),
    .B(_14965_),
    .Y(_06473_));
 XOR2x2_ASAP7_75t_SL _28901_ (.A(_06473_),
    .B(_12190_),
    .Y(_06474_));
 NOR2x1_ASAP7_75t_R _28902_ (.A(_00574_),
    .B(_00532_),
    .Y(_06475_));
 AO21x1_ASAP7_75t_R _28903_ (.A1(_06474_),
    .A2(_00574_),
    .B(_06475_),
    .Y(_06476_));
 NOR2x1_ASAP7_75t_R _28904_ (.A(_00929_),
    .B(_06476_),
    .Y(_06477_));
 AND2x2_ASAP7_75t_R _28905_ (.A(_06476_),
    .B(_00929_),
    .Y(_06478_));
 NOR2x2_ASAP7_75t_SL _28906_ (.A(_06477_),
    .B(_06478_),
    .Y(_06479_));
 INVx1_ASAP7_75t_SL _28907_ (.A(_06479_),
    .Y(_06480_));
 OAI21x1_ASAP7_75t_SL _28909_ (.A1(_06466_),
    .A2(_06471_),
    .B(_06480_),
    .Y(_06482_));
 AOI21x1_ASAP7_75t_SL _28910_ (.A1(_06433_),
    .A2(_06461_),
    .B(_06482_),
    .Y(_06483_));
 INVx1_ASAP7_75t_SL _28912_ (.A(_06415_),
    .Y(_06485_));
 NOR3x1_ASAP7_75t_R _28913_ (.A(_06414_),
    .B(_08790_),
    .C(_06406_),
    .Y(_06486_));
 OAI21x1_ASAP7_75t_R _28914_ (.A1(_06485_),
    .A2(_06486_),
    .B(_01370_),
    .Y(_06487_));
 INVx1_ASAP7_75t_SL _28915_ (.A(_06487_),
    .Y(_06488_));
 NOR2x1p5_ASAP7_75t_SL _28916_ (.A(_06451_),
    .B(_06448_),
    .Y(_06489_));
 AO21x1_ASAP7_75t_SL _28917_ (.A1(_06420_),
    .A2(_06415_),
    .B(_01364_),
    .Y(_06490_));
 AOI22x1_ASAP7_75t_SL _28918_ (.A1(_06448_),
    .A2(_06488_),
    .B1(_06489_),
    .B2(_06490_),
    .Y(_06491_));
 AOI21x1_ASAP7_75t_SL _28919_ (.A1(_06426_),
    .A2(_06427_),
    .B(_06456_),
    .Y(_06492_));
 AND2x2_ASAP7_75t_SL _28920_ (.A(_06492_),
    .B(_06448_),
    .Y(_06493_));
 NOR2x1_ASAP7_75t_SL _28921_ (.A(_06469_),
    .B(_06493_),
    .Y(_06494_));
 AND2x2_ASAP7_75t_SL _28922_ (.A(_06491_),
    .B(_06494_),
    .Y(_06495_));
 NOR2x2_ASAP7_75t_SL _28924_ (.A(_06428_),
    .B(_06392_),
    .Y(_06497_));
 AND2x4_ASAP7_75t_SL _28925_ (.A(_06448_),
    .B(_06451_),
    .Y(_06498_));
 AOI21x1_ASAP7_75t_SL _28926_ (.A1(_06415_),
    .A2(_06420_),
    .B(_06450_),
    .Y(_06499_));
 NOR2x1p5_ASAP7_75t_SL _28927_ (.A(_06499_),
    .B(_06448_),
    .Y(_06500_));
 AOI211x1_ASAP7_75t_SL _28928_ (.A1(_06448_),
    .A2(_06497_),
    .B(_06500_),
    .C(_06498_),
    .Y(_06501_));
 OAI21x1_ASAP7_75t_SL _28930_ (.A1(_06501_),
    .A2(_06433_),
    .B(_06479_),
    .Y(_06503_));
 XOR2x2_ASAP7_75t_SL _28931_ (.A(_00596_),
    .B(_00597_),
    .Y(_06504_));
 XOR2x2_ASAP7_75t_R _28932_ (.A(_06504_),
    .B(_15007_),
    .Y(_06505_));
 XOR2x2_ASAP7_75t_R _28933_ (.A(_06505_),
    .B(_12223_),
    .Y(_06506_));
 NOR2x1_ASAP7_75t_R _28934_ (.A(_00574_),
    .B(_00531_),
    .Y(_06507_));
 AO21x1_ASAP7_75t_SL _28935_ (.A1(_06506_),
    .A2(_00574_),
    .B(_06507_),
    .Y(_06508_));
 XOR2x2_ASAP7_75t_SL _28936_ (.A(_06508_),
    .B(_00930_),
    .Y(_06509_));
 OAI21x1_ASAP7_75t_SL _28938_ (.A1(_06503_),
    .A2(_06495_),
    .B(_06509_),
    .Y(_06511_));
 NOR2x1_ASAP7_75t_SL _28939_ (.A(_06511_),
    .B(_06483_),
    .Y(_06512_));
 XOR2x2_ASAP7_75t_SL _28940_ (.A(_06447_),
    .B(_00927_),
    .Y(_06513_));
 OAI21x1_ASAP7_75t_SL _28942_ (.A1(_06421_),
    .A2(_06450_),
    .B(_06513_),
    .Y(_06515_));
 INVx1_ASAP7_75t_SL _28944_ (.A(_01373_),
    .Y(_06517_));
 NOR2x1_ASAP7_75t_SL _28945_ (.A(_06517_),
    .B(_06428_),
    .Y(_06518_));
 OA21x2_ASAP7_75t_SL _28946_ (.A1(_06515_),
    .A2(_06518_),
    .B(_06469_),
    .Y(_06519_));
 NOR2x1_ASAP7_75t_SL _28947_ (.A(_06421_),
    .B(_06424_),
    .Y(_06520_));
 AOI21x1_ASAP7_75t_SL _28948_ (.A1(_06424_),
    .A2(_06392_),
    .B(_06428_),
    .Y(_06521_));
 OAI21x1_ASAP7_75t_SL _28950_ (.A1(_06520_),
    .A2(_06521_),
    .B(_06448_),
    .Y(_06523_));
 AND2x2_ASAP7_75t_SL _28951_ (.A(_06519_),
    .B(_06523_),
    .Y(_06524_));
 INVx1_ASAP7_75t_SL _28954_ (.A(_01368_),
    .Y(_06527_));
 OAI21x1_ASAP7_75t_SL _28956_ (.A1(_06527_),
    .A2(_06421_),
    .B(_06513_),
    .Y(_06529_));
 NAND2x1_ASAP7_75t_SL _28957_ (.A(_06421_),
    .B(_06424_),
    .Y(_06530_));
 NOR2x1_ASAP7_75t_SL _28958_ (.A(_06439_),
    .B(_06530_),
    .Y(_06531_));
 OAI21x1_ASAP7_75t_SL _28960_ (.A1(_06428_),
    .A2(_06405_),
    .B(_06448_),
    .Y(_06533_));
 OAI21x1_ASAP7_75t_SL _28961_ (.A1(_06529_),
    .A2(_06531_),
    .B(_06533_),
    .Y(_06534_));
 OAI21x1_ASAP7_75t_SL _28964_ (.A1(_06469_),
    .A2(_06534_),
    .B(_06480_),
    .Y(_06537_));
 INVx1_ASAP7_75t_SL _28965_ (.A(_06509_),
    .Y(_06538_));
 OAI21x1_ASAP7_75t_SL _28967_ (.A1(_06524_),
    .A2(_06537_),
    .B(_06538_),
    .Y(_06540_));
 AOI21x1_ASAP7_75t_SL _28969_ (.A1(_06426_),
    .A2(_06427_),
    .B(_01366_),
    .Y(_06542_));
 OAI21x1_ASAP7_75t_SL _28970_ (.A1(_06542_),
    .A2(_06497_),
    .B(_06448_),
    .Y(_06543_));
 AOI21x1_ASAP7_75t_SL _28971_ (.A1(_06421_),
    .A2(_06424_),
    .B(_06448_),
    .Y(_06544_));
 NAND2x1_ASAP7_75t_SL _28972_ (.A(_06392_),
    .B(_06520_),
    .Y(_06545_));
 AOI21x1_ASAP7_75t_SL _28974_ (.A1(_06544_),
    .A2(_06545_),
    .B(_06469_),
    .Y(_06547_));
 AO21x1_ASAP7_75t_SL _28976_ (.A1(_06439_),
    .A2(_06428_),
    .B(_06513_),
    .Y(_06549_));
 NOR2x1_ASAP7_75t_SL _28977_ (.A(_06549_),
    .B(_06531_),
    .Y(_06550_));
 AO21x1_ASAP7_75t_R _28978_ (.A1(_06427_),
    .A2(_06426_),
    .B(_06517_),
    .Y(_06551_));
 AO21x1_ASAP7_75t_SL _28980_ (.A1(_06544_),
    .A2(_06551_),
    .B(_06433_),
    .Y(_06553_));
 OAI21x1_ASAP7_75t_SL _28981_ (.A1(_06550_),
    .A2(_06553_),
    .B(_06479_),
    .Y(_06554_));
 AOI21x1_ASAP7_75t_SL _28982_ (.A1(_06543_),
    .A2(_06547_),
    .B(_06554_),
    .Y(_06555_));
 XOR2x2_ASAP7_75t_R _28983_ (.A(_00597_),
    .B(_00598_),
    .Y(_06556_));
 XOR2x2_ASAP7_75t_SL _28984_ (.A(_06556_),
    .B(_00693_),
    .Y(_06557_));
 XOR2x2_ASAP7_75t_SL _28985_ (.A(_06557_),
    .B(_12270_),
    .Y(_06558_));
 NOR2x1_ASAP7_75t_SL _28986_ (.A(_00574_),
    .B(_00530_),
    .Y(_06559_));
 AO21x1_ASAP7_75t_SL _28987_ (.A1(_06558_),
    .A2(_00574_),
    .B(_06559_),
    .Y(_06560_));
 XOR2x2_ASAP7_75t_SL _28988_ (.A(_06560_),
    .B(_00931_),
    .Y(_06561_));
 OAI21x1_ASAP7_75t_SL _28990_ (.A1(_06540_),
    .A2(_06555_),
    .B(_06561_),
    .Y(_06563_));
 OAI21x1_ASAP7_75t_SL _28992_ (.A1(_06405_),
    .A2(_06439_),
    .B(_06428_),
    .Y(_06565_));
 AOI21x1_ASAP7_75t_SL _28993_ (.A1(_06415_),
    .A2(_06420_),
    .B(_01368_),
    .Y(_06566_));
 NAND2x1p5_ASAP7_75t_SL _28994_ (.A(_06566_),
    .B(_06448_),
    .Y(_06567_));
 OAI21x1_ASAP7_75t_SL _28995_ (.A1(_06513_),
    .A2(_06565_),
    .B(_06567_),
    .Y(_06568_));
 AO21x1_ASAP7_75t_SL _28996_ (.A1(_06420_),
    .A2(_06415_),
    .B(_01366_),
    .Y(_06569_));
 INVx1_ASAP7_75t_SL _28997_ (.A(_06569_),
    .Y(_06570_));
 NAND2x1_ASAP7_75t_SL _28998_ (.A(_06448_),
    .B(_06570_),
    .Y(_06571_));
 AND3x1_ASAP7_75t_SL _28999_ (.A(_06405_),
    .B(_06421_),
    .C(_06513_),
    .Y(_06572_));
 AO21x1_ASAP7_75t_SL _29000_ (.A1(_06492_),
    .A2(_06513_),
    .B(_06469_),
    .Y(_06573_));
 NOR2x1_ASAP7_75t_SL _29001_ (.A(_06572_),
    .B(_06573_),
    .Y(_06574_));
 NAND2x1_ASAP7_75t_SL _29002_ (.A(_06571_),
    .B(_06574_),
    .Y(_06575_));
 INVx1_ASAP7_75t_SL _29004_ (.A(_01378_),
    .Y(_06577_));
 AOI21x1_ASAP7_75t_SL _29005_ (.A1(_06415_),
    .A2(_06420_),
    .B(_01365_),
    .Y(_06578_));
 NOR2x1p5_ASAP7_75t_SL _29006_ (.A(_06578_),
    .B(_06513_),
    .Y(_06579_));
 INVx2_ASAP7_75t_SL _29007_ (.A(_06579_),
    .Y(_06580_));
 OAI21x1_ASAP7_75t_SL _29008_ (.A1(_06577_),
    .A2(_06448_),
    .B(_06580_),
    .Y(_06581_));
 AOI21x1_ASAP7_75t_SL _29009_ (.A1(_06469_),
    .A2(_06581_),
    .B(_06480_),
    .Y(_06582_));
 OAI21x1_ASAP7_75t_SL _29010_ (.A1(_06568_),
    .A2(_06575_),
    .B(_06582_),
    .Y(_06583_));
 NOR2x1_ASAP7_75t_SL _29011_ (.A(_06421_),
    .B(_06439_),
    .Y(_06584_));
 NAND2x1_ASAP7_75t_SL _29012_ (.A(_06424_),
    .B(_06584_),
    .Y(_06585_));
 AOI21x1_ASAP7_75t_SL _29014_ (.A1(_06454_),
    .A2(_06421_),
    .B(_06513_),
    .Y(_06587_));
 AO21x1_ASAP7_75t_SL _29016_ (.A1(_06542_),
    .A2(_06513_),
    .B(_06433_),
    .Y(_06589_));
 AO21x1_ASAP7_75t_SL _29017_ (.A1(_06585_),
    .A2(_06587_),
    .B(_06589_),
    .Y(_06590_));
 AOI21x1_ASAP7_75t_SL _29019_ (.A1(_06448_),
    .A2(_06542_),
    .B(_06469_),
    .Y(_06592_));
 AOI21x1_ASAP7_75t_SL _29021_ (.A1(_01371_),
    .A2(_06421_),
    .B(_06448_),
    .Y(_06594_));
 NAND2x1_ASAP7_75t_SL _29022_ (.A(_06594_),
    .B(_06585_),
    .Y(_06595_));
 AOI21x1_ASAP7_75t_SL _29024_ (.A1(_06592_),
    .A2(_06595_),
    .B(_06479_),
    .Y(_06597_));
 AOI21x1_ASAP7_75t_SL _29025_ (.A1(_06590_),
    .A2(_06597_),
    .B(_06538_),
    .Y(_06598_));
 NAND2x1_ASAP7_75t_SL _29026_ (.A(_06598_),
    .B(_06583_),
    .Y(_06599_));
 OAI21x1_ASAP7_75t_SL _29027_ (.A1(_06542_),
    .A2(_06457_),
    .B(_06448_),
    .Y(_06600_));
 AOI21x1_ASAP7_75t_SL _29029_ (.A1(_01368_),
    .A2(_06428_),
    .B(_06448_),
    .Y(_06602_));
 NOR2x1_ASAP7_75t_SL _29030_ (.A(_06433_),
    .B(_06602_),
    .Y(_06603_));
 AOI21x1_ASAP7_75t_SL _29031_ (.A1(_06600_),
    .A2(_06603_),
    .B(_06479_),
    .Y(_06604_));
 INVx2_ASAP7_75t_SL _29032_ (.A(_06578_),
    .Y(_06605_));
 AOI21x1_ASAP7_75t_SL _29033_ (.A1(_06428_),
    .A2(_06392_),
    .B(_06513_),
    .Y(_06606_));
 AOI21x1_ASAP7_75t_SL _29034_ (.A1(_06605_),
    .A2(_06606_),
    .B(_06469_),
    .Y(_06607_));
 NAND2x1_ASAP7_75t_SL _29035_ (.A(_06428_),
    .B(_06405_),
    .Y(_06608_));
 AO21x1_ASAP7_75t_SL _29036_ (.A1(_06608_),
    .A2(_06487_),
    .B(_06448_),
    .Y(_06609_));
 NAND2x1_ASAP7_75t_SL _29037_ (.A(_06607_),
    .B(_06609_),
    .Y(_06610_));
 AOI21x1_ASAP7_75t_SL _29038_ (.A1(_06604_),
    .A2(_06610_),
    .B(_06509_),
    .Y(_06611_));
 AOI21x1_ASAP7_75t_SL _29039_ (.A1(_06426_),
    .A2(_06427_),
    .B(_01371_),
    .Y(_06612_));
 NOR2x1p5_ASAP7_75t_SL _29040_ (.A(_06566_),
    .B(_06612_),
    .Y(_06613_));
 NOR2x1_ASAP7_75t_SL _29041_ (.A(_06513_),
    .B(_06613_),
    .Y(_06614_));
 NAND2x1_ASAP7_75t_SL _29042_ (.A(_06469_),
    .B(_06515_),
    .Y(_06615_));
 OA21x2_ASAP7_75t_SL _29044_ (.A1(_06614_),
    .A2(_06615_),
    .B(_06479_),
    .Y(_06617_));
 NAND2x1_ASAP7_75t_SL _29045_ (.A(_06567_),
    .B(_06547_),
    .Y(_06618_));
 NAND2x1_ASAP7_75t_SL _29046_ (.A(_06617_),
    .B(_06618_),
    .Y(_06619_));
 AOI21x1_ASAP7_75t_SL _29047_ (.A1(_06611_),
    .A2(_06619_),
    .B(_06561_),
    .Y(_06620_));
 NAND2x1_ASAP7_75t_SL _29048_ (.A(_06599_),
    .B(_06620_),
    .Y(_06621_));
 OAI21x1_ASAP7_75t_SL _29049_ (.A1(_06512_),
    .A2(_06563_),
    .B(_06621_),
    .Y(_00144_));
 AOI21x1_ASAP7_75t_SL _29050_ (.A1(_06405_),
    .A2(_06392_),
    .B(_06421_),
    .Y(_06622_));
 NOR2x1_ASAP7_75t_SL _29051_ (.A(_06622_),
    .B(_06521_),
    .Y(_06623_));
 NAND2x1_ASAP7_75t_SL _29052_ (.A(_06428_),
    .B(_06424_),
    .Y(_06624_));
 AOI21x1_ASAP7_75t_R _29053_ (.A1(_06456_),
    .A2(_06421_),
    .B(_06513_),
    .Y(_06625_));
 AOI21x1_ASAP7_75t_R _29054_ (.A1(_06624_),
    .A2(_06625_),
    .B(_06479_),
    .Y(_06626_));
 OAI21x1_ASAP7_75t_R _29055_ (.A1(_06448_),
    .A2(_06623_),
    .B(_06626_),
    .Y(_06627_));
 AOI21x1_ASAP7_75t_R _29056_ (.A1(_06428_),
    .A2(_06405_),
    .B(_06513_),
    .Y(_06628_));
 NOR2x1_ASAP7_75t_SL _29057_ (.A(_06428_),
    .B(_06439_),
    .Y(_06629_));
 INVx1_ASAP7_75t_SL _29058_ (.A(_06629_),
    .Y(_06630_));
 NAND2x1_ASAP7_75t_SL _29059_ (.A(_06628_),
    .B(_06630_),
    .Y(_06631_));
 NAND2x1_ASAP7_75t_SL _29060_ (.A(_06421_),
    .B(_06439_),
    .Y(_06632_));
 NAND2x1_ASAP7_75t_SL _29061_ (.A(_06632_),
    .B(_06602_),
    .Y(_06633_));
 NAND3x1_ASAP7_75t_SL _29062_ (.A(_06631_),
    .B(_06633_),
    .C(_06479_),
    .Y(_06634_));
 NAND2x1_ASAP7_75t_SL _29063_ (.A(_06627_),
    .B(_06634_),
    .Y(_06635_));
 NAND2x1_ASAP7_75t_SL _29064_ (.A(_06405_),
    .B(_06392_),
    .Y(_06636_));
 OAI21x1_ASAP7_75t_SL _29065_ (.A1(_06421_),
    .A2(_06636_),
    .B(_06587_),
    .Y(_06637_));
 INVx1_ASAP7_75t_R _29066_ (.A(_01380_),
    .Y(_06638_));
 NOR2x1_ASAP7_75t_R _29067_ (.A(_06638_),
    .B(_06448_),
    .Y(_06639_));
 AOI21x1_ASAP7_75t_R _29068_ (.A1(_06639_),
    .A2(_06479_),
    .B(_06469_),
    .Y(_06640_));
 AO21x1_ASAP7_75t_R _29069_ (.A1(_06637_),
    .A2(_06640_),
    .B(_06538_),
    .Y(_06641_));
 AOI21x1_ASAP7_75t_R _29070_ (.A1(_06469_),
    .A2(_06635_),
    .B(_06641_),
    .Y(_06642_));
 NAND2x1_ASAP7_75t_R _29071_ (.A(_01366_),
    .B(_06421_),
    .Y(_06643_));
 AOI21x1_ASAP7_75t_R _29072_ (.A1(_01373_),
    .A2(_06428_),
    .B(_06513_),
    .Y(_06644_));
 AOI21x1_ASAP7_75t_R _29073_ (.A1(_06643_),
    .A2(_06644_),
    .B(_06433_),
    .Y(_06645_));
 AOI21x1_ASAP7_75t_SL _29074_ (.A1(_06405_),
    .A2(_06392_),
    .B(_06428_),
    .Y(_06646_));
 OAI21x1_ASAP7_75t_SL _29076_ (.A1(_06451_),
    .A2(_06646_),
    .B(_06513_),
    .Y(_06648_));
 NAND2x1_ASAP7_75t_SL _29077_ (.A(_06645_),
    .B(_06648_),
    .Y(_06649_));
 NOR2x1_ASAP7_75t_L _29078_ (.A(_06469_),
    .B(_06489_),
    .Y(_06650_));
 AOI21x1_ASAP7_75t_SL _29079_ (.A1(_06421_),
    .A2(_06424_),
    .B(_06513_),
    .Y(_06651_));
 OAI21x1_ASAP7_75t_R _29080_ (.A1(_06421_),
    .A2(_06636_),
    .B(_06651_),
    .Y(_06652_));
 AOI21x1_ASAP7_75t_SL _29081_ (.A1(_06652_),
    .A2(_06650_),
    .B(_06480_),
    .Y(_06653_));
 NAND2x1_ASAP7_75t_L _29082_ (.A(_06649_),
    .B(_06653_),
    .Y(_06654_));
 NAND2x1_ASAP7_75t_R _29083_ (.A(_06490_),
    .B(_06628_),
    .Y(_06655_));
 AOI21x1_ASAP7_75t_R _29084_ (.A1(_06633_),
    .A2(_06655_),
    .B(_06469_),
    .Y(_06656_));
 OAI21x1_ASAP7_75t_R _29086_ (.A1(_06492_),
    .A2(_06578_),
    .B(_06513_),
    .Y(_06658_));
 OAI21x1_ASAP7_75t_R _29087_ (.A1(_06542_),
    .A2(_06467_),
    .B(_06448_),
    .Y(_06659_));
 AOI21x1_ASAP7_75t_R _29088_ (.A1(_06658_),
    .A2(_06659_),
    .B(_06433_),
    .Y(_06660_));
 OAI21x1_ASAP7_75t_R _29089_ (.A1(_06656_),
    .A2(_06660_),
    .B(_06480_),
    .Y(_06661_));
 AOI21x1_ASAP7_75t_R _29090_ (.A1(_06654_),
    .A2(_06661_),
    .B(_06509_),
    .Y(_06662_));
 OAI21x1_ASAP7_75t_SL _29091_ (.A1(_06642_),
    .A2(_06662_),
    .B(_06561_),
    .Y(_06663_));
 NOR2x1_ASAP7_75t_R _29092_ (.A(_06566_),
    .B(_06515_),
    .Y(_06664_));
 AOI211x1_ASAP7_75t_R _29094_ (.A1(_06405_),
    .A2(_06421_),
    .B(_06513_),
    .C(_06492_),
    .Y(_06666_));
 OAI21x1_ASAP7_75t_R _29095_ (.A1(_06664_),
    .A2(_06666_),
    .B(_06469_),
    .Y(_06667_));
 NOR2x1_ASAP7_75t_SL _29096_ (.A(_06421_),
    .B(_06405_),
    .Y(_06668_));
 NOR2x1_ASAP7_75t_SL _29097_ (.A(_06424_),
    .B(_06439_),
    .Y(_06669_));
 OAI21x1_ASAP7_75t_R _29098_ (.A1(_06668_),
    .A2(_06669_),
    .B(_06513_),
    .Y(_06670_));
 AOI21x1_ASAP7_75t_SL _29099_ (.A1(_06624_),
    .A2(_06579_),
    .B(_06469_),
    .Y(_06671_));
 AOI21x1_ASAP7_75t_R _29100_ (.A1(_06670_),
    .A2(_06671_),
    .B(_06480_),
    .Y(_06672_));
 NAND2x1_ASAP7_75t_SL _29101_ (.A(_06667_),
    .B(_06672_),
    .Y(_06673_));
 NAND2x1_ASAP7_75t_L _29102_ (.A(_06448_),
    .B(_06622_),
    .Y(_06674_));
 NAND2x1_ASAP7_75t_SL _29103_ (.A(_06428_),
    .B(_06439_),
    .Y(_06675_));
 AOI21x1_ASAP7_75t_SL _29104_ (.A1(_01373_),
    .A2(_06421_),
    .B(_06448_),
    .Y(_06676_));
 AOI21x1_ASAP7_75t_SL _29105_ (.A1(_06675_),
    .A2(_06676_),
    .B(_06433_),
    .Y(_06677_));
 NAND2x1_ASAP7_75t_R _29106_ (.A(_06674_),
    .B(_06677_),
    .Y(_06678_));
 AO21x1_ASAP7_75t_R _29107_ (.A1(_06427_),
    .A2(_06426_),
    .B(_01368_),
    .Y(_06679_));
 OA21x2_ASAP7_75t_R _29108_ (.A1(_06679_),
    .A2(_06513_),
    .B(_06433_),
    .Y(_06680_));
 AOI21x1_ASAP7_75t_R _29109_ (.A1(_06680_),
    .A2(_06648_),
    .B(_06479_),
    .Y(_06681_));
 NAND2x1_ASAP7_75t_R _29110_ (.A(_06678_),
    .B(_06681_),
    .Y(_06682_));
 AOI21x1_ASAP7_75t_R _29111_ (.A1(_06673_),
    .A2(_06682_),
    .B(_06509_),
    .Y(_06683_));
 AOI21x1_ASAP7_75t_R _29112_ (.A1(_06544_),
    .A2(_06452_),
    .B(_06433_),
    .Y(_06684_));
 AO21x1_ASAP7_75t_R _29113_ (.A1(_06530_),
    .A2(_06679_),
    .B(_06513_),
    .Y(_06685_));
 NAND2x1_ASAP7_75t_L _29114_ (.A(_06685_),
    .B(_06684_),
    .Y(_06686_));
 NOR2x2_ASAP7_75t_SL _29115_ (.A(_06448_),
    .B(_06428_),
    .Y(_06687_));
 NAND2x1_ASAP7_75t_SL _29116_ (.A(_06424_),
    .B(_06392_),
    .Y(_06688_));
 NAND2x1_ASAP7_75t_SL _29117_ (.A(_06687_),
    .B(_06688_),
    .Y(_06689_));
 NAND2x1_ASAP7_75t_SL _29118_ (.A(_06424_),
    .B(_06439_),
    .Y(_06690_));
 AOI21x1_ASAP7_75t_R _29119_ (.A1(_06690_),
    .A2(_06606_),
    .B(_06469_),
    .Y(_06691_));
 AOI21x1_ASAP7_75t_R _29120_ (.A1(_06689_),
    .A2(_06691_),
    .B(_06479_),
    .Y(_06692_));
 NAND2x1_ASAP7_75t_SL _29121_ (.A(_06686_),
    .B(_06692_),
    .Y(_06693_));
 INVx1_ASAP7_75t_SL _29122_ (.A(_06675_),
    .Y(_06694_));
 AOI21x1_ASAP7_75t_SL _29123_ (.A1(_06421_),
    .A2(_06392_),
    .B(_06448_),
    .Y(_06695_));
 NOR2x1_ASAP7_75t_SL _29124_ (.A(_06694_),
    .B(_06695_),
    .Y(_06696_));
 NAND3x1_ASAP7_75t_R _29126_ (.A(_06696_),
    .B(_06469_),
    .C(_06567_),
    .Y(_06698_));
 AOI21x1_ASAP7_75t_SL _29127_ (.A1(_06500_),
    .A2(_06551_),
    .B(_06469_),
    .Y(_06699_));
 AOI21x1_ASAP7_75t_R _29128_ (.A1(_06424_),
    .A2(_06392_),
    .B(_06421_),
    .Y(_06700_));
 OAI21x1_ASAP7_75t_R _29129_ (.A1(_06566_),
    .A2(_06700_),
    .B(_06448_),
    .Y(_06701_));
 AOI21x1_ASAP7_75t_SL _29130_ (.A1(_06701_),
    .A2(_06699_),
    .B(_06480_),
    .Y(_06702_));
 NAND2x1_ASAP7_75t_SL _29131_ (.A(_06702_),
    .B(_06698_),
    .Y(_06703_));
 AOI21x1_ASAP7_75t_SL _29132_ (.A1(_06703_),
    .A2(_06693_),
    .B(_06538_),
    .Y(_06704_));
 INVx1_ASAP7_75t_SL _29133_ (.A(_06561_),
    .Y(_06705_));
 OAI21x1_ASAP7_75t_SL _29134_ (.A1(_06704_),
    .A2(_06683_),
    .B(_06705_),
    .Y(_06706_));
 NAND2x1_ASAP7_75t_SL _29135_ (.A(_06706_),
    .B(_06663_),
    .Y(_00145_));
 OAI21x1_ASAP7_75t_SL _29136_ (.A1(_06428_),
    .A2(_06392_),
    .B(_06513_),
    .Y(_06707_));
 NOR2x1_ASAP7_75t_R _29137_ (.A(_06612_),
    .B(_06707_),
    .Y(_06708_));
 NOR2x1_ASAP7_75t_SL _29138_ (.A(_01373_),
    .B(_06428_),
    .Y(_06709_));
 OAI21x1_ASAP7_75t_SL _29139_ (.A1(_06709_),
    .A2(_06465_),
    .B(_06469_),
    .Y(_06710_));
 NOR2x1_ASAP7_75t_SL _29140_ (.A(_06708_),
    .B(_06710_),
    .Y(_06711_));
 AOI21x1_ASAP7_75t_SL _29141_ (.A1(_01371_),
    .A2(_06421_),
    .B(_06513_),
    .Y(_06712_));
 NAND2x1_ASAP7_75t_SL _29142_ (.A(_06624_),
    .B(_06712_),
    .Y(_06713_));
 NAND2x1_ASAP7_75t_L _29143_ (.A(_06605_),
    .B(_06489_),
    .Y(_06714_));
 AOI21x1_ASAP7_75t_R _29144_ (.A1(_06713_),
    .A2(_06714_),
    .B(_06469_),
    .Y(_06715_));
 OA21x2_ASAP7_75t_SL _29145_ (.A1(_06711_),
    .A2(_06715_),
    .B(_06480_),
    .Y(_06716_));
 INVx1_ASAP7_75t_L _29146_ (.A(_06612_),
    .Y(_06717_));
 AO21x1_ASAP7_75t_R _29147_ (.A1(_06420_),
    .A2(_06415_),
    .B(_01373_),
    .Y(_06718_));
 AOI21x1_ASAP7_75t_R _29148_ (.A1(_06717_),
    .A2(_06718_),
    .B(_06513_),
    .Y(_06719_));
 INVx2_ASAP7_75t_SL _29149_ (.A(_06566_),
    .Y(_06720_));
 AOI21x1_ASAP7_75t_R _29150_ (.A1(_06720_),
    .A2(_06608_),
    .B(_06448_),
    .Y(_06721_));
 OAI21x1_ASAP7_75t_R _29151_ (.A1(_06719_),
    .A2(_06721_),
    .B(_06469_),
    .Y(_06722_));
 NAND2x1_ASAP7_75t_SL _29152_ (.A(_06428_),
    .B(_06392_),
    .Y(_06723_));
 AOI21x1_ASAP7_75t_R _29153_ (.A1(_06720_),
    .A2(_06723_),
    .B(_06448_),
    .Y(_06724_));
 OAI21x1_ASAP7_75t_R _29154_ (.A1(_06614_),
    .A2(_06724_),
    .B(_06433_),
    .Y(_06725_));
 AOI21x1_ASAP7_75t_R _29155_ (.A1(_06722_),
    .A2(_06725_),
    .B(_06480_),
    .Y(_06726_));
 NOR3x1_ASAP7_75t_L _29156_ (.A(_06716_),
    .B(_06509_),
    .C(_06726_),
    .Y(_06727_));
 OAI21x1_ASAP7_75t_R _29157_ (.A1(_06527_),
    .A2(_06421_),
    .B(_06448_),
    .Y(_06728_));
 NOR2x1_ASAP7_75t_SL _29158_ (.A(_06518_),
    .B(_06728_),
    .Y(_06729_));
 OAI21x1_ASAP7_75t_SL _29159_ (.A1(_06694_),
    .A2(_06521_),
    .B(_06513_),
    .Y(_06730_));
 INVx1_ASAP7_75t_SL _29160_ (.A(_06730_),
    .Y(_06731_));
 OAI21x1_ASAP7_75t_R _29161_ (.A1(_06729_),
    .A2(_06731_),
    .B(_06469_),
    .Y(_06732_));
 NAND2x1p5_ASAP7_75t_L _29162_ (.A(_06606_),
    .B(_06605_),
    .Y(_06733_));
 OAI21x1_ASAP7_75t_R _29163_ (.A1(_06421_),
    .A2(_06424_),
    .B(_06513_),
    .Y(_06734_));
 NOR2x1_ASAP7_75t_SL _29164_ (.A(_06566_),
    .B(_06734_),
    .Y(_06735_));
 AOI21x1_ASAP7_75t_SL _29165_ (.A1(_06675_),
    .A2(_06735_),
    .B(_06469_),
    .Y(_06736_));
 NAND2x1_ASAP7_75t_L _29166_ (.A(_06733_),
    .B(_06736_),
    .Y(_06737_));
 AOI21x1_ASAP7_75t_R _29167_ (.A1(_06732_),
    .A2(_06737_),
    .B(_06480_),
    .Y(_06738_));
 AOI21x1_ASAP7_75t_SL _29168_ (.A1(_06426_),
    .A2(_06427_),
    .B(_01365_),
    .Y(_06739_));
 OAI21x1_ASAP7_75t_R _29169_ (.A1(_06428_),
    .A2(_06392_),
    .B(_06448_),
    .Y(_06740_));
 NOR2x1_ASAP7_75t_L _29170_ (.A(_06740_),
    .B(_06739_),
    .Y(_06741_));
 NOR2x1_ASAP7_75t_R _29171_ (.A(_06570_),
    .B(_06734_),
    .Y(_06742_));
 OA21x2_ASAP7_75t_R _29172_ (.A1(_06741_),
    .A2(_06742_),
    .B(_06469_),
    .Y(_06743_));
 OAI21x1_ASAP7_75t_SL _29173_ (.A1(_06439_),
    .A2(_06530_),
    .B(_06448_),
    .Y(_06744_));
 NAND2x1_ASAP7_75t_R _29174_ (.A(_06433_),
    .B(_06744_),
    .Y(_06745_));
 NOR2x1_ASAP7_75t_SL _29175_ (.A(_01373_),
    .B(_06421_),
    .Y(_06746_));
 OA21x2_ASAP7_75t_R _29176_ (.A1(_06646_),
    .A2(_06746_),
    .B(_06513_),
    .Y(_06747_));
 OAI21x1_ASAP7_75t_R _29177_ (.A1(_06745_),
    .A2(_06747_),
    .B(_06480_),
    .Y(_06748_));
 OAI21x1_ASAP7_75t_R _29178_ (.A1(_06743_),
    .A2(_06748_),
    .B(_06509_),
    .Y(_06749_));
 OAI21x1_ASAP7_75t_R _29179_ (.A1(_06738_),
    .A2(_06749_),
    .B(_06561_),
    .Y(_06750_));
 NAND2x1_ASAP7_75t_SL _29180_ (.A(_01377_),
    .B(_06513_),
    .Y(_06751_));
 AOI21x1_ASAP7_75t_R _29181_ (.A1(_06751_),
    .A2(_06744_),
    .B(_06469_),
    .Y(_06752_));
 OR2x2_ASAP7_75t_R _29182_ (.A(_06513_),
    .B(_01382_),
    .Y(_06753_));
 AOI21x1_ASAP7_75t_R _29183_ (.A1(_06753_),
    .A2(_06730_),
    .B(_06433_),
    .Y(_06754_));
 OAI21x1_ASAP7_75t_SL _29184_ (.A1(_06752_),
    .A2(_06754_),
    .B(_06479_),
    .Y(_06755_));
 INVx2_ASAP7_75t_SL _29185_ (.A(_06739_),
    .Y(_06756_));
 AO21x1_ASAP7_75t_SL _29186_ (.A1(_06720_),
    .A2(_06756_),
    .B(_06448_),
    .Y(_06757_));
 AOI21x1_ASAP7_75t_SL _29187_ (.A1(_06494_),
    .A2(_06757_),
    .B(_06479_),
    .Y(_06758_));
 AOI22x1_ASAP7_75t_R _29188_ (.A1(_01366_),
    .A2(_01368_),
    .B1(_06427_),
    .B2(_06426_),
    .Y(_06759_));
 OAI21x1_ASAP7_75t_R _29189_ (.A1(_06759_),
    .A2(_06646_),
    .B(_06513_),
    .Y(_06760_));
 AOI21x1_ASAP7_75t_R _29190_ (.A1(_06587_),
    .A2(_06545_),
    .B(_06433_),
    .Y(_06761_));
 NAND2x1_ASAP7_75t_SL _29191_ (.A(_06760_),
    .B(_06761_),
    .Y(_06762_));
 AOI21x1_ASAP7_75t_SL _29192_ (.A1(_06758_),
    .A2(_06762_),
    .B(_06538_),
    .Y(_06763_));
 NAND2x1_ASAP7_75t_SL _29193_ (.A(_06763_),
    .B(_06755_),
    .Y(_06764_));
 NAND2x1_ASAP7_75t_R _29194_ (.A(_06513_),
    .B(_06455_),
    .Y(_06765_));
 NOR2x1_ASAP7_75t_R _29195_ (.A(_06578_),
    .B(_06765_),
    .Y(_06766_));
 AND2x2_ASAP7_75t_SL _29196_ (.A(_06606_),
    .B(_06458_),
    .Y(_06767_));
 OAI21x1_ASAP7_75t_R _29197_ (.A1(_06766_),
    .A2(_06767_),
    .B(_06469_),
    .Y(_06768_));
 AOI21x1_ASAP7_75t_R _29198_ (.A1(_06424_),
    .A2(_06439_),
    .B(_06448_),
    .Y(_06769_));
 NOR2x1_ASAP7_75t_R _29199_ (.A(_06638_),
    .B(_06513_),
    .Y(_06770_));
 AOI21x1_ASAP7_75t_R _29200_ (.A1(_06723_),
    .A2(_06769_),
    .B(_06770_),
    .Y(_06771_));
 AOI21x1_ASAP7_75t_R _29201_ (.A1(_06433_),
    .A2(_06771_),
    .B(_06480_),
    .Y(_06772_));
 NAND2x1_ASAP7_75t_SL _29202_ (.A(_06768_),
    .B(_06772_),
    .Y(_06773_));
 AOI21x1_ASAP7_75t_R _29203_ (.A1(_06421_),
    .A2(_06439_),
    .B(_06448_),
    .Y(_06774_));
 NAND2x1_ASAP7_75t_SL _29204_ (.A(_06624_),
    .B(_06774_),
    .Y(_06775_));
 AOI21x1_ASAP7_75t_SL _29205_ (.A1(_06605_),
    .A2(_06606_),
    .B(_06433_),
    .Y(_06776_));
 NAND2x1_ASAP7_75t_SL _29206_ (.A(_06775_),
    .B(_06776_),
    .Y(_06777_));
 OA21x2_ASAP7_75t_R _29207_ (.A1(_01378_),
    .A2(_06513_),
    .B(_06433_),
    .Y(_06778_));
 OAI21x1_ASAP7_75t_SL _29208_ (.A1(_06421_),
    .A2(_06688_),
    .B(_06500_),
    .Y(_06779_));
 AOI21x1_ASAP7_75t_SL _29209_ (.A1(_06779_),
    .A2(_06778_),
    .B(_06479_),
    .Y(_06780_));
 AOI21x1_ASAP7_75t_SL _29210_ (.A1(_06780_),
    .A2(_06777_),
    .B(_06509_),
    .Y(_06781_));
 AOI21x1_ASAP7_75t_SL _29211_ (.A1(_06781_),
    .A2(_06773_),
    .B(_06561_),
    .Y(_06782_));
 NAND2x1_ASAP7_75t_SL _29212_ (.A(_06782_),
    .B(_06764_),
    .Y(_06783_));
 OAI21x1_ASAP7_75t_SL _29213_ (.A1(_06727_),
    .A2(_06750_),
    .B(_06783_),
    .Y(_00146_));
 OAI21x1_ASAP7_75t_SL _29214_ (.A1(_06709_),
    .A2(_06759_),
    .B(_06513_),
    .Y(_06784_));
 AOI21x1_ASAP7_75t_SL _29215_ (.A1(_06452_),
    .A2(_06651_),
    .B(_06480_),
    .Y(_06785_));
 NAND2x1_ASAP7_75t_SL _29216_ (.A(_06784_),
    .B(_06785_),
    .Y(_06786_));
 AND2x2_ASAP7_75t_L _29217_ (.A(_06612_),
    .B(_06513_),
    .Y(_06787_));
 NOR2x1_ASAP7_75t_SL _29218_ (.A(_06479_),
    .B(_06787_),
    .Y(_06788_));
 AOI21x1_ASAP7_75t_SL _29219_ (.A1(_06713_),
    .A2(_06788_),
    .B(_06469_),
    .Y(_06789_));
 NAND2x1_ASAP7_75t_SL _29220_ (.A(_06786_),
    .B(_06789_),
    .Y(_06790_));
 AND2x2_ASAP7_75t_SL _29221_ (.A(_06542_),
    .B(_06513_),
    .Y(_06791_));
 AO21x1_ASAP7_75t_SL _29222_ (.A1(_06498_),
    .A2(_06480_),
    .B(_06791_),
    .Y(_06792_));
 NAND2x1p5_ASAP7_75t_SL _29223_ (.A(_06499_),
    .B(_06513_),
    .Y(_06793_));
 NAND2x1_ASAP7_75t_SL _29224_ (.A(_06723_),
    .B(_06587_),
    .Y(_06794_));
 AOI21x1_ASAP7_75t_SL _29225_ (.A1(_06793_),
    .A2(_06794_),
    .B(_06480_),
    .Y(_06795_));
 OAI21x1_ASAP7_75t_SL _29226_ (.A1(_06792_),
    .A2(_06795_),
    .B(_06469_),
    .Y(_06796_));
 AOI21x1_ASAP7_75t_SL _29227_ (.A1(_06790_),
    .A2(_06796_),
    .B(_06538_),
    .Y(_06797_));
 NAND2x1_ASAP7_75t_SL _29228_ (.A(_06479_),
    .B(_06710_),
    .Y(_06798_));
 NOR2x1_ASAP7_75t_SL _29229_ (.A(_01371_),
    .B(_06428_),
    .Y(_06799_));
 OAI21x1_ASAP7_75t_SL _29230_ (.A1(_06799_),
    .A2(_06759_),
    .B(_06513_),
    .Y(_06800_));
 AOI21x1_ASAP7_75t_SL _29231_ (.A1(_06800_),
    .A2(_06637_),
    .B(_06469_),
    .Y(_06801_));
 OAI21x1_ASAP7_75t_SL _29232_ (.A1(_06798_),
    .A2(_06801_),
    .B(_06538_),
    .Y(_06802_));
 OAI21x1_ASAP7_75t_SL _29233_ (.A1(_06739_),
    .A2(_06709_),
    .B(_06448_),
    .Y(_06803_));
 NAND2x1_ASAP7_75t_SL _29234_ (.A(_06424_),
    .B(_06687_),
    .Y(_06804_));
 AOI21x1_ASAP7_75t_SL _29235_ (.A1(_06513_),
    .A2(_06612_),
    .B(_06433_),
    .Y(_06805_));
 NAND3x1_ASAP7_75t_SL _29236_ (.A(_06803_),
    .B(_06804_),
    .C(_06805_),
    .Y(_06806_));
 NAND2x1_ASAP7_75t_SL _29237_ (.A(_06690_),
    .B(_06606_),
    .Y(_06807_));
 NAND2x1_ASAP7_75t_SL _29238_ (.A(_06807_),
    .B(_06574_),
    .Y(_06808_));
 AOI21x1_ASAP7_75t_SL _29239_ (.A1(_06806_),
    .A2(_06808_),
    .B(_06479_),
    .Y(_06809_));
 NOR2x1_ASAP7_75t_SL _29240_ (.A(_06802_),
    .B(_06809_),
    .Y(_06810_));
 OAI21x1_ASAP7_75t_SL _29241_ (.A1(_06797_),
    .A2(_06810_),
    .B(_06561_),
    .Y(_06811_));
 OAI21x1_ASAP7_75t_SL _29242_ (.A1(_06629_),
    .A2(_06465_),
    .B(_06793_),
    .Y(_06812_));
 AOI21x1_ASAP7_75t_SL _29243_ (.A1(_06469_),
    .A2(_06812_),
    .B(_06480_),
    .Y(_06813_));
 NAND2x1_ASAP7_75t_SL _29244_ (.A(_06608_),
    .B(_06688_),
    .Y(_06814_));
 OA21x2_ASAP7_75t_SL _29245_ (.A1(_06515_),
    .A2(_06497_),
    .B(_06433_),
    .Y(_06815_));
 OAI21x1_ASAP7_75t_SL _29246_ (.A1(_06513_),
    .A2(_06814_),
    .B(_06815_),
    .Y(_06816_));
 AOI21x1_ASAP7_75t_SL _29247_ (.A1(_06816_),
    .A2(_06813_),
    .B(_06538_),
    .Y(_06817_));
 INVx2_ASAP7_75t_SL _29248_ (.A(_06492_),
    .Y(_06818_));
 AND2x2_ASAP7_75t_SL _29249_ (.A(_06500_),
    .B(_06818_),
    .Y(_06819_));
 AND3x1_ASAP7_75t_SL _29250_ (.A(_06440_),
    .B(_06448_),
    .C(_06455_),
    .Y(_06820_));
 OAI21x1_ASAP7_75t_SL _29251_ (.A1(_06819_),
    .A2(_06820_),
    .B(_06469_),
    .Y(_06821_));
 NOR2x1p5_ASAP7_75t_SL _29252_ (.A(_06739_),
    .B(_06513_),
    .Y(_06822_));
 AO21x1_ASAP7_75t_SL _29253_ (.A1(_06632_),
    .A2(_06822_),
    .B(_06469_),
    .Y(_06823_));
 OA21x2_ASAP7_75t_SL _29254_ (.A1(_06746_),
    .A2(_06566_),
    .B(_06513_),
    .Y(_06824_));
 OA21x2_ASAP7_75t_SL _29255_ (.A1(_06824_),
    .A2(_06823_),
    .B(_06480_),
    .Y(_06825_));
 NAND2x1p5_ASAP7_75t_SL _29256_ (.A(_06825_),
    .B(_06821_),
    .Y(_06826_));
 NAND2x1p5_ASAP7_75t_SL _29257_ (.A(_06826_),
    .B(_06817_),
    .Y(_06827_));
 NOR2x1_ASAP7_75t_SL _29258_ (.A(_06448_),
    .B(_06421_),
    .Y(_06828_));
 NOR2x1_ASAP7_75t_SL _29259_ (.A(_06469_),
    .B(_06828_),
    .Y(_06829_));
 NAND2x1_ASAP7_75t_SL _29260_ (.A(_06829_),
    .B(_06814_),
    .Y(_06830_));
 OAI21x1_ASAP7_75t_SL _29261_ (.A1(_06485_),
    .A2(_06486_),
    .B(_01371_),
    .Y(_06831_));
 NAND2x1p5_ASAP7_75t_SL _29262_ (.A(_06822_),
    .B(_06831_),
    .Y(_06832_));
 AOI21x1_ASAP7_75t_SL _29263_ (.A1(_06677_),
    .A2(_06832_),
    .B(_06480_),
    .Y(_06833_));
 AOI21x1_ASAP7_75t_SL _29264_ (.A1(_06833_),
    .A2(_06830_),
    .B(_06509_),
    .Y(_06834_));
 NOR2x1_ASAP7_75t_SL _29265_ (.A(_06622_),
    .B(_06580_),
    .Y(_06835_));
 OAI21x1_ASAP7_75t_SL _29266_ (.A1(_06521_),
    .A2(_06765_),
    .B(_06433_),
    .Y(_06836_));
 NOR2x1_ASAP7_75t_SL _29267_ (.A(_06835_),
    .B(_06836_),
    .Y(_06837_));
 NOR2x1_ASAP7_75t_SL _29268_ (.A(_06488_),
    .B(_06453_),
    .Y(_06838_));
 NOR2x1_ASAP7_75t_SL _29269_ (.A(_06838_),
    .B(_06471_),
    .Y(_06839_));
 OAI21x1_ASAP7_75t_SL _29270_ (.A1(_06837_),
    .A2(_06839_),
    .B(_06480_),
    .Y(_06840_));
 AOI21x1_ASAP7_75t_SL _29271_ (.A1(_06840_),
    .A2(_06834_),
    .B(_06561_),
    .Y(_06841_));
 NAND2x1_ASAP7_75t_SL _29272_ (.A(_06841_),
    .B(_06827_),
    .Y(_06842_));
 NAND2x1_ASAP7_75t_SL _29273_ (.A(_06842_),
    .B(_06811_),
    .Y(_00147_));
 NAND2x1_ASAP7_75t_R _29274_ (.A(_06392_),
    .B(_06687_),
    .Y(_06843_));
 AOI21x1_ASAP7_75t_R _29275_ (.A1(_06513_),
    .A2(_06492_),
    .B(_06469_),
    .Y(_06844_));
 NAND2x1_ASAP7_75t_R _29276_ (.A(_06843_),
    .B(_06844_),
    .Y(_06845_));
 OAI21x1_ASAP7_75t_R _29277_ (.A1(_06845_),
    .A2(_06568_),
    .B(_06479_),
    .Y(_06846_));
 AOI211x1_ASAP7_75t_R _29278_ (.A1(_06585_),
    .A2(_06774_),
    .B(_06433_),
    .C(_06729_),
    .Y(_06847_));
 NOR2x1_ASAP7_75t_SL _29279_ (.A(_06846_),
    .B(_06847_),
    .Y(_06848_));
 INVx1_ASAP7_75t_R _29280_ (.A(_06805_),
    .Y(_06849_));
 NAND2x1p5_ASAP7_75t_SL _29281_ (.A(_06513_),
    .B(_06578_),
    .Y(_06850_));
 OAI21x1_ASAP7_75t_SL _29282_ (.A1(_06513_),
    .A2(_06613_),
    .B(_06850_),
    .Y(_06851_));
 OAI21x1_ASAP7_75t_R _29283_ (.A1(_06849_),
    .A2(_06851_),
    .B(_06480_),
    .Y(_06852_));
 OA21x2_ASAP7_75t_SL _29284_ (.A1(_06723_),
    .A2(_06405_),
    .B(_06594_),
    .Y(_06853_));
 INVx1_ASAP7_75t_SL _29285_ (.A(_06499_),
    .Y(_06854_));
 AO21x1_ASAP7_75t_SL _29286_ (.A1(_06854_),
    .A2(_06644_),
    .B(_06469_),
    .Y(_06855_));
 NOR2x1_ASAP7_75t_SL _29287_ (.A(_06853_),
    .B(_06855_),
    .Y(_06856_));
 OAI21x1_ASAP7_75t_SL _29288_ (.A1(_06856_),
    .A2(_06852_),
    .B(_06509_),
    .Y(_06857_));
 OAI21x1_ASAP7_75t_SL _29289_ (.A1(_06848_),
    .A2(_06857_),
    .B(_06705_),
    .Y(_06858_));
 AND3x1_ASAP7_75t_L _29290_ (.A(_06675_),
    .B(_06513_),
    .C(_06490_),
    .Y(_06859_));
 OAI21x1_ASAP7_75t_R _29291_ (.A1(_06669_),
    .A2(_06549_),
    .B(_06469_),
    .Y(_06860_));
 NOR2x1_ASAP7_75t_R _29292_ (.A(_06859_),
    .B(_06860_),
    .Y(_06861_));
 INVx1_ASAP7_75t_SL _29293_ (.A(_06631_),
    .Y(_06862_));
 OAI21x1_ASAP7_75t_R _29294_ (.A1(_06405_),
    .A2(_06392_),
    .B(_06513_),
    .Y(_06863_));
 OAI21x1_ASAP7_75t_R _29295_ (.A1(_06584_),
    .A2(_06863_),
    .B(_06433_),
    .Y(_06864_));
 OAI21x1_ASAP7_75t_R _29296_ (.A1(_06862_),
    .A2(_06864_),
    .B(_06479_),
    .Y(_06865_));
 OAI21x1_ASAP7_75t_R _29297_ (.A1(_06428_),
    .A2(_06439_),
    .B(_06513_),
    .Y(_06866_));
 INVx1_ASAP7_75t_R _29298_ (.A(_06625_),
    .Y(_06867_));
 AOI21x1_ASAP7_75t_R _29299_ (.A1(_06866_),
    .A2(_06867_),
    .B(_06668_),
    .Y(_06868_));
 AOI21x1_ASAP7_75t_SL _29300_ (.A1(_06513_),
    .A2(_06831_),
    .B(_06542_),
    .Y(_06869_));
 AOI21x1_ASAP7_75t_R _29301_ (.A1(_06469_),
    .A2(_06869_),
    .B(_06479_),
    .Y(_06870_));
 OAI21x1_ASAP7_75t_R _29302_ (.A1(_06469_),
    .A2(_06868_),
    .B(_06870_),
    .Y(_06871_));
 OAI21x1_ASAP7_75t_SL _29303_ (.A1(_06861_),
    .A2(_06865_),
    .B(_06871_),
    .Y(_06872_));
 NOR2x1_ASAP7_75t_R _29304_ (.A(_06509_),
    .B(_06872_),
    .Y(_06873_));
 AOI21x1_ASAP7_75t_R _29305_ (.A1(_01366_),
    .A2(_06421_),
    .B(_06513_),
    .Y(_06874_));
 NOR2x1_ASAP7_75t_R _29306_ (.A(_06433_),
    .B(_06874_),
    .Y(_06875_));
 OA21x2_ASAP7_75t_R _29307_ (.A1(_06441_),
    .A2(_06448_),
    .B(_06875_),
    .Y(_06876_));
 OAI21x1_ASAP7_75t_R _29308_ (.A1(_06578_),
    .A2(_06728_),
    .B(_06433_),
    .Y(_06877_));
 AOI21x1_ASAP7_75t_R _29309_ (.A1(_06544_),
    .A2(_06545_),
    .B(_06877_),
    .Y(_06878_));
 OAI21x1_ASAP7_75t_R _29310_ (.A1(_06876_),
    .A2(_06878_),
    .B(_06538_),
    .Y(_06879_));
 NAND2x1_ASAP7_75t_SL _29311_ (.A(_06675_),
    .B(_06594_),
    .Y(_06880_));
 NAND2x1_ASAP7_75t_R _29312_ (.A(_06448_),
    .B(_06700_),
    .Y(_06881_));
 NAND2x1_ASAP7_75t_R _29313_ (.A(_06880_),
    .B(_06881_),
    .Y(_06882_));
 OA21x2_ASAP7_75t_R _29314_ (.A1(_01372_),
    .A2(_06513_),
    .B(_06433_),
    .Y(_06883_));
 AO21x1_ASAP7_75t_SL _29315_ (.A1(_06850_),
    .A2(_06883_),
    .B(_06538_),
    .Y(_06884_));
 AO21x1_ASAP7_75t_SL _29316_ (.A1(_06469_),
    .A2(_06882_),
    .B(_06884_),
    .Y(_06885_));
 AOI21x1_ASAP7_75t_SL _29317_ (.A1(_06885_),
    .A2(_06879_),
    .B(_06479_),
    .Y(_06886_));
 AOI21x1_ASAP7_75t_R _29318_ (.A1(_06818_),
    .A2(_06632_),
    .B(_06513_),
    .Y(_06887_));
 OAI21x1_ASAP7_75t_SL _29319_ (.A1(_06497_),
    .A2(_06529_),
    .B(_06469_),
    .Y(_06888_));
 NOR2x1_ASAP7_75t_R _29320_ (.A(_06887_),
    .B(_06888_),
    .Y(_06889_));
 AO21x1_ASAP7_75t_R _29321_ (.A1(_06421_),
    .A2(_06513_),
    .B(_06469_),
    .Y(_06890_));
 NOR2x1_ASAP7_75t_R _29322_ (.A(_06518_),
    .B(_06465_),
    .Y(_06891_));
 OAI21x1_ASAP7_75t_R _29323_ (.A1(_06890_),
    .A2(_06891_),
    .B(_06538_),
    .Y(_06892_));
 OAI21x1_ASAP7_75t_R _29324_ (.A1(_06889_),
    .A2(_06892_),
    .B(_06479_),
    .Y(_06893_));
 INVx1_ASAP7_75t_R _29325_ (.A(_06600_),
    .Y(_06894_));
 AOI21x1_ASAP7_75t_R _29326_ (.A1(_06608_),
    .A2(_06690_),
    .B(_06448_),
    .Y(_06895_));
 OAI21x1_ASAP7_75t_R _29327_ (.A1(_06894_),
    .A2(_06895_),
    .B(_06433_),
    .Y(_06896_));
 NAND2x1_ASAP7_75t_R _29328_ (.A(_06513_),
    .B(_06831_),
    .Y(_06897_));
 NOR2x1_ASAP7_75t_R _29329_ (.A(_06520_),
    .B(_06897_),
    .Y(_06898_));
 INVx1_ASAP7_75t_SL _29330_ (.A(_06688_),
    .Y(_06899_));
 NOR2x1_ASAP7_75t_SL _29331_ (.A(_06740_),
    .B(_06899_),
    .Y(_06900_));
 OAI21x1_ASAP7_75t_R _29332_ (.A1(_06898_),
    .A2(_06900_),
    .B(_06469_),
    .Y(_06901_));
 AOI21x1_ASAP7_75t_R _29333_ (.A1(_06896_),
    .A2(_06901_),
    .B(_06538_),
    .Y(_06902_));
 OAI21x1_ASAP7_75t_R _29334_ (.A1(_06893_),
    .A2(_06902_),
    .B(_06561_),
    .Y(_06903_));
 OAI22x1_ASAP7_75t_SL _29335_ (.A1(_06858_),
    .A2(_06873_),
    .B1(_06903_),
    .B2(_06886_),
    .Y(_00148_));
 OAI21x1_ASAP7_75t_R _29336_ (.A1(_06739_),
    .A2(_06488_),
    .B(_06513_),
    .Y(_06904_));
 INVx2_ASAP7_75t_L _29337_ (.A(_06518_),
    .Y(_06905_));
 NAND2x1p5_ASAP7_75t_SL _29338_ (.A(_06822_),
    .B(_06905_),
    .Y(_06906_));
 AOI21x1_ASAP7_75t_SL _29339_ (.A1(_06904_),
    .A2(_06906_),
    .B(_06433_),
    .Y(_06907_));
 NAND2x1_ASAP7_75t_R _29340_ (.A(_01370_),
    .B(_06513_),
    .Y(_06908_));
 NOR2x1_ASAP7_75t_R _29341_ (.A(_06513_),
    .B(_06405_),
    .Y(_06909_));
 NOR2x1_ASAP7_75t_SL _29342_ (.A(_06909_),
    .B(_06606_),
    .Y(_06910_));
 AOI21x1_ASAP7_75t_R _29343_ (.A1(_06908_),
    .A2(_06910_),
    .B(_06469_),
    .Y(_06911_));
 OAI21x1_ASAP7_75t_SL _29344_ (.A1(_06911_),
    .A2(_06907_),
    .B(_06479_),
    .Y(_06912_));
 AND3x1_ASAP7_75t_R _29345_ (.A(_06428_),
    .B(_01366_),
    .C(_01368_),
    .Y(_06913_));
 OAI21x1_ASAP7_75t_R _29346_ (.A1(_06448_),
    .A2(_06913_),
    .B(_06433_),
    .Y(_06914_));
 NOR2x1_ASAP7_75t_SL _29347_ (.A(_06513_),
    .B(_06623_),
    .Y(_06915_));
 INVx1_ASAP7_75t_SL _29348_ (.A(_06676_),
    .Y(_06916_));
 AOI21x1_ASAP7_75t_R _29349_ (.A1(_06448_),
    .A2(_06566_),
    .B(_06433_),
    .Y(_06917_));
 AOI21x1_ASAP7_75t_R _29350_ (.A1(_06916_),
    .A2(_06917_),
    .B(_06479_),
    .Y(_06918_));
 OAI21x1_ASAP7_75t_R _29351_ (.A1(_06914_),
    .A2(_06915_),
    .B(_06918_),
    .Y(_06919_));
 NAND3x1_ASAP7_75t_SL _29352_ (.A(_06919_),
    .B(_06509_),
    .C(_06912_),
    .Y(_06920_));
 OA21x2_ASAP7_75t_R _29353_ (.A1(_06487_),
    .A2(_06448_),
    .B(_06469_),
    .Y(_06921_));
 OAI21x1_ASAP7_75t_R _29354_ (.A1(_06909_),
    .A2(_06606_),
    .B(_06905_),
    .Y(_06922_));
 AOI21x1_ASAP7_75t_R _29355_ (.A1(_06921_),
    .A2(_06922_),
    .B(_06480_),
    .Y(_06923_));
 AO21x1_ASAP7_75t_SL _29356_ (.A1(_06720_),
    .A2(_06608_),
    .B(_06513_),
    .Y(_06924_));
 NAND2x1_ASAP7_75t_SL _29357_ (.A(_06924_),
    .B(_06547_),
    .Y(_06925_));
 NAND2x1_ASAP7_75t_R _29358_ (.A(_06923_),
    .B(_06925_),
    .Y(_06926_));
 AOI21x1_ASAP7_75t_R _29359_ (.A1(_06675_),
    .A2(_06712_),
    .B(_06433_),
    .Y(_06927_));
 OAI21x1_ASAP7_75t_L _29360_ (.A1(_06515_),
    .A2(_06531_),
    .B(_06927_),
    .Y(_06928_));
 NOR2x1_ASAP7_75t_R _29361_ (.A(_06448_),
    .B(_06424_),
    .Y(_06929_));
 AOI21x1_ASAP7_75t_R _29362_ (.A1(_06690_),
    .A2(_06628_),
    .B(_06929_),
    .Y(_06930_));
 AOI21x1_ASAP7_75t_R _29363_ (.A1(_06433_),
    .A2(_06930_),
    .B(_06479_),
    .Y(_06931_));
 AOI21x1_ASAP7_75t_R _29364_ (.A1(_06928_),
    .A2(_06931_),
    .B(_06509_),
    .Y(_06932_));
 AOI21x1_ASAP7_75t_L _29365_ (.A1(_06926_),
    .A2(_06932_),
    .B(_06705_),
    .Y(_06933_));
 NAND2x1_ASAP7_75t_SL _29366_ (.A(_06933_),
    .B(_06920_),
    .Y(_06934_));
 NAND2x1_ASAP7_75t_SL _29367_ (.A(_06723_),
    .B(_06874_),
    .Y(_06935_));
 AOI21x1_ASAP7_75t_R _29368_ (.A1(_06850_),
    .A2(_06935_),
    .B(_06433_),
    .Y(_06936_));
 NOR2x1_ASAP7_75t_L _29369_ (.A(_06457_),
    .B(_06515_),
    .Y(_06937_));
 AO21x1_ASAP7_75t_R _29370_ (.A1(_06718_),
    .A2(_06448_),
    .B(_06469_),
    .Y(_06938_));
 NOR2x1_ASAP7_75t_R _29371_ (.A(_06937_),
    .B(_06938_),
    .Y(_06939_));
 OAI21x1_ASAP7_75t_R _29372_ (.A1(_06936_),
    .A2(_06939_),
    .B(_06479_),
    .Y(_06940_));
 AO21x1_ASAP7_75t_R _29373_ (.A1(_06439_),
    .A2(_06513_),
    .B(_06469_),
    .Y(_06941_));
 NOR2x1_ASAP7_75t_R _29374_ (.A(_06941_),
    .B(_06900_),
    .Y(_06942_));
 OAI21x1_ASAP7_75t_R _29375_ (.A1(_06421_),
    .A2(_06392_),
    .B(_06513_),
    .Y(_06943_));
 OAI21x1_ASAP7_75t_R _29376_ (.A1(_06405_),
    .A2(_06421_),
    .B(_06487_),
    .Y(_06944_));
 NOR2x1_ASAP7_75t_SL _29377_ (.A(_06943_),
    .B(_06944_),
    .Y(_06945_));
 OAI21x1_ASAP7_75t_R _29378_ (.A1(_06669_),
    .A2(_06533_),
    .B(_06469_),
    .Y(_06946_));
 NOR2x1_ASAP7_75t_SL _29379_ (.A(_06945_),
    .B(_06946_),
    .Y(_06947_));
 OAI21x1_ASAP7_75t_R _29380_ (.A1(_06942_),
    .A2(_06947_),
    .B(_06480_),
    .Y(_06948_));
 AOI21x1_ASAP7_75t_R _29381_ (.A1(_06940_),
    .A2(_06948_),
    .B(_06538_),
    .Y(_06949_));
 AOI21x1_ASAP7_75t_SL _29382_ (.A1(_06424_),
    .A2(_06687_),
    .B(_06469_),
    .Y(_06950_));
 INVx1_ASAP7_75t_R _29383_ (.A(_06787_),
    .Y(_06951_));
 NAND3x1_ASAP7_75t_SL _29384_ (.A(_06950_),
    .B(_06453_),
    .C(_06951_),
    .Y(_06952_));
 AND2x2_ASAP7_75t_SL _29385_ (.A(_06728_),
    .B(_06469_),
    .Y(_06953_));
 AOI21x1_ASAP7_75t_SL _29386_ (.A1(_06689_),
    .A2(_06953_),
    .B(_06480_),
    .Y(_06954_));
 NAND2x1_ASAP7_75t_SL _29387_ (.A(_06952_),
    .B(_06954_),
    .Y(_06955_));
 NAND2x1_ASAP7_75t_SL _29388_ (.A(_06602_),
    .B(_06905_),
    .Y(_06956_));
 AOI21x1_ASAP7_75t_R _29389_ (.A1(_06956_),
    .A2(_06543_),
    .B(_06469_),
    .Y(_06957_));
 OAI21x1_ASAP7_75t_R _29390_ (.A1(_06527_),
    .A2(_06542_),
    .B(_06513_),
    .Y(_06958_));
 OAI21x1_ASAP7_75t_R _29391_ (.A1(_06421_),
    .A2(_06688_),
    .B(_06712_),
    .Y(_06959_));
 AOI21x1_ASAP7_75t_R _29392_ (.A1(_06958_),
    .A2(_06959_),
    .B(_06433_),
    .Y(_06960_));
 OAI21x1_ASAP7_75t_R _29393_ (.A1(_06957_),
    .A2(_06960_),
    .B(_06480_),
    .Y(_06961_));
 AOI21x1_ASAP7_75t_SL _29394_ (.A1(_06961_),
    .A2(_06955_),
    .B(_06509_),
    .Y(_06962_));
 OAI21x1_ASAP7_75t_SL _29395_ (.A1(_06949_),
    .A2(_06962_),
    .B(_06705_),
    .Y(_06963_));
 NAND2x1_ASAP7_75t_SL _29396_ (.A(_06934_),
    .B(_06963_),
    .Y(_00149_));
 NAND2x1_ASAP7_75t_SL _29397_ (.A(_06448_),
    .B(_06439_),
    .Y(_06964_));
 AOI21x1_ASAP7_75t_SL _29398_ (.A1(_06964_),
    .A2(_06814_),
    .B(_06469_),
    .Y(_06965_));
 AO21x1_ASAP7_75t_SL _29399_ (.A1(_06405_),
    .A2(_06421_),
    .B(_06433_),
    .Y(_06966_));
 NOR2x1_ASAP7_75t_SL _29400_ (.A(_06644_),
    .B(_06769_),
    .Y(_06967_));
 OAI21x1_ASAP7_75t_SL _29401_ (.A1(_06966_),
    .A2(_06967_),
    .B(_06480_),
    .Y(_06968_));
 OAI21x1_ASAP7_75t_SL _29402_ (.A1(_06965_),
    .A2(_06968_),
    .B(_06538_),
    .Y(_06969_));
 NOR2x1_ASAP7_75t_SL _29403_ (.A(_06433_),
    .B(_06695_),
    .Y(_06970_));
 NAND2x1_ASAP7_75t_SL _29404_ (.A(_06970_),
    .B(_06523_),
    .Y(_06971_));
 AO21x1_ASAP7_75t_SL _29405_ (.A1(_06513_),
    .A2(_06717_),
    .B(_06822_),
    .Y(_06972_));
 NAND2x1_ASAP7_75t_SL _29406_ (.A(_06972_),
    .B(_06950_),
    .Y(_06973_));
 AOI21x1_ASAP7_75t_SL _29407_ (.A1(_06971_),
    .A2(_06973_),
    .B(_06480_),
    .Y(_06974_));
 OAI21x1_ASAP7_75t_SL _29408_ (.A1(_06974_),
    .A2(_06969_),
    .B(_06561_),
    .Y(_06975_));
 INVx1_ASAP7_75t_SL _29409_ (.A(_06587_),
    .Y(_06976_));
 AOI21x1_ASAP7_75t_SL _29410_ (.A1(_06976_),
    .A2(_06880_),
    .B(_06433_),
    .Y(_06977_));
 OAI21x1_ASAP7_75t_SL _29411_ (.A1(_06977_),
    .A2(_06736_),
    .B(_06479_),
    .Y(_06978_));
 OA21x2_ASAP7_75t_SL _29412_ (.A1(_06440_),
    .A2(_06513_),
    .B(_06469_),
    .Y(_06979_));
 OAI21x1_ASAP7_75t_SL _29413_ (.A1(_06739_),
    .A2(_06916_),
    .B(_06979_),
    .Y(_06980_));
 AND2x2_ASAP7_75t_SL _29414_ (.A(_06712_),
    .B(_06675_),
    .Y(_06981_));
 AO21x1_ASAP7_75t_SL _29415_ (.A1(_01376_),
    .A2(_06513_),
    .B(_06469_),
    .Y(_06982_));
 OA21x2_ASAP7_75t_SL _29416_ (.A1(_06981_),
    .A2(_06982_),
    .B(_06480_),
    .Y(_06983_));
 NAND2x1_ASAP7_75t_SL _29417_ (.A(_06980_),
    .B(_06983_),
    .Y(_06984_));
 AOI21x1_ASAP7_75t_SL _29418_ (.A1(_06978_),
    .A2(_06984_),
    .B(_06538_),
    .Y(_06985_));
 NOR2x1_ASAP7_75t_SL _29419_ (.A(_06985_),
    .B(_06975_),
    .Y(_06986_));
 AO21x1_ASAP7_75t_R _29420_ (.A1(_01375_),
    .A2(_01381_),
    .B(_06513_),
    .Y(_06987_));
 AND2x2_ASAP7_75t_SL _29421_ (.A(_06987_),
    .B(_06433_),
    .Y(_06988_));
 OAI21x1_ASAP7_75t_SL _29422_ (.A1(_06899_),
    .A2(_06707_),
    .B(_06988_),
    .Y(_06989_));
 OAI21x1_ASAP7_75t_R _29423_ (.A1(_06448_),
    .A2(_06569_),
    .B(_06469_),
    .Y(_06990_));
 INVx1_ASAP7_75t_SL _29424_ (.A(_06990_),
    .Y(_06991_));
 NOR2x1_ASAP7_75t_SL _29425_ (.A(_06493_),
    .B(_06787_),
    .Y(_06992_));
 AOI21x1_ASAP7_75t_SL _29426_ (.A1(_06991_),
    .A2(_06992_),
    .B(_06479_),
    .Y(_06993_));
 AOI21x1_ASAP7_75t_SL _29427_ (.A1(_06989_),
    .A2(_06993_),
    .B(_06509_),
    .Y(_06994_));
 AOI21x1_ASAP7_75t_SL _29428_ (.A1(_06551_),
    .A2(_06712_),
    .B(_06469_),
    .Y(_06995_));
 OAI21x1_ASAP7_75t_SL _29429_ (.A1(_06542_),
    .A2(_06646_),
    .B(_06513_),
    .Y(_06996_));
 NAND2x1_ASAP7_75t_SL _29430_ (.A(_06995_),
    .B(_06996_),
    .Y(_06997_));
 NAND2x1_ASAP7_75t_SL _29431_ (.A(_06608_),
    .B(_06579_),
    .Y(_06998_));
 AOI21x1_ASAP7_75t_R _29432_ (.A1(_06720_),
    .A2(_06717_),
    .B(_06448_),
    .Y(_06999_));
 NOR2x1_ASAP7_75t_SL _29433_ (.A(_06999_),
    .B(_06990_),
    .Y(_07000_));
 AOI21x1_ASAP7_75t_SL _29434_ (.A1(_06998_),
    .A2(_07000_),
    .B(_06480_),
    .Y(_07001_));
 NAND2x1_ASAP7_75t_SL _29435_ (.A(_06997_),
    .B(_07001_),
    .Y(_07002_));
 NAND2x1_ASAP7_75t_SL _29436_ (.A(_06994_),
    .B(_07002_),
    .Y(_07003_));
 AOI21x1_ASAP7_75t_SL _29437_ (.A1(_06751_),
    .A2(_06744_),
    .B(_06498_),
    .Y(_07004_));
 AOI21x1_ASAP7_75t_SL _29438_ (.A1(_06643_),
    .A2(_06822_),
    .B(_06469_),
    .Y(_07005_));
 OAI21x1_ASAP7_75t_SL _29439_ (.A1(_06584_),
    .A2(_06521_),
    .B(_06513_),
    .Y(_07006_));
 AOI21x1_ASAP7_75t_SL _29440_ (.A1(_07005_),
    .A2(_07006_),
    .B(_06479_),
    .Y(_07007_));
 OAI21x1_ASAP7_75t_SL _29441_ (.A1(_06433_),
    .A2(_07004_),
    .B(_07007_),
    .Y(_07008_));
 OA21x2_ASAP7_75t_SL _29442_ (.A1(_06487_),
    .A2(_06513_),
    .B(_06469_),
    .Y(_07009_));
 OAI21x1_ASAP7_75t_SL _29443_ (.A1(_06439_),
    .A2(_06520_),
    .B(_06513_),
    .Y(_07010_));
 AOI21x1_ASAP7_75t_SL _29444_ (.A1(_07009_),
    .A2(_07010_),
    .B(_06480_),
    .Y(_07011_));
 OAI21x1_ASAP7_75t_SL _29445_ (.A1(_06520_),
    .A2(_06462_),
    .B(_06513_),
    .Y(_07012_));
 OAI21x1_ASAP7_75t_SL _29446_ (.A1(_06499_),
    .A2(_06759_),
    .B(_06448_),
    .Y(_07013_));
 NAND3x1_ASAP7_75t_SL _29447_ (.A(_07012_),
    .B(_06950_),
    .C(_07013_),
    .Y(_07014_));
 AOI21x1_ASAP7_75t_SL _29448_ (.A1(_07011_),
    .A2(_07014_),
    .B(_06538_),
    .Y(_07015_));
 NAND2x1_ASAP7_75t_SL _29449_ (.A(_07008_),
    .B(_07015_),
    .Y(_07016_));
 AOI21x1_ASAP7_75t_SL _29450_ (.A1(_07003_),
    .A2(_07016_),
    .B(_06561_),
    .Y(_07017_));
 NOR2x1_ASAP7_75t_SL _29451_ (.A(_06986_),
    .B(_07017_),
    .Y(_00150_));
 NOR2x1_ASAP7_75t_R _29452_ (.A(_06469_),
    .B(_06644_),
    .Y(_07018_));
 AOI21x1_ASAP7_75t_R _29453_ (.A1(_06880_),
    .A2(_07018_),
    .B(_06479_),
    .Y(_07019_));
 OAI21x1_ASAP7_75t_R _29454_ (.A1(_06492_),
    .A2(_06646_),
    .B(_06513_),
    .Y(_07020_));
 AOI21x1_ASAP7_75t_R _29455_ (.A1(_06651_),
    .A2(_06585_),
    .B(_06433_),
    .Y(_07021_));
 NAND2x1_ASAP7_75t_R _29456_ (.A(_07020_),
    .B(_07021_),
    .Y(_07022_));
 AOI21x1_ASAP7_75t_R _29457_ (.A1(_07019_),
    .A2(_07022_),
    .B(_06705_),
    .Y(_07023_));
 AOI21x1_ASAP7_75t_R _29458_ (.A1(_06775_),
    .A2(_06995_),
    .B(_06480_),
    .Y(_07024_));
 AO21x1_ASAP7_75t_SL _29459_ (.A1(_06551_),
    .A2(_06500_),
    .B(_06433_),
    .Y(_07025_));
 AO21x1_ASAP7_75t_SL _29460_ (.A1(_06452_),
    .A2(_06651_),
    .B(_07025_),
    .Y(_07026_));
 NAND2x1_ASAP7_75t_SL _29461_ (.A(_07026_),
    .B(_07024_),
    .Y(_07027_));
 NAND2x1_ASAP7_75t_SL _29462_ (.A(_07027_),
    .B(_07023_),
    .Y(_07028_));
 NAND2x1_ASAP7_75t_L _29463_ (.A(_06636_),
    .B(_06606_),
    .Y(_07029_));
 AOI21x1_ASAP7_75t_R _29464_ (.A1(_06800_),
    .A2(_07029_),
    .B(_06433_),
    .Y(_07030_));
 NOR2x1_ASAP7_75t_R _29465_ (.A(_06492_),
    .B(_06646_),
    .Y(_07031_));
 OAI21x1_ASAP7_75t_R _29466_ (.A1(_06488_),
    .A2(_06515_),
    .B(_06433_),
    .Y(_07032_));
 AOI21x1_ASAP7_75t_SL _29467_ (.A1(_06448_),
    .A2(_07031_),
    .B(_07032_),
    .Y(_07033_));
 OAI21x1_ASAP7_75t_R _29468_ (.A1(_07030_),
    .A2(_07033_),
    .B(_06480_),
    .Y(_07034_));
 AO21x1_ASAP7_75t_R _29469_ (.A1(_06527_),
    .A2(_06448_),
    .B(_06433_),
    .Y(_07035_));
 AO21x1_ASAP7_75t_R _29470_ (.A1(_06688_),
    .A2(_06774_),
    .B(_07035_),
    .Y(_07036_));
 NOR2x1_ASAP7_75t_R _29471_ (.A(_06492_),
    .B(_06469_),
    .Y(_07037_));
 OAI21x1_ASAP7_75t_R _29472_ (.A1(_06513_),
    .A2(_06570_),
    .B(_06707_),
    .Y(_07038_));
 AOI21x1_ASAP7_75t_R _29473_ (.A1(_07037_),
    .A2(_07038_),
    .B(_06480_),
    .Y(_07039_));
 AOI21x1_ASAP7_75t_R _29474_ (.A1(_07036_),
    .A2(_07039_),
    .B(_06561_),
    .Y(_07040_));
 AOI21x1_ASAP7_75t_R _29475_ (.A1(_07034_),
    .A2(_07040_),
    .B(_06509_),
    .Y(_07041_));
 NAND2x1_ASAP7_75t_SL _29476_ (.A(_07028_),
    .B(_07041_),
    .Y(_07042_));
 NOR2x1_ASAP7_75t_R _29477_ (.A(_06549_),
    .B(_06441_),
    .Y(_07043_));
 AO21x1_ASAP7_75t_SL _29478_ (.A1(_06695_),
    .A2(_06624_),
    .B(_06909_),
    .Y(_07044_));
 AOI21x1_ASAP7_75t_R _29479_ (.A1(_06469_),
    .A2(_07044_),
    .B(_06479_),
    .Y(_07045_));
 OA21x2_ASAP7_75t_SL _29480_ (.A1(_06864_),
    .A2(_07043_),
    .B(_07045_),
    .Y(_07046_));
 AOI211x1_ASAP7_75t_R _29481_ (.A1(_06636_),
    .A2(_06828_),
    .B(_06498_),
    .C(_06469_),
    .Y(_07047_));
 OA21x2_ASAP7_75t_SL _29482_ (.A1(_06439_),
    .A2(_06440_),
    .B(_06822_),
    .Y(_07048_));
 AO21x1_ASAP7_75t_R _29483_ (.A1(_06585_),
    .A2(_06513_),
    .B(_06433_),
    .Y(_07049_));
 OAI21x1_ASAP7_75t_R _29484_ (.A1(_07048_),
    .A2(_07049_),
    .B(_06479_),
    .Y(_07050_));
 OAI21x1_ASAP7_75t_R _29485_ (.A1(_07047_),
    .A2(_07050_),
    .B(_06561_),
    .Y(_07051_));
 AOI21x1_ASAP7_75t_SL _29486_ (.A1(_06500_),
    .A2(_06756_),
    .B(_06433_),
    .Y(_07052_));
 OAI21x1_ASAP7_75t_SL _29487_ (.A1(_06694_),
    .A2(_06533_),
    .B(_07052_),
    .Y(_07053_));
 NAND2x1_ASAP7_75t_R _29488_ (.A(_06448_),
    .B(_06499_),
    .Y(_07054_));
 OAI21x1_ASAP7_75t_R _29489_ (.A1(_01381_),
    .A2(_06448_),
    .B(_06433_),
    .Y(_07055_));
 AOI21x1_ASAP7_75t_R _29490_ (.A1(_06448_),
    .A2(_06612_),
    .B(_07055_),
    .Y(_07056_));
 AOI21x1_ASAP7_75t_R _29491_ (.A1(_07054_),
    .A2(_07056_),
    .B(_06480_),
    .Y(_07057_));
 NAND2x1_ASAP7_75t_L _29492_ (.A(_07053_),
    .B(_07057_),
    .Y(_07058_));
 AOI21x1_ASAP7_75t_R _29493_ (.A1(_01372_),
    .A2(_06513_),
    .B(_06469_),
    .Y(_07059_));
 AOI21x1_ASAP7_75t_R _29494_ (.A1(_07059_),
    .A2(_06571_),
    .B(_06479_),
    .Y(_07060_));
 AO21x1_ASAP7_75t_R _29495_ (.A1(_06608_),
    .A2(_06392_),
    .B(_06513_),
    .Y(_07061_));
 INVx1_ASAP7_75t_SL _29496_ (.A(_06888_),
    .Y(_07062_));
 NAND2x1_ASAP7_75t_SL _29497_ (.A(_07061_),
    .B(_07062_),
    .Y(_07063_));
 AOI21x1_ASAP7_75t_SL _29498_ (.A1(_07060_),
    .A2(_07063_),
    .B(_06561_),
    .Y(_07064_));
 AOI21x1_ASAP7_75t_SL _29499_ (.A1(_07064_),
    .A2(_07058_),
    .B(_06538_),
    .Y(_07065_));
 OAI21x1_ASAP7_75t_SL _29500_ (.A1(_07046_),
    .A2(_07051_),
    .B(_07065_),
    .Y(_07066_));
 NAND2x1_ASAP7_75t_SL _29501_ (.A(_07066_),
    .B(_07042_),
    .Y(_00151_));
 NOR2x1_ASAP7_75t_R _29502_ (.A(_00574_),
    .B(_00408_),
    .Y(_07067_));
 XOR2x2_ASAP7_75t_L _29503_ (.A(_12768_),
    .B(_00664_),
    .Y(_07068_));
 XOR2x2_ASAP7_75t_L _29504_ (.A(_12805_),
    .B(_04364_),
    .Y(_07069_));
 NAND2x1_ASAP7_75t_SL _29505_ (.A(_07068_),
    .B(_07069_),
    .Y(_07070_));
 XNOR2x2_ASAP7_75t_SL _29506_ (.A(_00664_),
    .B(_12768_),
    .Y(_07071_));
 XOR2x2_ASAP7_75t_L _29507_ (.A(_12807_),
    .B(_04364_),
    .Y(_07072_));
 NAND2x1p5_ASAP7_75t_L _29508_ (.A(_07071_),
    .B(_07072_),
    .Y(_07073_));
 AOI21x1_ASAP7_75t_SL _29509_ (.A1(_07070_),
    .A2(_07073_),
    .B(_10675_),
    .Y(_07074_));
 OAI21x1_ASAP7_75t_R _29510_ (.A1(_07067_),
    .A2(_07074_),
    .B(_00945_),
    .Y(_07075_));
 AND2x2_ASAP7_75t_R _29511_ (.A(_10675_),
    .B(_00408_),
    .Y(_07076_));
 NAND2x1_ASAP7_75t_L _29512_ (.A(_07068_),
    .B(_07072_),
    .Y(_07077_));
 NAND2x1_ASAP7_75t_L _29513_ (.A(_07071_),
    .B(_07069_),
    .Y(_07078_));
 AOI21x1_ASAP7_75t_SL _29514_ (.A1(_07077_),
    .A2(_07078_),
    .B(_10675_),
    .Y(_07079_));
 OAI21x1_ASAP7_75t_R _29515_ (.A1(_07076_),
    .A2(_07079_),
    .B(_08867_),
    .Y(_07080_));
 NAND2x2_ASAP7_75t_SL _29516_ (.A(_07075_),
    .B(_07080_),
    .Y(_07081_));
 NOR2x1_ASAP7_75t_L _29518_ (.A(_00574_),
    .B(_00409_),
    .Y(_07082_));
 XOR2x2_ASAP7_75t_SL _29519_ (.A(_12768_),
    .B(_12791_),
    .Y(_07083_));
 NAND2x1_ASAP7_75t_L _29520_ (.A(_00569_),
    .B(_07083_),
    .Y(_07084_));
 XOR2x2_ASAP7_75t_SL _29521_ (.A(_12774_),
    .B(_12791_),
    .Y(_07085_));
 NAND2x1_ASAP7_75t_L _29522_ (.A(_04537_),
    .B(_07085_),
    .Y(_07086_));
 AOI21x1_ASAP7_75t_SL _29523_ (.A1(_07086_),
    .A2(_07084_),
    .B(_10675_),
    .Y(_07087_));
 OAI21x1_ASAP7_75t_R _29524_ (.A1(_07082_),
    .A2(_07087_),
    .B(_00934_),
    .Y(_07088_));
 AND2x2_ASAP7_75t_L _29525_ (.A(_10675_),
    .B(_00409_),
    .Y(_07089_));
 NAND2x1_ASAP7_75t_L _29526_ (.A(_04537_),
    .B(_07083_),
    .Y(_07090_));
 NAND2x1_ASAP7_75t_L _29527_ (.A(_00569_),
    .B(_07085_),
    .Y(_07091_));
 AOI21x1_ASAP7_75t_SL _29528_ (.A1(_07091_),
    .A2(_07090_),
    .B(_10675_),
    .Y(_07092_));
 OAI21x1_ASAP7_75t_R _29529_ (.A1(_07089_),
    .A2(_07092_),
    .B(_08862_),
    .Y(_07093_));
 NAND2x1p5_ASAP7_75t_SL _29530_ (.A(_07088_),
    .B(_07093_),
    .Y(_07094_));
 XOR2x2_ASAP7_75t_L _29532_ (.A(_00600_),
    .B(_00665_),
    .Y(_07095_));
 NAND2x1_ASAP7_75t_SL _29533_ (.A(_12772_),
    .B(_07095_),
    .Y(_07096_));
 XNOR2x2_ASAP7_75t_L _29534_ (.A(_00600_),
    .B(_00665_),
    .Y(_07097_));
 NAND2x1_ASAP7_75t_R _29535_ (.A(_00696_),
    .B(_07097_),
    .Y(_07098_));
 AOI21x1_ASAP7_75t_SL _29536_ (.A1(_07096_),
    .A2(_07098_),
    .B(_04390_),
    .Y(_07099_));
 XOR2x2_ASAP7_75t_SL _29537_ (.A(_00665_),
    .B(_00696_),
    .Y(_07100_));
 NAND2x1_ASAP7_75t_R _29538_ (.A(_00600_),
    .B(_07100_),
    .Y(_07101_));
 XNOR2x2_ASAP7_75t_SL _29539_ (.A(_00665_),
    .B(_00696_),
    .Y(_07102_));
 NAND2x1_ASAP7_75t_R _29540_ (.A(_01578_),
    .B(_07102_),
    .Y(_07103_));
 AOI21x1_ASAP7_75t_R _29541_ (.A1(_07101_),
    .A2(_07103_),
    .B(_04389_),
    .Y(_07104_));
 OAI21x1_ASAP7_75t_SL _29542_ (.A1(_07099_),
    .A2(_07104_),
    .B(_00574_),
    .Y(_07105_));
 NOR2x1_ASAP7_75t_R _29543_ (.A(_00574_),
    .B(_00410_),
    .Y(_07106_));
 INVx1_ASAP7_75t_R _29544_ (.A(_07106_),
    .Y(_07107_));
 NAND3x1_ASAP7_75t_SL _29545_ (.A(_07105_),
    .B(_00956_),
    .C(_07107_),
    .Y(_07108_));
 INVx2_ASAP7_75t_SL _29546_ (.A(_07105_),
    .Y(_07109_));
 INVx1_ASAP7_75t_R _29547_ (.A(_00956_),
    .Y(_07110_));
 OAI21x1_ASAP7_75t_SL _29548_ (.A1(_07106_),
    .A2(_07109_),
    .B(_07110_),
    .Y(_07111_));
 NAND2x1_ASAP7_75t_SL _29549_ (.A(_07108_),
    .B(_07111_),
    .Y(_07112_));
 OAI21x1_ASAP7_75t_SL _29552_ (.A1(_07092_),
    .A2(_07089_),
    .B(_00934_),
    .Y(_07114_));
 OAI21x1_ASAP7_75t_SL _29553_ (.A1(_07087_),
    .A2(_07082_),
    .B(_08862_),
    .Y(_07115_));
 NAND2x2_ASAP7_75t_SL _29554_ (.A(_07115_),
    .B(_07114_),
    .Y(_07116_));
 NAND3x1_ASAP7_75t_L _29556_ (.A(_07105_),
    .B(_07110_),
    .C(_07107_),
    .Y(_07117_));
 OAI21x1_ASAP7_75t_SL _29557_ (.A1(_07106_),
    .A2(_07109_),
    .B(_00956_),
    .Y(_07118_));
 NAND2x2_ASAP7_75t_SL _29558_ (.A(_07117_),
    .B(_07118_),
    .Y(_07119_));
 AO21x2_ASAP7_75t_SL _29561_ (.A1(_07118_),
    .A2(_07117_),
    .B(_01386_),
    .Y(_07121_));
 INVx2_ASAP7_75t_SL _29562_ (.A(_01385_),
    .Y(_07122_));
 AO21x1_ASAP7_75t_R _29563_ (.A1(_07111_),
    .A2(_07108_),
    .B(_07122_),
    .Y(_07123_));
 XNOR2x2_ASAP7_75t_SL _29564_ (.A(_04415_),
    .B(_04414_),
    .Y(_07124_));
 XOR2x2_ASAP7_75t_SL _29565_ (.A(_12833_),
    .B(_00666_),
    .Y(_07125_));
 AND2x2_ASAP7_75t_SL _29566_ (.A(_07124_),
    .B(_07125_),
    .Y(_07126_));
 OAI21x1_ASAP7_75t_SL _29567_ (.A1(_07125_),
    .A2(_07124_),
    .B(_00574_),
    .Y(_07127_));
 NAND2x1_ASAP7_75t_SL _29568_ (.A(_00529_),
    .B(_10675_),
    .Y(_07128_));
 OAI21x1_ASAP7_75t_SL _29569_ (.A1(_07126_),
    .A2(_07127_),
    .B(_07128_),
    .Y(_07129_));
 XOR2x2_ASAP7_75t_SL _29570_ (.A(_07129_),
    .B(_08880_),
    .Y(_07130_));
 AO21x1_ASAP7_75t_SL _29573_ (.A1(_07121_),
    .A2(_07123_),
    .B(_07130_),
    .Y(_07133_));
 INVx1_ASAP7_75t_R _29574_ (.A(_01391_),
    .Y(_07134_));
 AO21x1_ASAP7_75t_SL _29575_ (.A1(_07111_),
    .A2(_07108_),
    .B(_07134_),
    .Y(_07135_));
 AO21x1_ASAP7_75t_R _29576_ (.A1(_07118_),
    .A2(_07117_),
    .B(_07122_),
    .Y(_07136_));
 XOR2x2_ASAP7_75t_SL _29578_ (.A(_07129_),
    .B(_00959_),
    .Y(_07138_));
 AO21x1_ASAP7_75t_SL _29581_ (.A1(_07135_),
    .A2(_07136_),
    .B(_07138_),
    .Y(_07141_));
 XOR2x2_ASAP7_75t_SL _29582_ (.A(_12850_),
    .B(_00667_),
    .Y(_07142_));
 XOR2x2_ASAP7_75t_L _29583_ (.A(_04437_),
    .B(_07142_),
    .Y(_07143_));
 NOR2x1_ASAP7_75t_R _29584_ (.A(_00574_),
    .B(_00523_),
    .Y(_07144_));
 AOI21x1_ASAP7_75t_R _29585_ (.A1(_00574_),
    .A2(_07143_),
    .B(_07144_),
    .Y(_07145_));
 XNOR2x2_ASAP7_75t_SL _29586_ (.A(_00960_),
    .B(_07145_),
    .Y(_07146_));
 INVx3_ASAP7_75t_SL _29587_ (.A(_07146_),
    .Y(_07147_));
 AO21x1_ASAP7_75t_SL _29590_ (.A1(_07133_),
    .A2(_07141_),
    .B(_07147_),
    .Y(_07150_));
 NAND2x1_ASAP7_75t_SL _29592_ (.A(_07112_),
    .B(_07081_),
    .Y(_07152_));
 AO21x1_ASAP7_75t_SL _29593_ (.A1(_07152_),
    .A2(_07121_),
    .B(_07138_),
    .Y(_07153_));
 INVx1_ASAP7_75t_SL _29595_ (.A(_01386_),
    .Y(_07155_));
 NOR2x1_ASAP7_75t_SL _29596_ (.A(_07155_),
    .B(_07119_),
    .Y(_07156_));
 NAND2x1_ASAP7_75t_SL _29597_ (.A(_07138_),
    .B(_07156_),
    .Y(_07157_));
 AO21x1_ASAP7_75t_SL _29600_ (.A1(_07153_),
    .A2(_07157_),
    .B(_07146_),
    .Y(_07160_));
 OR2x2_ASAP7_75t_R _29601_ (.A(_00574_),
    .B(_00516_),
    .Y(_07161_));
 XOR2x2_ASAP7_75t_R _29602_ (.A(_00603_),
    .B(_00604_),
    .Y(_07162_));
 XOR2x2_ASAP7_75t_L _29603_ (.A(_12870_),
    .B(_00699_),
    .Y(_07163_));
 NOR2x1_ASAP7_75t_R _29604_ (.A(_07162_),
    .B(_07163_),
    .Y(_07164_));
 AND2x2_ASAP7_75t_R _29605_ (.A(_07163_),
    .B(_07162_),
    .Y(_07165_));
 OAI21x1_ASAP7_75t_R _29606_ (.A1(_07164_),
    .A2(_07165_),
    .B(_00574_),
    .Y(_07166_));
 NAND2x1_ASAP7_75t_R _29607_ (.A(_07161_),
    .B(_07166_),
    .Y(_07167_));
 XNOR2x2_ASAP7_75t_SL _29608_ (.A(_00961_),
    .B(_07167_),
    .Y(_07168_));
 AOI21x1_ASAP7_75t_SL _29611_ (.A1(_07150_),
    .A2(_07160_),
    .B(_07168_),
    .Y(_07171_));
 NOR2x1_ASAP7_75t_SL _29612_ (.A(_07094_),
    .B(_07081_),
    .Y(_07172_));
 OAI21x1_ASAP7_75t_SL _29613_ (.A1(_07112_),
    .A2(_07116_),
    .B(_07130_),
    .Y(_07173_));
 NOR2x1_ASAP7_75t_SL _29614_ (.A(_07172_),
    .B(_07173_),
    .Y(_07174_));
 NOR2x1_ASAP7_75t_SL _29615_ (.A(_07112_),
    .B(_07116_),
    .Y(_07175_));
 OAI21x1_ASAP7_75t_SL _29616_ (.A1(_07175_),
    .A2(_07172_),
    .B(_07138_),
    .Y(_07176_));
 NAND2x1_ASAP7_75t_SL _29617_ (.A(_07147_),
    .B(_07176_),
    .Y(_07177_));
 OAI21x1_ASAP7_75t_SL _29618_ (.A1(_07174_),
    .A2(_07177_),
    .B(_07168_),
    .Y(_07178_));
 OAI21x1_ASAP7_75t_SL _29619_ (.A1(_07067_),
    .A2(_07074_),
    .B(_08867_),
    .Y(_07179_));
 OAI21x1_ASAP7_75t_SL _29620_ (.A1(_07076_),
    .A2(_07079_),
    .B(_00945_),
    .Y(_07180_));
 NAND2x2_ASAP7_75t_SL _29621_ (.A(_07180_),
    .B(_07179_),
    .Y(_01384_));
 NOR2x2_ASAP7_75t_SL _29622_ (.A(_07119_),
    .B(_01384_),
    .Y(_07181_));
 NAND2x1_ASAP7_75t_SL _29623_ (.A(_07094_),
    .B(_07181_),
    .Y(_07182_));
 NOR2x1p5_ASAP7_75t_SL _29626_ (.A(_07155_),
    .B(_07112_),
    .Y(_07185_));
 NOR2x1_ASAP7_75t_SL _29627_ (.A(_07138_),
    .B(_07185_),
    .Y(_07186_));
 NOR2x1_ASAP7_75t_SL _29628_ (.A(_07122_),
    .B(_07119_),
    .Y(_07187_));
 NOR2x1_ASAP7_75t_SL _29629_ (.A(_07134_),
    .B(_07112_),
    .Y(_07188_));
 OA21x2_ASAP7_75t_SL _29631_ (.A1(_07187_),
    .A2(_07188_),
    .B(_07138_),
    .Y(_07190_));
 AOI211x1_ASAP7_75t_SL _29632_ (.A1(_07182_),
    .A2(_07186_),
    .B(_07190_),
    .C(_07147_),
    .Y(_07191_));
 XOR2x2_ASAP7_75t_R _29633_ (.A(_00604_),
    .B(_00605_),
    .Y(_07192_));
 XOR2x2_ASAP7_75t_R _29634_ (.A(_07192_),
    .B(_01713_),
    .Y(_07193_));
 XOR2x2_ASAP7_75t_R _29635_ (.A(_07193_),
    .B(_12906_),
    .Y(_07194_));
 NOR2x1_ASAP7_75t_R _29636_ (.A(_00574_),
    .B(_00508_),
    .Y(_07195_));
 AO21x1_ASAP7_75t_R _29637_ (.A1(_07194_),
    .A2(_00574_),
    .B(_07195_),
    .Y(_07196_));
 XNOR2x2_ASAP7_75t_SL _29638_ (.A(_00962_),
    .B(_07196_),
    .Y(_07197_));
 INVx2_ASAP7_75t_SL _29639_ (.A(_07197_),
    .Y(_07198_));
 OAI21x1_ASAP7_75t_SL _29641_ (.A1(_07178_),
    .A2(_07191_),
    .B(_07198_),
    .Y(_07200_));
 NOR2x1_ASAP7_75t_SL _29642_ (.A(_07171_),
    .B(_07200_),
    .Y(_07201_));
 NAND2x2_ASAP7_75t_L _29643_ (.A(_07112_),
    .B(_01384_),
    .Y(_07202_));
 AO21x1_ASAP7_75t_R _29644_ (.A1(_07118_),
    .A2(_07117_),
    .B(_01387_),
    .Y(_07203_));
 AO21x1_ASAP7_75t_SL _29646_ (.A1(_07202_),
    .A2(_07203_),
    .B(_07138_),
    .Y(_07205_));
 AOI21x1_ASAP7_75t_SL _29647_ (.A1(_07112_),
    .A2(_07116_),
    .B(_07130_),
    .Y(_07206_));
 NOR2x2_ASAP7_75t_SL _29648_ (.A(_07112_),
    .B(_01384_),
    .Y(_07207_));
 NAND2x1_ASAP7_75t_SL _29649_ (.A(_07094_),
    .B(_07207_),
    .Y(_07208_));
 NAND2x1_ASAP7_75t_SL _29650_ (.A(_07206_),
    .B(_07208_),
    .Y(_07209_));
 AND2x2_ASAP7_75t_SL _29651_ (.A(_07209_),
    .B(_07146_),
    .Y(_07210_));
 NAND2x1_ASAP7_75t_SL _29653_ (.A(_01394_),
    .B(_07119_),
    .Y(_07212_));
 AO21x1_ASAP7_75t_SL _29655_ (.A1(_07206_),
    .A2(_07212_),
    .B(_07146_),
    .Y(_07214_));
 NOR2x1_ASAP7_75t_SL _29656_ (.A(_07112_),
    .B(_07081_),
    .Y(_07215_));
 OAI21x1_ASAP7_75t_SL _29658_ (.A1(_07094_),
    .A2(_07152_),
    .B(_07130_),
    .Y(_07217_));
 NOR2x1_ASAP7_75t_SL _29659_ (.A(_07215_),
    .B(_07217_),
    .Y(_07218_));
 INVx1_ASAP7_75t_SL _29660_ (.A(_07168_),
    .Y(_07219_));
 OAI21x1_ASAP7_75t_SL _29663_ (.A1(_07214_),
    .A2(_07218_),
    .B(_07219_),
    .Y(_07222_));
 AOI21x1_ASAP7_75t_SL _29664_ (.A1(_07205_),
    .A2(_07210_),
    .B(_07222_),
    .Y(_07223_));
 NOR2x1_ASAP7_75t_SL _29666_ (.A(_07119_),
    .B(_07094_),
    .Y(_07225_));
 NOR2x1_ASAP7_75t_SL _29667_ (.A(_07138_),
    .B(_07225_),
    .Y(_07226_));
 NOR2x1_ASAP7_75t_SL _29668_ (.A(_07147_),
    .B(_07226_),
    .Y(_07227_));
 AOI21x1_ASAP7_75t_SL _29670_ (.A1(_01389_),
    .A2(_07119_),
    .B(_07130_),
    .Y(_07229_));
 NAND2x1_ASAP7_75t_SL _29671_ (.A(_07116_),
    .B(_07181_),
    .Y(_07230_));
 NAND2x1_ASAP7_75t_SL _29672_ (.A(_07229_),
    .B(_07230_),
    .Y(_07231_));
 AO21x1_ASAP7_75t_SL _29674_ (.A1(_07227_),
    .A2(_07231_),
    .B(_07219_),
    .Y(_07233_));
 AOI21x1_ASAP7_75t_SL _29675_ (.A1(_07116_),
    .A2(_07081_),
    .B(_07119_),
    .Y(_07234_));
 OAI21x1_ASAP7_75t_SL _29677_ (.A1(_07175_),
    .A2(_07234_),
    .B(_07130_),
    .Y(_07236_));
 AO21x2_ASAP7_75t_SL _29678_ (.A1(_07118_),
    .A2(_07117_),
    .B(_07155_),
    .Y(_07237_));
 AOI21x1_ASAP7_75t_R _29681_ (.A1(_01394_),
    .A2(_07112_),
    .B(_07130_),
    .Y(_07240_));
 NAND2x1_ASAP7_75t_SL _29682_ (.A(_07237_),
    .B(_07240_),
    .Y(_07241_));
 AND3x1_ASAP7_75t_SL _29683_ (.A(_07236_),
    .B(_07147_),
    .C(_07241_),
    .Y(_07242_));
 OAI21x1_ASAP7_75t_SL _29685_ (.A1(_07233_),
    .A2(_07242_),
    .B(_07197_),
    .Y(_07244_));
 XOR2x2_ASAP7_75t_SL _29686_ (.A(_00605_),
    .B(_00606_),
    .Y(_07245_));
 XOR2x2_ASAP7_75t_R _29687_ (.A(_07245_),
    .B(_00701_),
    .Y(_07246_));
 XOR2x2_ASAP7_75t_SL _29688_ (.A(_07246_),
    .B(_12914_),
    .Y(_07247_));
 NOR2x1_ASAP7_75t_SL _29689_ (.A(_00574_),
    .B(_00500_),
    .Y(_07248_));
 AO21x1_ASAP7_75t_SL _29690_ (.A1(_07247_),
    .A2(_00574_),
    .B(_07248_),
    .Y(_07249_));
 XOR2x2_ASAP7_75t_SL _29691_ (.A(_07249_),
    .B(_00963_),
    .Y(_07250_));
 OAI21x1_ASAP7_75t_SL _29693_ (.A1(_07223_),
    .A2(_07244_),
    .B(_07250_),
    .Y(_07252_));
 NOR2x1_ASAP7_75t_SL _29694_ (.A(_01389_),
    .B(_07119_),
    .Y(_07253_));
 AOI21x1_ASAP7_75t_SL _29695_ (.A1(_07116_),
    .A2(_07081_),
    .B(_07112_),
    .Y(_07254_));
 OAI21x1_ASAP7_75t_SL _29696_ (.A1(_07253_),
    .A2(_07254_),
    .B(_07130_),
    .Y(_07255_));
 NAND2x2_ASAP7_75t_SL _29697_ (.A(_07112_),
    .B(_07094_),
    .Y(_07256_));
 AO21x1_ASAP7_75t_SL _29698_ (.A1(_07256_),
    .A2(_07136_),
    .B(_07130_),
    .Y(_07257_));
 AO21x1_ASAP7_75t_SL _29699_ (.A1(_07111_),
    .A2(_07108_),
    .B(_01387_),
    .Y(_07258_));
 OA21x2_ASAP7_75t_SL _29700_ (.A1(_07258_),
    .A2(_07138_),
    .B(_07146_),
    .Y(_07259_));
 AND2x2_ASAP7_75t_SL _29701_ (.A(_07257_),
    .B(_07259_),
    .Y(_07260_));
 AO21x1_ASAP7_75t_SL _29702_ (.A1(_07111_),
    .A2(_07108_),
    .B(_01386_),
    .Y(_07261_));
 AND2x2_ASAP7_75t_SL _29704_ (.A(_07138_),
    .B(_01399_),
    .Y(_07263_));
 AO21x1_ASAP7_75t_SL _29705_ (.A1(_07130_),
    .A2(_07261_),
    .B(_07263_),
    .Y(_07264_));
 AO21x1_ASAP7_75t_SL _29707_ (.A1(_07264_),
    .A2(_07147_),
    .B(_07168_),
    .Y(_07266_));
 AOI21x1_ASAP7_75t_SL _29708_ (.A1(_07255_),
    .A2(_07260_),
    .B(_07266_),
    .Y(_07267_));
 NAND2x1_ASAP7_75t_SL _29709_ (.A(_07116_),
    .B(_07207_),
    .Y(_07268_));
 AOI21x1_ASAP7_75t_SL _29710_ (.A1(_07134_),
    .A2(_07112_),
    .B(_07138_),
    .Y(_07269_));
 NOR2x1_ASAP7_75t_SL _29711_ (.A(_01387_),
    .B(_07112_),
    .Y(_07270_));
 AO21x1_ASAP7_75t_SL _29712_ (.A1(_07270_),
    .A2(_07138_),
    .B(_07146_),
    .Y(_07271_));
 AO21x1_ASAP7_75t_SL _29713_ (.A1(_07268_),
    .A2(_07269_),
    .B(_07271_),
    .Y(_07272_));
 OA21x2_ASAP7_75t_SL _29714_ (.A1(_07203_),
    .A2(_07138_),
    .B(_07146_),
    .Y(_07273_));
 AOI21x1_ASAP7_75t_SL _29715_ (.A1(_01392_),
    .A2(_07112_),
    .B(_07130_),
    .Y(_07274_));
 NAND2x1_ASAP7_75t_SL _29716_ (.A(_07274_),
    .B(_07268_),
    .Y(_07275_));
 AOI21x1_ASAP7_75t_SL _29717_ (.A1(_07273_),
    .A2(_07275_),
    .B(_07219_),
    .Y(_07276_));
 AO21x1_ASAP7_75t_SL _29718_ (.A1(_07272_),
    .A2(_07276_),
    .B(_07197_),
    .Y(_07277_));
 NAND2x1_ASAP7_75t_SL _29719_ (.A(_07119_),
    .B(_07116_),
    .Y(_07278_));
 INVx1_ASAP7_75t_L _29720_ (.A(_07278_),
    .Y(_07279_));
 AO21x1_ASAP7_75t_SL _29721_ (.A1(_07112_),
    .A2(_07134_),
    .B(_07130_),
    .Y(_07280_));
 NOR2x1_ASAP7_75t_SL _29722_ (.A(_07279_),
    .B(_07280_),
    .Y(_07281_));
 AOI21x1_ASAP7_75t_SL _29723_ (.A1(_07119_),
    .A2(_07081_),
    .B(_07138_),
    .Y(_07282_));
 AO21x1_ASAP7_75t_SL _29725_ (.A1(_07282_),
    .A2(_07261_),
    .B(_07147_),
    .Y(_07284_));
 OAI21x1_ASAP7_75t_SL _29726_ (.A1(_07187_),
    .A2(_07270_),
    .B(_07130_),
    .Y(_07285_));
 NOR2x1_ASAP7_75t_SL _29727_ (.A(_07146_),
    .B(_07229_),
    .Y(_07286_));
 AOI21x1_ASAP7_75t_SL _29728_ (.A1(_07285_),
    .A2(_07286_),
    .B(_07219_),
    .Y(_07287_));
 OAI21x1_ASAP7_75t_SL _29729_ (.A1(_07281_),
    .A2(_07284_),
    .B(_07287_),
    .Y(_07288_));
 AOI21x1_ASAP7_75t_SL _29730_ (.A1(_07138_),
    .A2(_07237_),
    .B(_07146_),
    .Y(_07289_));
 AO21x1_ASAP7_75t_R _29731_ (.A1(_07118_),
    .A2(_07117_),
    .B(_01392_),
    .Y(_07290_));
 INVx1_ASAP7_75t_SL _29733_ (.A(_07290_),
    .Y(_07292_));
 OAI21x1_ASAP7_75t_SL _29734_ (.A1(_07253_),
    .A2(_07292_),
    .B(_07130_),
    .Y(_07293_));
 AOI21x1_ASAP7_75t_SL _29735_ (.A1(_07289_),
    .A2(_07293_),
    .B(_07168_),
    .Y(_07294_));
 AO21x2_ASAP7_75t_L _29737_ (.A1(_07111_),
    .A2(_07108_),
    .B(_01389_),
    .Y(_07296_));
 NOR2x1_ASAP7_75t_L _29738_ (.A(_07138_),
    .B(_07296_),
    .Y(_07297_));
 NOR2x1_ASAP7_75t_SL _29739_ (.A(_07147_),
    .B(_07297_),
    .Y(_07298_));
 NAND2x1_ASAP7_75t_SL _29740_ (.A(_07298_),
    .B(_07209_),
    .Y(_07299_));
 AOI21x1_ASAP7_75t_SL _29741_ (.A1(_07294_),
    .A2(_07299_),
    .B(_07198_),
    .Y(_07300_));
 AOI21x1_ASAP7_75t_SL _29742_ (.A1(_07288_),
    .A2(_07300_),
    .B(_07250_),
    .Y(_07301_));
 OAI21x1_ASAP7_75t_SL _29743_ (.A1(_07267_),
    .A2(_07277_),
    .B(_07301_),
    .Y(_07302_));
 OAI21x1_ASAP7_75t_SL _29744_ (.A1(_07201_),
    .A2(_07252_),
    .B(_07302_),
    .Y(_00152_));
 AOI21x1_ASAP7_75t_R _29745_ (.A1(_07094_),
    .A2(_07081_),
    .B(_07112_),
    .Y(_07303_));
 NAND2x1_ASAP7_75t_SL _29746_ (.A(_07130_),
    .B(_07303_),
    .Y(_07304_));
 NAND2x1_ASAP7_75t_SL _29747_ (.A(_07119_),
    .B(_01384_),
    .Y(_07305_));
 AOI21x1_ASAP7_75t_SL _29748_ (.A1(_07305_),
    .A2(_07240_),
    .B(_07146_),
    .Y(_07306_));
 AO21x1_ASAP7_75t_R _29749_ (.A1(_07118_),
    .A2(_07117_),
    .B(_01389_),
    .Y(_07307_));
 OA21x2_ASAP7_75t_SL _29750_ (.A1(_07307_),
    .A2(_07138_),
    .B(_07146_),
    .Y(_07308_));
 AOI21x1_ASAP7_75t_SL _29751_ (.A1(_07094_),
    .A2(_07081_),
    .B(_07119_),
    .Y(_07309_));
 OAI21x1_ASAP7_75t_SL _29753_ (.A1(_07185_),
    .A2(_07309_),
    .B(_07138_),
    .Y(_07311_));
 AOI221x1_ASAP7_75t_SL _29754_ (.A1(_07304_),
    .A2(_07306_),
    .B1(_07308_),
    .B2(_07311_),
    .C(_07219_),
    .Y(_07312_));
 AO21x1_ASAP7_75t_SL _29755_ (.A1(_07256_),
    .A2(_07136_),
    .B(_07138_),
    .Y(_07313_));
 AO21x1_ASAP7_75t_SL _29756_ (.A1(_07237_),
    .A2(_07296_),
    .B(_07130_),
    .Y(_07314_));
 AO21x1_ASAP7_75t_SL _29757_ (.A1(_07314_),
    .A2(_07313_),
    .B(_07146_),
    .Y(_07315_));
 NAND2x1_ASAP7_75t_SL _29758_ (.A(_07094_),
    .B(_07081_),
    .Y(_07316_));
 AO21x1_ASAP7_75t_SL _29759_ (.A1(_07316_),
    .A2(_07278_),
    .B(_07130_),
    .Y(_07317_));
 NOR2x1_ASAP7_75t_SL _29760_ (.A(_01386_),
    .B(_07119_),
    .Y(_07318_));
 NOR2x1_ASAP7_75t_SL _29761_ (.A(_07138_),
    .B(_07318_),
    .Y(_07319_));
 NAND2x1_ASAP7_75t_SL _29762_ (.A(_07278_),
    .B(_07319_),
    .Y(_07320_));
 AO21x1_ASAP7_75t_SL _29763_ (.A1(_07317_),
    .A2(_07320_),
    .B(_07147_),
    .Y(_07321_));
 AOI21x1_ASAP7_75t_SL _29764_ (.A1(_07315_),
    .A2(_07321_),
    .B(_07168_),
    .Y(_07322_));
 OAI21x1_ASAP7_75t_SL _29765_ (.A1(_07322_),
    .A2(_07312_),
    .B(_07197_),
    .Y(_07323_));
 AO21x1_ASAP7_75t_R _29766_ (.A1(_07081_),
    .A2(_07112_),
    .B(_07130_),
    .Y(_07324_));
 AND3x1_ASAP7_75t_SL _29767_ (.A(_07324_),
    .B(_07147_),
    .C(_07305_),
    .Y(_07325_));
 AO21x1_ASAP7_75t_SL _29768_ (.A1(_07118_),
    .A2(_07117_),
    .B(_01394_),
    .Y(_07326_));
 AO21x1_ASAP7_75t_SL _29769_ (.A1(_07261_),
    .A2(_07326_),
    .B(_07130_),
    .Y(_07327_));
 NAND2x1_ASAP7_75t_SL _29770_ (.A(_07130_),
    .B(_07254_),
    .Y(_07328_));
 AND3x1_ASAP7_75t_SL _29771_ (.A(_07327_),
    .B(_07146_),
    .C(_07328_),
    .Y(_07329_));
 NOR2x1_ASAP7_75t_SL _29772_ (.A(_07168_),
    .B(_07297_),
    .Y(_07330_));
 OAI21x1_ASAP7_75t_SL _29773_ (.A1(_07325_),
    .A2(_07329_),
    .B(_07330_),
    .Y(_07331_));
 NAND2x1_ASAP7_75t_R _29774_ (.A(_07112_),
    .B(_07116_),
    .Y(_07332_));
 AOI21x1_ASAP7_75t_SL _29775_ (.A1(_07307_),
    .A2(_07332_),
    .B(_07138_),
    .Y(_07333_));
 AO21x1_ASAP7_75t_SL _29777_ (.A1(_07206_),
    .A2(_07237_),
    .B(_07146_),
    .Y(_07335_));
 NOR2x1_ASAP7_75t_SL _29778_ (.A(_07119_),
    .B(_07130_),
    .Y(_07336_));
 NAND2x1_ASAP7_75t_R _29779_ (.A(_07116_),
    .B(_07081_),
    .Y(_07337_));
 NAND2x1_ASAP7_75t_SL _29780_ (.A(_07336_),
    .B(_07337_),
    .Y(_07338_));
 INVx1_ASAP7_75t_SL _29781_ (.A(_07172_),
    .Y(_07339_));
 AOI21x1_ASAP7_75t_SL _29782_ (.A1(_07282_),
    .A2(_07339_),
    .B(_07147_),
    .Y(_07340_));
 NAND2x1_ASAP7_75t_SL _29783_ (.A(_07338_),
    .B(_07340_),
    .Y(_07341_));
 OAI21x1_ASAP7_75t_SL _29784_ (.A1(_07333_),
    .A2(_07335_),
    .B(_07341_),
    .Y(_07342_));
 AOI21x1_ASAP7_75t_SL _29785_ (.A1(_07168_),
    .A2(_07342_),
    .B(_07197_),
    .Y(_07343_));
 AOI21x1_ASAP7_75t_SL _29786_ (.A1(_07331_),
    .A2(_07343_),
    .B(_07250_),
    .Y(_07344_));
 NOR2x1_ASAP7_75t_SL _29787_ (.A(_07130_),
    .B(_07168_),
    .Y(_07345_));
 AOI21x1_ASAP7_75t_SL _29788_ (.A1(_01401_),
    .A2(_07345_),
    .B(_07197_),
    .Y(_07346_));
 NAND2x1_ASAP7_75t_SL _29789_ (.A(_07269_),
    .B(_07208_),
    .Y(_07347_));
 AO21x1_ASAP7_75t_SL _29790_ (.A1(_07346_),
    .A2(_07347_),
    .B(_07147_),
    .Y(_07348_));
 AO21x1_ASAP7_75t_SL _29791_ (.A1(_07116_),
    .A2(_07112_),
    .B(_07138_),
    .Y(_07349_));
 INVx1_ASAP7_75t_SL _29792_ (.A(_07208_),
    .Y(_07350_));
 AOI21x1_ASAP7_75t_SL _29793_ (.A1(_07138_),
    .A2(_07237_),
    .B(_07168_),
    .Y(_07351_));
 OAI21x1_ASAP7_75t_SL _29794_ (.A1(_07349_),
    .A2(_07350_),
    .B(_07351_),
    .Y(_07352_));
 AOI21x1_ASAP7_75t_SL _29795_ (.A1(_07202_),
    .A2(_07229_),
    .B(_07219_),
    .Y(_07353_));
 AO21x1_ASAP7_75t_SL _29797_ (.A1(_07278_),
    .A2(_07123_),
    .B(_07138_),
    .Y(_07355_));
 NAND2x1_ASAP7_75t_SL _29798_ (.A(_07353_),
    .B(_07355_),
    .Y(_07356_));
 AOI21x1_ASAP7_75t_SL _29799_ (.A1(_07352_),
    .A2(_07356_),
    .B(_07198_),
    .Y(_07357_));
 OAI21x1_ASAP7_75t_SL _29800_ (.A1(_07348_),
    .A2(_07357_),
    .B(_07250_),
    .Y(_07358_));
 INVx1_ASAP7_75t_SL _29801_ (.A(_01387_),
    .Y(_07359_));
 AO21x1_ASAP7_75t_SL _29802_ (.A1(_07111_),
    .A2(_07108_),
    .B(_07359_),
    .Y(_07360_));
 AOI21x1_ASAP7_75t_SL _29803_ (.A1(_01394_),
    .A2(_07119_),
    .B(_07138_),
    .Y(_07361_));
 AOI21x1_ASAP7_75t_SL _29804_ (.A1(_07360_),
    .A2(_07361_),
    .B(_07168_),
    .Y(_07362_));
 AOI21x1_ASAP7_75t_SL _29805_ (.A1(_07362_),
    .A2(_07311_),
    .B(_07198_),
    .Y(_07363_));
 AOI21x1_ASAP7_75t_SL _29806_ (.A1(_07130_),
    .A2(_07270_),
    .B(_07219_),
    .Y(_07364_));
 NOR2x1_ASAP7_75t_SL _29807_ (.A(_07122_),
    .B(_07112_),
    .Y(_07365_));
 OAI21x1_ASAP7_75t_SL _29808_ (.A1(_07365_),
    .A2(_07318_),
    .B(_07138_),
    .Y(_07366_));
 OR3x1_ASAP7_75t_SL _29809_ (.A(_07116_),
    .B(_07119_),
    .C(_07138_),
    .Y(_07367_));
 NAND3x1_ASAP7_75t_SL _29810_ (.A(_07364_),
    .B(_07366_),
    .C(_07367_),
    .Y(_07368_));
 NAND2x1_ASAP7_75t_SL _29811_ (.A(_07363_),
    .B(_07368_),
    .Y(_07369_));
 NAND2x1_ASAP7_75t_SL _29812_ (.A(_07202_),
    .B(_07229_),
    .Y(_07370_));
 OA21x2_ASAP7_75t_SL _29813_ (.A1(_07173_),
    .A2(_07181_),
    .B(_07219_),
    .Y(_07371_));
 NAND2x1_ASAP7_75t_SL _29814_ (.A(_07370_),
    .B(_07371_),
    .Y(_07372_));
 AOI21x1_ASAP7_75t_SL _29815_ (.A1(_07122_),
    .A2(_07112_),
    .B(_07138_),
    .Y(_07373_));
 AOI21x1_ASAP7_75t_SL _29816_ (.A1(_07278_),
    .A2(_07373_),
    .B(_07219_),
    .Y(_07374_));
 OAI21x1_ASAP7_75t_SL _29817_ (.A1(_07303_),
    .A2(_07234_),
    .B(_07138_),
    .Y(_07375_));
 AOI21x1_ASAP7_75t_SL _29819_ (.A1(_07374_),
    .A2(_07375_),
    .B(_07197_),
    .Y(_07377_));
 NAND2x1_ASAP7_75t_SL _29820_ (.A(_07372_),
    .B(_07377_),
    .Y(_07378_));
 AOI21x1_ASAP7_75t_SL _29821_ (.A1(_07369_),
    .A2(_07378_),
    .B(_07146_),
    .Y(_07379_));
 NOR2x1_ASAP7_75t_SL _29822_ (.A(_07358_),
    .B(_07379_),
    .Y(_07380_));
 AOI21x1_ASAP7_75t_SL _29823_ (.A1(_07323_),
    .A2(_07344_),
    .B(_07380_),
    .Y(_00153_));
 NAND2x1_ASAP7_75t_SL _29824_ (.A(_01398_),
    .B(_07138_),
    .Y(_07381_));
 AO21x1_ASAP7_75t_R _29825_ (.A1(_07217_),
    .A2(_07381_),
    .B(_07147_),
    .Y(_07382_));
 NOR2x1_ASAP7_75t_SL _29826_ (.A(_07130_),
    .B(_07207_),
    .Y(_07383_));
 NAND2x1_ASAP7_75t_R _29827_ (.A(_07337_),
    .B(_07383_),
    .Y(_07384_));
 OR2x2_ASAP7_75t_R _29828_ (.A(_07138_),
    .B(_01403_),
    .Y(_07385_));
 AO21x1_ASAP7_75t_R _29829_ (.A1(_07384_),
    .A2(_07385_),
    .B(_07146_),
    .Y(_07386_));
 AOI21x1_ASAP7_75t_R _29830_ (.A1(_07382_),
    .A2(_07386_),
    .B(_07197_),
    .Y(_07387_));
 INVx1_ASAP7_75t_R _29831_ (.A(_01401_),
    .Y(_07388_));
 AOI21x1_ASAP7_75t_SL _29832_ (.A1(_07339_),
    .A2(_07383_),
    .B(_07147_),
    .Y(_07389_));
 OA21x2_ASAP7_75t_R _29833_ (.A1(_07388_),
    .A2(_07138_),
    .B(_07389_),
    .Y(_07390_));
 NOR2x1_ASAP7_75t_SL _29834_ (.A(_07130_),
    .B(_07188_),
    .Y(_07391_));
 AOI22x1_ASAP7_75t_R _29835_ (.A1(_07123_),
    .A2(_07282_),
    .B1(_07391_),
    .B2(_07261_),
    .Y(_07392_));
 OAI21x1_ASAP7_75t_R _29836_ (.A1(_07146_),
    .A2(_07392_),
    .B(_07197_),
    .Y(_07393_));
 INVx1_ASAP7_75t_SL _29837_ (.A(_07250_),
    .Y(_07394_));
 OAI21x1_ASAP7_75t_R _29838_ (.A1(_07390_),
    .A2(_07393_),
    .B(_07394_),
    .Y(_07395_));
 NOR2x1_ASAP7_75t_SL _29839_ (.A(_07387_),
    .B(_07395_),
    .Y(_07396_));
 OAI21x1_ASAP7_75t_R _29840_ (.A1(_07253_),
    .A2(_07254_),
    .B(_07138_),
    .Y(_07397_));
 NAND2x1_ASAP7_75t_SL _29841_ (.A(_07119_),
    .B(_07081_),
    .Y(_07398_));
 AO21x1_ASAP7_75t_SL _29842_ (.A1(_07398_),
    .A2(_07261_),
    .B(_07138_),
    .Y(_07399_));
 AOI21x1_ASAP7_75t_R _29843_ (.A1(_07397_),
    .A2(_07399_),
    .B(_07147_),
    .Y(_07400_));
 AOI21x1_ASAP7_75t_SL _29844_ (.A1(_01389_),
    .A2(_07119_),
    .B(_07138_),
    .Y(_07401_));
 AOI21x1_ASAP7_75t_R _29845_ (.A1(_01394_),
    .A2(_07112_),
    .B(_07146_),
    .Y(_07402_));
 AOI21x1_ASAP7_75t_SL _29846_ (.A1(_07401_),
    .A2(_07402_),
    .B(_07197_),
    .Y(_07403_));
 OAI21x1_ASAP7_75t_R _29847_ (.A1(_07146_),
    .A2(_07384_),
    .B(_07403_),
    .Y(_07404_));
 NOR2x1_ASAP7_75t_SL _29848_ (.A(_07400_),
    .B(_07404_),
    .Y(_07405_));
 AO21x2_ASAP7_75t_SL _29849_ (.A1(_07111_),
    .A2(_07108_),
    .B(_01394_),
    .Y(_07406_));
 AND2x2_ASAP7_75t_SL _29850_ (.A(_07406_),
    .B(_07130_),
    .Y(_07407_));
 OAI21x1_ASAP7_75t_SL _29851_ (.A1(_07112_),
    .A2(_07116_),
    .B(_07138_),
    .Y(_07408_));
 NOR2x1_ASAP7_75t_SL _29852_ (.A(_07253_),
    .B(_07408_),
    .Y(_07409_));
 NOR2x1_ASAP7_75t_SL _29854_ (.A(_07138_),
    .B(_07290_),
    .Y(_07411_));
 NOR2x1_ASAP7_75t_R _29855_ (.A(_07146_),
    .B(_07411_),
    .Y(_07412_));
 OAI21x1_ASAP7_75t_R _29856_ (.A1(_07407_),
    .A2(_07409_),
    .B(_07412_),
    .Y(_07413_));
 AO21x1_ASAP7_75t_R _29857_ (.A1(_07398_),
    .A2(_07296_),
    .B(_07130_),
    .Y(_07414_));
 NAND2x1_ASAP7_75t_SL _29858_ (.A(_07296_),
    .B(_07290_),
    .Y(_07415_));
 AOI21x1_ASAP7_75t_R _29859_ (.A1(_07130_),
    .A2(_07415_),
    .B(_07147_),
    .Y(_07416_));
 NAND2x1_ASAP7_75t_R _29860_ (.A(_07414_),
    .B(_07416_),
    .Y(_07417_));
 AOI21x1_ASAP7_75t_R _29861_ (.A1(_07413_),
    .A2(_07417_),
    .B(_07198_),
    .Y(_07418_));
 NOR2x1_ASAP7_75t_SL _29862_ (.A(_07405_),
    .B(_07418_),
    .Y(_07419_));
 OAI21x1_ASAP7_75t_R _29863_ (.A1(_07394_),
    .A2(_07419_),
    .B(_07219_),
    .Y(_07420_));
 INVx1_ASAP7_75t_R _29864_ (.A(_07326_),
    .Y(_07421_));
 OAI21x1_ASAP7_75t_R _29865_ (.A1(_07421_),
    .A2(_07309_),
    .B(_07138_),
    .Y(_07422_));
 AOI21x1_ASAP7_75t_R _29866_ (.A1(_07217_),
    .A2(_07422_),
    .B(_07147_),
    .Y(_07423_));
 INVx1_ASAP7_75t_R _29867_ (.A(_07258_),
    .Y(_07424_));
 OAI21x1_ASAP7_75t_R _29868_ (.A1(_07424_),
    .A2(_07408_),
    .B(_07147_),
    .Y(_07425_));
 AND3x1_ASAP7_75t_R _29870_ (.A(_07202_),
    .B(_07130_),
    .C(_07121_),
    .Y(_07427_));
 OAI21x1_ASAP7_75t_R _29871_ (.A1(_07425_),
    .A2(_07427_),
    .B(_07198_),
    .Y(_07428_));
 NOR2x1_ASAP7_75t_L _29872_ (.A(_07423_),
    .B(_07428_),
    .Y(_07429_));
 AOI21x1_ASAP7_75t_SL _29873_ (.A1(_01392_),
    .A2(_07112_),
    .B(_07138_),
    .Y(_07430_));
 NAND2x1_ASAP7_75t_SL _29874_ (.A(_07278_),
    .B(_07430_),
    .Y(_07431_));
 AO21x2_ASAP7_75t_SL _29875_ (.A1(_07111_),
    .A2(_07108_),
    .B(_07155_),
    .Y(_07432_));
 AO21x1_ASAP7_75t_SL _29876_ (.A1(_07432_),
    .A2(_07121_),
    .B(_07130_),
    .Y(_07433_));
 AOI21x1_ASAP7_75t_R _29877_ (.A1(_07431_),
    .A2(_07433_),
    .B(_07147_),
    .Y(_07434_));
 INVx1_ASAP7_75t_R _29878_ (.A(_07406_),
    .Y(_07435_));
 OAI21x1_ASAP7_75t_SL _29879_ (.A1(_07435_),
    .A2(_07173_),
    .B(_07147_),
    .Y(_07436_));
 AND3x1_ASAP7_75t_R _29880_ (.A(_07202_),
    .B(_07138_),
    .C(_07290_),
    .Y(_07437_));
 OAI21x1_ASAP7_75t_R _29881_ (.A1(_07436_),
    .A2(_07437_),
    .B(_07197_),
    .Y(_07438_));
 NOR2x1_ASAP7_75t_SL _29882_ (.A(_07434_),
    .B(_07438_),
    .Y(_07439_));
 OAI21x1_ASAP7_75t_SL _29883_ (.A1(_07439_),
    .A2(_07429_),
    .B(_07250_),
    .Y(_07440_));
 AOI21x1_ASAP7_75t_R _29884_ (.A1(_07261_),
    .A2(_07282_),
    .B(_07146_),
    .Y(_07441_));
 NAND2x1_ASAP7_75t_SL _29885_ (.A(_07119_),
    .B(_07094_),
    .Y(_07442_));
 AO21x1_ASAP7_75t_SL _29886_ (.A1(_07152_),
    .A2(_07442_),
    .B(_07130_),
    .Y(_07443_));
 NAND2x1_ASAP7_75t_R _29887_ (.A(_07441_),
    .B(_07443_),
    .Y(_07444_));
 OA21x2_ASAP7_75t_R _29888_ (.A1(_01399_),
    .A2(_07138_),
    .B(_07146_),
    .Y(_07445_));
 OAI21x1_ASAP7_75t_SL _29889_ (.A1(_07318_),
    .A2(_07254_),
    .B(_07138_),
    .Y(_07446_));
 AOI21x1_ASAP7_75t_R _29890_ (.A1(_07445_),
    .A2(_07446_),
    .B(_07198_),
    .Y(_07447_));
 NAND2x1_ASAP7_75t_L _29891_ (.A(_07444_),
    .B(_07447_),
    .Y(_07448_));
 AO21x1_ASAP7_75t_SL _29892_ (.A1(_07296_),
    .A2(_07121_),
    .B(_07130_),
    .Y(_07449_));
 NOR2x1_ASAP7_75t_SL _29893_ (.A(_07138_),
    .B(_07136_),
    .Y(_07450_));
 NOR2x1_ASAP7_75t_R _29894_ (.A(_07147_),
    .B(_07450_),
    .Y(_07451_));
 AOI21x1_ASAP7_75t_R _29895_ (.A1(_07449_),
    .A2(_07451_),
    .B(_07197_),
    .Y(_07452_));
 AND2x2_ASAP7_75t_R _29896_ (.A(_01387_),
    .B(_01389_),
    .Y(_07453_));
 NOR2x1_ASAP7_75t_L _29897_ (.A(_07453_),
    .B(_07112_),
    .Y(_07454_));
 OAI21x1_ASAP7_75t_R _29898_ (.A1(_07454_),
    .A2(_07309_),
    .B(_07138_),
    .Y(_07455_));
 AOI21x1_ASAP7_75t_R _29899_ (.A1(_07269_),
    .A2(_07208_),
    .B(_07146_),
    .Y(_07456_));
 NAND2x1_ASAP7_75t_R _29900_ (.A(_07455_),
    .B(_07456_),
    .Y(_07457_));
 AOI21x1_ASAP7_75t_R _29901_ (.A1(_07452_),
    .A2(_07457_),
    .B(_07250_),
    .Y(_07458_));
 AOI21x1_ASAP7_75t_R _29902_ (.A1(_07448_),
    .A2(_07458_),
    .B(_07219_),
    .Y(_07459_));
 NAND2x1_ASAP7_75t_SL _29903_ (.A(_07440_),
    .B(_07459_),
    .Y(_07460_));
 OAI21x1_ASAP7_75t_SL _29904_ (.A1(_07396_),
    .A2(_07420_),
    .B(_07460_),
    .Y(_00154_));
 NAND2x1_ASAP7_75t_SL _29905_ (.A(_07257_),
    .B(_07340_),
    .Y(_07461_));
 AO21x1_ASAP7_75t_R _29906_ (.A1(_07121_),
    .A2(_07406_),
    .B(_07138_),
    .Y(_07462_));
 NAND2x1_ASAP7_75t_SL _29907_ (.A(_07290_),
    .B(_07332_),
    .Y(_07463_));
 AOI21x1_ASAP7_75t_R _29908_ (.A1(_07138_),
    .A2(_07463_),
    .B(_07146_),
    .Y(_07464_));
 NAND2x1_ASAP7_75t_R _29909_ (.A(_07462_),
    .B(_07464_),
    .Y(_07465_));
 AOI21x1_ASAP7_75t_R _29910_ (.A1(_07461_),
    .A2(_07465_),
    .B(_07219_),
    .Y(_07466_));
 NAND2x1_ASAP7_75t_SL _29911_ (.A(_07219_),
    .B(_07436_),
    .Y(_07467_));
 NAND2x1_ASAP7_75t_L _29912_ (.A(_07453_),
    .B(_07119_),
    .Y(_07468_));
 NAND2x1_ASAP7_75t_L _29913_ (.A(_07468_),
    .B(_07274_),
    .Y(_07469_));
 AOI21x1_ASAP7_75t_R _29914_ (.A1(_07469_),
    .A2(_07347_),
    .B(_07147_),
    .Y(_07470_));
 OAI21x1_ASAP7_75t_R _29915_ (.A1(_07467_),
    .A2(_07470_),
    .B(_07197_),
    .Y(_07471_));
 OAI21x1_ASAP7_75t_SL _29916_ (.A1(_07466_),
    .A2(_07471_),
    .B(_07250_),
    .Y(_07472_));
 NOR2x1_ASAP7_75t_SL _29917_ (.A(_07130_),
    .B(_07290_),
    .Y(_07473_));
 NOR2x1_ASAP7_75t_R _29918_ (.A(_07219_),
    .B(_07473_),
    .Y(_07474_));
 NAND2x1_ASAP7_75t_R _29919_ (.A(_07431_),
    .B(_07474_),
    .Y(_07475_));
 AO21x1_ASAP7_75t_SL _29920_ (.A1(_07256_),
    .A2(_07121_),
    .B(_07138_),
    .Y(_07476_));
 OAI21x1_ASAP7_75t_R _29921_ (.A1(_07454_),
    .A2(_07435_),
    .B(_07138_),
    .Y(_07477_));
 NAND3x1_ASAP7_75t_SL _29922_ (.A(_07476_),
    .B(_07219_),
    .C(_07477_),
    .Y(_07478_));
 AOI21x1_ASAP7_75t_R _29923_ (.A1(_07475_),
    .A2(_07478_),
    .B(_07147_),
    .Y(_07479_));
 NOR2x1_ASAP7_75t_SL _29924_ (.A(_07138_),
    .B(_07237_),
    .Y(_07480_));
 AOI21x1_ASAP7_75t_R _29925_ (.A1(_07168_),
    .A2(_07480_),
    .B(_07271_),
    .Y(_07481_));
 NAND2x1_ASAP7_75t_R _29926_ (.A(_07398_),
    .B(_07269_),
    .Y(_07482_));
 AO21x1_ASAP7_75t_SL _29927_ (.A1(_07482_),
    .A2(_07157_),
    .B(_07168_),
    .Y(_07483_));
 AO21x1_ASAP7_75t_R _29928_ (.A1(_07481_),
    .A2(_07483_),
    .B(_07197_),
    .Y(_07484_));
 NOR2x1_ASAP7_75t_R _29929_ (.A(_07479_),
    .B(_07484_),
    .Y(_07485_));
 NOR2x1_ASAP7_75t_SL _29930_ (.A(_07472_),
    .B(_07485_),
    .Y(_07486_));
 AND3x1_ASAP7_75t_R _29931_ (.A(_07136_),
    .B(_07432_),
    .C(_07138_),
    .Y(_07487_));
 AO21x1_ASAP7_75t_R _29932_ (.A1(_07118_),
    .A2(_07117_),
    .B(_07134_),
    .Y(_07488_));
 AND3x1_ASAP7_75t_SL _29933_ (.A(_07256_),
    .B(_07130_),
    .C(_07488_),
    .Y(_07489_));
 OAI21x1_ASAP7_75t_R _29934_ (.A1(_07487_),
    .A2(_07489_),
    .B(_07147_),
    .Y(_07490_));
 AO21x1_ASAP7_75t_R _29935_ (.A1(_07326_),
    .A2(_07296_),
    .B(_07130_),
    .Y(_07491_));
 NOR2x1_ASAP7_75t_SL _29936_ (.A(_01386_),
    .B(_07112_),
    .Y(_07492_));
 NOR2x1_ASAP7_75t_SL _29937_ (.A(_07138_),
    .B(_07492_),
    .Y(_07493_));
 AOI21x1_ASAP7_75t_R _29938_ (.A1(_07202_),
    .A2(_07493_),
    .B(_07147_),
    .Y(_07494_));
 AOI21x1_ASAP7_75t_R _29939_ (.A1(_07491_),
    .A2(_07494_),
    .B(_07219_),
    .Y(_07495_));
 NAND2x1_ASAP7_75t_R _29940_ (.A(_07490_),
    .B(_07495_),
    .Y(_07496_));
 AO21x1_ASAP7_75t_SL _29941_ (.A1(_07081_),
    .A2(_07116_),
    .B(_07173_),
    .Y(_07497_));
 NOR2x1_ASAP7_75t_SL _29942_ (.A(_07130_),
    .B(_07185_),
    .Y(_07498_));
 AOI21x1_ASAP7_75t_R _29943_ (.A1(_07202_),
    .A2(_07498_),
    .B(_07147_),
    .Y(_07499_));
 NAND2x1_ASAP7_75t_SL _29944_ (.A(_07497_),
    .B(_07499_),
    .Y(_07500_));
 OAI21x1_ASAP7_75t_R _29945_ (.A1(_07181_),
    .A2(_07173_),
    .B(_07157_),
    .Y(_07501_));
 AOI21x1_ASAP7_75t_R _29946_ (.A1(_07147_),
    .A2(_07501_),
    .B(_07168_),
    .Y(_07502_));
 AOI21x1_ASAP7_75t_SL _29947_ (.A1(_07500_),
    .A2(_07502_),
    .B(_07197_),
    .Y(_07503_));
 NAND2x1_ASAP7_75t_R _29948_ (.A(_07496_),
    .B(_07503_),
    .Y(_07504_));
 AO21x1_ASAP7_75t_R _29949_ (.A1(_07119_),
    .A2(_07138_),
    .B(_07147_),
    .Y(_07505_));
 AO21x1_ASAP7_75t_R _29950_ (.A1(_07442_),
    .A2(_07337_),
    .B(_07505_),
    .Y(_07506_));
 INVx1_ASAP7_75t_R _29951_ (.A(_01392_),
    .Y(_07507_));
 OAI21x1_ASAP7_75t_R _29952_ (.A1(_07507_),
    .A2(_07119_),
    .B(_07493_),
    .Y(_07508_));
 AOI21x1_ASAP7_75t_R _29953_ (.A1(_07306_),
    .A2(_07508_),
    .B(_07168_),
    .Y(_07509_));
 AOI21x1_ASAP7_75t_R _29954_ (.A1(_07506_),
    .A2(_07509_),
    .B(_07198_),
    .Y(_07510_));
 AND3x1_ASAP7_75t_R _29955_ (.A(_07237_),
    .B(_07135_),
    .C(_07130_),
    .Y(_07511_));
 NOR2x1_ASAP7_75t_L _29956_ (.A(_07511_),
    .B(_07177_),
    .Y(_07512_));
 INVx1_ASAP7_75t_SL _29957_ (.A(_07303_),
    .Y(_07513_));
 NAND2x1_ASAP7_75t_R _29958_ (.A(_07138_),
    .B(_07488_),
    .Y(_07514_));
 OAI21x1_ASAP7_75t_SL _29959_ (.A1(_07234_),
    .A2(_07514_),
    .B(_07146_),
    .Y(_07515_));
 AOI21x1_ASAP7_75t_R _29960_ (.A1(_07513_),
    .A2(_07319_),
    .B(_07515_),
    .Y(_07516_));
 OAI21x1_ASAP7_75t_SL _29961_ (.A1(_07512_),
    .A2(_07516_),
    .B(_07168_),
    .Y(_07517_));
 NAND2x1_ASAP7_75t_SL _29962_ (.A(_07510_),
    .B(_07517_),
    .Y(_07518_));
 AOI21x1_ASAP7_75t_SL _29963_ (.A1(_07504_),
    .A2(_07518_),
    .B(_07250_),
    .Y(_07519_));
 NOR2x1_ASAP7_75t_SL _29964_ (.A(_07486_),
    .B(_07519_),
    .Y(_00155_));
 NOR2x1_ASAP7_75t_R _29965_ (.A(_07147_),
    .B(_07336_),
    .Y(_07520_));
 AO21x1_ASAP7_75t_R _29966_ (.A1(_07278_),
    .A2(_07406_),
    .B(_07138_),
    .Y(_07521_));
 NAND2x1_ASAP7_75t_R _29967_ (.A(_07520_),
    .B(_07521_),
    .Y(_07522_));
 AOI21x1_ASAP7_75t_SL _29968_ (.A1(_07202_),
    .A2(_07229_),
    .B(_07146_),
    .Y(_07523_));
 AO21x1_ASAP7_75t_R _29969_ (.A1(_07202_),
    .A2(_07136_),
    .B(_07138_),
    .Y(_07524_));
 AOI21x1_ASAP7_75t_SL _29970_ (.A1(_07523_),
    .A2(_07524_),
    .B(_07168_),
    .Y(_07525_));
 NAND2x1_ASAP7_75t_SL _29971_ (.A(_07522_),
    .B(_07525_),
    .Y(_07526_));
 AOI21x1_ASAP7_75t_R _29972_ (.A1(_07261_),
    .A2(_07401_),
    .B(_07147_),
    .Y(_07527_));
 NAND2x1_ASAP7_75t_R _29973_ (.A(_07527_),
    .B(_07209_),
    .Y(_07528_));
 OA21x2_ASAP7_75t_SL _29974_ (.A1(_07119_),
    .A2(_07359_),
    .B(_07130_),
    .Y(_07529_));
 NOR2x1_ASAP7_75t_R _29975_ (.A(_07146_),
    .B(_07529_),
    .Y(_07530_));
 AO21x1_ASAP7_75t_R _29976_ (.A1(_07181_),
    .A2(_07094_),
    .B(_07130_),
    .Y(_07531_));
 AOI21x1_ASAP7_75t_R _29977_ (.A1(_07530_),
    .A2(_07531_),
    .B(_07219_),
    .Y(_07532_));
 NAND2x1_ASAP7_75t_SL _29978_ (.A(_07528_),
    .B(_07532_),
    .Y(_07533_));
 AOI21x1_ASAP7_75t_L _29979_ (.A1(_07526_),
    .A2(_07533_),
    .B(_07198_),
    .Y(_07534_));
 AOI21x1_ASAP7_75t_R _29980_ (.A1(_07285_),
    .A2(_07176_),
    .B(_07147_),
    .Y(_07535_));
 NAND2x1_ASAP7_75t_SL _29981_ (.A(_07442_),
    .B(_07274_),
    .Y(_07536_));
 NOR2x1_ASAP7_75t_R _29982_ (.A(_07116_),
    .B(_01384_),
    .Y(_07537_));
 OAI21x1_ASAP7_75t_SL _29983_ (.A1(_07215_),
    .A2(_07537_),
    .B(_07130_),
    .Y(_07538_));
 AOI21x1_ASAP7_75t_R _29984_ (.A1(_07536_),
    .A2(_07538_),
    .B(_07146_),
    .Y(_07539_));
 OAI21x1_ASAP7_75t_R _29985_ (.A1(_07535_),
    .A2(_07539_),
    .B(_07219_),
    .Y(_07540_));
 NAND2x1_ASAP7_75t_SL _29986_ (.A(_07305_),
    .B(_07274_),
    .Y(_07541_));
 AOI21x1_ASAP7_75t_R _29987_ (.A1(_07541_),
    .A2(_07328_),
    .B(_07146_),
    .Y(_07542_));
 NAND2x1_ASAP7_75t_R _29988_ (.A(_07138_),
    .B(_07318_),
    .Y(_07543_));
 OR2x2_ASAP7_75t_R _29989_ (.A(_07138_),
    .B(_01393_),
    .Y(_07544_));
 AND3x1_ASAP7_75t_SL _29990_ (.A(_07543_),
    .B(_07146_),
    .C(_07544_),
    .Y(_07545_));
 OAI21x1_ASAP7_75t_R _29991_ (.A1(_07542_),
    .A2(_07545_),
    .B(_07168_),
    .Y(_07546_));
 AOI21x1_ASAP7_75t_R _29992_ (.A1(_07540_),
    .A2(_07546_),
    .B(_07197_),
    .Y(_07547_));
 OAI21x1_ASAP7_75t_SL _29993_ (.A1(_07534_),
    .A2(_07547_),
    .B(_07250_),
    .Y(_07548_));
 AO21x1_ASAP7_75t_R _29994_ (.A1(_07406_),
    .A2(_07307_),
    .B(_07138_),
    .Y(_07549_));
 OAI21x1_ASAP7_75t_R _29995_ (.A1(_07181_),
    .A2(_07254_),
    .B(_07138_),
    .Y(_07550_));
 AOI21x1_ASAP7_75t_R _29996_ (.A1(_07549_),
    .A2(_07550_),
    .B(_07146_),
    .Y(_07551_));
 AO21x1_ASAP7_75t_R _29997_ (.A1(_07152_),
    .A2(_07136_),
    .B(_07130_),
    .Y(_07552_));
 AOI21x1_ASAP7_75t_SL _29998_ (.A1(_07255_),
    .A2(_07552_),
    .B(_07147_),
    .Y(_07553_));
 OAI21x1_ASAP7_75t_L _29999_ (.A1(_07551_),
    .A2(_07553_),
    .B(_07219_),
    .Y(_07554_));
 AOI21x1_ASAP7_75t_SL _30000_ (.A1(_07432_),
    .A2(_07361_),
    .B(_07147_),
    .Y(_07555_));
 AOI21x1_ASAP7_75t_SL _30001_ (.A1(_07555_),
    .A2(_07275_),
    .B(_07219_),
    .Y(_07556_));
 NOR2x1_ASAP7_75t_SL _30002_ (.A(_07146_),
    .B(_07297_),
    .Y(_07557_));
 NAND3x1_ASAP7_75t_R _30003_ (.A(_07557_),
    .B(_07290_),
    .C(_07543_),
    .Y(_07558_));
 AOI21x1_ASAP7_75t_R _30004_ (.A1(_07556_),
    .A2(_07558_),
    .B(_07197_),
    .Y(_07559_));
 AOI21x1_ASAP7_75t_R _30005_ (.A1(_07554_),
    .A2(_07559_),
    .B(_07250_),
    .Y(_07560_));
 AO21x1_ASAP7_75t_R _30006_ (.A1(_07202_),
    .A2(_07278_),
    .B(_07138_),
    .Y(_07561_));
 AOI21x1_ASAP7_75t_R _30007_ (.A1(_07561_),
    .A2(_07389_),
    .B(_07168_),
    .Y(_07562_));
 NAND2x1_ASAP7_75t_R _30008_ (.A(_07123_),
    .B(_07383_),
    .Y(_07563_));
 AO21x1_ASAP7_75t_R _30009_ (.A1(_07563_),
    .A2(_07538_),
    .B(_07146_),
    .Y(_07564_));
 NOR2x1_ASAP7_75t_SL _30010_ (.A(_07130_),
    .B(_07181_),
    .Y(_07565_));
 OAI21x1_ASAP7_75t_R _30011_ (.A1(_07373_),
    .A2(_07565_),
    .B(_07278_),
    .Y(_07566_));
 NAND2x1_ASAP7_75t_R _30012_ (.A(_07147_),
    .B(_07203_),
    .Y(_07567_));
 OAI21x1_ASAP7_75t_R _30013_ (.A1(_07274_),
    .A2(_07567_),
    .B(_07168_),
    .Y(_07568_));
 AOI21x1_ASAP7_75t_SL _30014_ (.A1(_07146_),
    .A2(_07566_),
    .B(_07568_),
    .Y(_07569_));
 AOI21x1_ASAP7_75t_SL _30015_ (.A1(_07562_),
    .A2(_07564_),
    .B(_07569_),
    .Y(_07570_));
 NAND2x1_ASAP7_75t_R _30016_ (.A(_07197_),
    .B(_07570_),
    .Y(_07571_));
 NAND2x1_ASAP7_75t_SL _30017_ (.A(_07560_),
    .B(_07571_),
    .Y(_07572_));
 NAND2x1_ASAP7_75t_SL _30018_ (.A(_07548_),
    .B(_07572_),
    .Y(_00156_));
 AOI21x1_ASAP7_75t_SL _30019_ (.A1(_07138_),
    .A2(_07468_),
    .B(_07147_),
    .Y(_07573_));
 OAI21x1_ASAP7_75t_SL _30020_ (.A1(_07217_),
    .A2(_07350_),
    .B(_07573_),
    .Y(_07574_));
 INVx1_ASAP7_75t_SL _30021_ (.A(_07240_),
    .Y(_07575_));
 AOI21x1_ASAP7_75t_SL _30022_ (.A1(_07575_),
    .A2(_07557_),
    .B(_07197_),
    .Y(_07576_));
 AOI21x1_ASAP7_75t_SL _30023_ (.A1(_07574_),
    .A2(_07576_),
    .B(_07219_),
    .Y(_07577_));
 AND2x2_ASAP7_75t_SL _30024_ (.A(_07230_),
    .B(_07498_),
    .Y(_07578_));
 AO21x1_ASAP7_75t_SL _30025_ (.A1(_07430_),
    .A2(_07305_),
    .B(_07146_),
    .Y(_07579_));
 AO21x1_ASAP7_75t_SL _30026_ (.A1(_07094_),
    .A2(_07138_),
    .B(_07147_),
    .Y(_07580_));
 OA21x2_ASAP7_75t_SL _30027_ (.A1(_07580_),
    .A2(_07174_),
    .B(_07197_),
    .Y(_07581_));
 OAI21x1_ASAP7_75t_SL _30028_ (.A1(_07578_),
    .A2(_07579_),
    .B(_07581_),
    .Y(_07582_));
 AOI21x1_ASAP7_75t_SL _30029_ (.A1(_07577_),
    .A2(_07582_),
    .B(_07394_),
    .Y(_07583_));
 OA21x2_ASAP7_75t_SL _30030_ (.A1(_07135_),
    .A2(_07130_),
    .B(_07147_),
    .Y(_07584_));
 AO21x1_ASAP7_75t_SL _30031_ (.A1(_07513_),
    .A2(_07406_),
    .B(_07138_),
    .Y(_07585_));
 AOI21x1_ASAP7_75t_SL _30032_ (.A1(_07584_),
    .A2(_07585_),
    .B(_07198_),
    .Y(_07586_));
 AO21x1_ASAP7_75t_SL _30033_ (.A1(_07442_),
    .A2(_07296_),
    .B(_07138_),
    .Y(_07587_));
 NAND2x1_ASAP7_75t_SL _30034_ (.A(_07587_),
    .B(_07210_),
    .Y(_07588_));
 NAND2x1_ASAP7_75t_SL _30035_ (.A(_07586_),
    .B(_07588_),
    .Y(_07589_));
 AO21x1_ASAP7_75t_SL _30036_ (.A1(_07237_),
    .A2(_07406_),
    .B(_07138_),
    .Y(_07590_));
 OA21x2_ASAP7_75t_SL _30037_ (.A1(_07280_),
    .A2(_07185_),
    .B(_07147_),
    .Y(_07591_));
 NAND2x1_ASAP7_75t_SL _30038_ (.A(_07590_),
    .B(_07591_),
    .Y(_07592_));
 OA21x2_ASAP7_75t_SL _30039_ (.A1(_07398_),
    .A2(_07116_),
    .B(_07130_),
    .Y(_07593_));
 AO21x1_ASAP7_75t_SL _30040_ (.A1(_01391_),
    .A2(_07138_),
    .B(_07147_),
    .Y(_07594_));
 OA21x2_ASAP7_75t_SL _30041_ (.A1(_07593_),
    .A2(_07594_),
    .B(_07198_),
    .Y(_07595_));
 AOI21x1_ASAP7_75t_SL _30042_ (.A1(_07592_),
    .A2(_07595_),
    .B(_07168_),
    .Y(_07596_));
 NAND2x1_ASAP7_75t_SL _30043_ (.A(_07589_),
    .B(_07596_),
    .Y(_07597_));
 NAND2x1_ASAP7_75t_SL _30044_ (.A(_07583_),
    .B(_07597_),
    .Y(_07598_));
 AND3x1_ASAP7_75t_SL _30045_ (.A(_07513_),
    .B(_07138_),
    .C(_07135_),
    .Y(_07599_));
 AO21x1_ASAP7_75t_SL _30046_ (.A1(_07226_),
    .A2(_07316_),
    .B(_07146_),
    .Y(_07600_));
 OA21x2_ASAP7_75t_SL _30047_ (.A1(_07081_),
    .A2(_07130_),
    .B(_07146_),
    .Y(_07601_));
 AOI21x1_ASAP7_75t_SL _30048_ (.A1(_07601_),
    .A2(_07538_),
    .B(_07197_),
    .Y(_07602_));
 OA21x2_ASAP7_75t_SL _30049_ (.A1(_07599_),
    .A2(_07600_),
    .B(_07602_),
    .Y(_07603_));
 NOR2x1_ASAP7_75t_SL _30050_ (.A(_07094_),
    .B(_07398_),
    .Y(_07604_));
 INVx1_ASAP7_75t_SL _30051_ (.A(_07430_),
    .Y(_07605_));
 NAND2x1_ASAP7_75t_R _30052_ (.A(_01389_),
    .B(_07203_),
    .Y(_07606_));
 AOI21x1_ASAP7_75t_SL _30053_ (.A1(_07138_),
    .A2(_07606_),
    .B(_07146_),
    .Y(_07607_));
 OAI21x1_ASAP7_75t_SL _30054_ (.A1(_07604_),
    .A2(_07605_),
    .B(_07607_),
    .Y(_07608_));
 AO21x1_ASAP7_75t_SL _30055_ (.A1(_07406_),
    .A2(_07307_),
    .B(_07130_),
    .Y(_07609_));
 NAND3x1_ASAP7_75t_SL _30056_ (.A(_07205_),
    .B(_07609_),
    .C(_07146_),
    .Y(_07610_));
 AOI21x1_ASAP7_75t_SL _30057_ (.A1(_07608_),
    .A2(_07610_),
    .B(_07198_),
    .Y(_07611_));
 NOR2x1_ASAP7_75t_SL _30058_ (.A(_07603_),
    .B(_07611_),
    .Y(_07612_));
 AO21x1_ASAP7_75t_SL _30059_ (.A1(_07463_),
    .A2(_07138_),
    .B(_07186_),
    .Y(_07613_));
 NOR2x1_ASAP7_75t_SL _30060_ (.A(_07146_),
    .B(_07401_),
    .Y(_07614_));
 AOI21x1_ASAP7_75t_SL _30061_ (.A1(_07338_),
    .A2(_07614_),
    .B(_07198_),
    .Y(_07615_));
 OAI21x1_ASAP7_75t_SL _30062_ (.A1(_07147_),
    .A2(_07613_),
    .B(_07615_),
    .Y(_07616_));
 OA21x2_ASAP7_75t_SL _30063_ (.A1(_07261_),
    .A2(_07130_),
    .B(_07147_),
    .Y(_07617_));
 NAND2x1_ASAP7_75t_SL _30064_ (.A(_07398_),
    .B(_07529_),
    .Y(_07618_));
 AOI21x1_ASAP7_75t_SL _30065_ (.A1(_07617_),
    .A2(_07618_),
    .B(_07197_),
    .Y(_07619_));
 AND3x1_ASAP7_75t_SL _30066_ (.A(_07237_),
    .B(_07123_),
    .C(_07138_),
    .Y(_07620_));
 OAI21x1_ASAP7_75t_SL _30067_ (.A1(_07407_),
    .A2(_07620_),
    .B(_07146_),
    .Y(_07621_));
 AOI21x1_ASAP7_75t_SL _30068_ (.A1(_07619_),
    .A2(_07621_),
    .B(_07168_),
    .Y(_07622_));
 AOI21x1_ASAP7_75t_SL _30069_ (.A1(_07616_),
    .A2(_07622_),
    .B(_07250_),
    .Y(_07623_));
 OAI21x1_ASAP7_75t_SL _30070_ (.A1(_07219_),
    .A2(_07612_),
    .B(_07623_),
    .Y(_07624_));
 NAND2x1_ASAP7_75t_SL _30071_ (.A(_07598_),
    .B(_07624_),
    .Y(_00157_));
 NAND2x1_ASAP7_75t_SL _30072_ (.A(_07256_),
    .B(_07361_),
    .Y(_07625_));
 AO21x1_ASAP7_75t_SL _30073_ (.A1(_07337_),
    .A2(_07442_),
    .B(_07130_),
    .Y(_07626_));
 AOI21x1_ASAP7_75t_SL _30074_ (.A1(_07625_),
    .A2(_07626_),
    .B(_07146_),
    .Y(_07627_));
 AOI22x1_ASAP7_75t_SL _30075_ (.A1(_07337_),
    .A2(_07442_),
    .B1(_01384_),
    .B2(_07130_),
    .Y(_07628_));
 OAI21x1_ASAP7_75t_SL _30076_ (.A1(_07147_),
    .A2(_07628_),
    .B(_07168_),
    .Y(_07629_));
 NOR2x1_ASAP7_75t_SL _30077_ (.A(_07627_),
    .B(_07629_),
    .Y(_07630_));
 NOR2x1_ASAP7_75t_SL _30078_ (.A(_07146_),
    .B(_07565_),
    .Y(_07631_));
 NAND2x1_ASAP7_75t_SL _30079_ (.A(_07236_),
    .B(_07631_),
    .Y(_07632_));
 NOR2x1_ASAP7_75t_SL _30080_ (.A(_07138_),
    .B(_07121_),
    .Y(_07633_));
 AOI21x1_ASAP7_75t_SL _30081_ (.A1(_07138_),
    .A2(_07463_),
    .B(_07633_),
    .Y(_07634_));
 NAND2x1_ASAP7_75t_SL _30082_ (.A(_07146_),
    .B(_07634_),
    .Y(_07635_));
 AOI21x1_ASAP7_75t_SL _30083_ (.A1(_07632_),
    .A2(_07635_),
    .B(_07168_),
    .Y(_07636_));
 OAI21x1_ASAP7_75t_SL _30084_ (.A1(_07630_),
    .A2(_07636_),
    .B(_07250_),
    .Y(_07637_));
 OA21x2_ASAP7_75t_SL _30085_ (.A1(_07450_),
    .A2(_07473_),
    .B(_07168_),
    .Y(_07638_));
 NAND2x1_ASAP7_75t_SL _30086_ (.A(_07345_),
    .B(_07415_),
    .Y(_07639_));
 NOR2x1_ASAP7_75t_SL _30087_ (.A(_07168_),
    .B(_07175_),
    .Y(_07640_));
 NOR2x1_ASAP7_75t_SL _30088_ (.A(_07130_),
    .B(_07258_),
    .Y(_07641_));
 AOI21x1_ASAP7_75t_SL _30089_ (.A1(_07319_),
    .A2(_07640_),
    .B(_07641_),
    .Y(_07642_));
 NAND2x1_ASAP7_75t_SL _30090_ (.A(_07639_),
    .B(_07642_),
    .Y(_07643_));
 OAI21x1_ASAP7_75t_SL _30091_ (.A1(_07638_),
    .A2(_07643_),
    .B(_07147_),
    .Y(_07644_));
 NAND2x1_ASAP7_75t_SL _30092_ (.A(_07212_),
    .B(_07430_),
    .Y(_07645_));
 AOI21x1_ASAP7_75t_SL _30093_ (.A1(_07138_),
    .A2(_07270_),
    .B(_07168_),
    .Y(_07646_));
 NAND2x1_ASAP7_75t_SL _30094_ (.A(_07336_),
    .B(_07316_),
    .Y(_07647_));
 NAND3x1_ASAP7_75t_SL _30095_ (.A(_07645_),
    .B(_07646_),
    .C(_07647_),
    .Y(_07648_));
 AO21x1_ASAP7_75t_SL _30096_ (.A1(_07316_),
    .A2(_07305_),
    .B(_07130_),
    .Y(_07649_));
 AO21x1_ASAP7_75t_SL _30097_ (.A1(_01402_),
    .A2(_01396_),
    .B(_07138_),
    .Y(_07650_));
 AND2x2_ASAP7_75t_SL _30098_ (.A(_07650_),
    .B(_07168_),
    .Y(_07651_));
 AOI21x1_ASAP7_75t_SL _30099_ (.A1(_07649_),
    .A2(_07651_),
    .B(_07147_),
    .Y(_07652_));
 AOI21x1_ASAP7_75t_SL _30100_ (.A1(_07648_),
    .A2(_07652_),
    .B(_07250_),
    .Y(_07653_));
 AOI21x1_ASAP7_75t_SL _30101_ (.A1(_07644_),
    .A2(_07653_),
    .B(_07198_),
    .Y(_07654_));
 NAND2x1_ASAP7_75t_SL _30102_ (.A(_07637_),
    .B(_07654_),
    .Y(_07655_));
 AO21x1_ASAP7_75t_SL _30103_ (.A1(_07237_),
    .A2(_07258_),
    .B(_07138_),
    .Y(_07656_));
 OAI21x1_ASAP7_75t_SL _30104_ (.A1(_07207_),
    .A2(_07234_),
    .B(_07138_),
    .Y(_07657_));
 AOI21x1_ASAP7_75t_SL _30105_ (.A1(_07656_),
    .A2(_07657_),
    .B(_07147_),
    .Y(_07658_));
 AO21x1_ASAP7_75t_SL _30106_ (.A1(_07185_),
    .A2(_07130_),
    .B(_07146_),
    .Y(_07659_));
 AOI21x1_ASAP7_75t_SL _30107_ (.A1(_07217_),
    .A2(_07381_),
    .B(_07659_),
    .Y(_07660_));
 OAI21x1_ASAP7_75t_SL _30108_ (.A1(_07658_),
    .A2(_07660_),
    .B(_07168_),
    .Y(_07661_));
 OAI21x1_ASAP7_75t_SL _30109_ (.A1(_07225_),
    .A2(_07254_),
    .B(_07138_),
    .Y(_07662_));
 AOI21x1_ASAP7_75t_SL _30110_ (.A1(_07468_),
    .A2(_07319_),
    .B(_07147_),
    .Y(_07663_));
 NAND2x1_ASAP7_75t_SL _30111_ (.A(_07662_),
    .B(_07663_),
    .Y(_07664_));
 OA21x2_ASAP7_75t_SL _30112_ (.A1(_07135_),
    .A2(_07138_),
    .B(_07147_),
    .Y(_07665_));
 AO21x1_ASAP7_75t_SL _30113_ (.A1(_07442_),
    .A2(_07081_),
    .B(_07130_),
    .Y(_07666_));
 AOI21x1_ASAP7_75t_SL _30114_ (.A1(_07665_),
    .A2(_07666_),
    .B(_07168_),
    .Y(_07667_));
 AOI21x1_ASAP7_75t_SL _30115_ (.A1(_07664_),
    .A2(_07667_),
    .B(_07250_),
    .Y(_07668_));
 AOI21x1_ASAP7_75t_SL _30116_ (.A1(_07661_),
    .A2(_07668_),
    .B(_07197_),
    .Y(_07669_));
 NAND2x1_ASAP7_75t_SL _30117_ (.A(_01397_),
    .B(_07138_),
    .Y(_07670_));
 NAND2x1_ASAP7_75t_SL _30118_ (.A(_07305_),
    .B(_07430_),
    .Y(_07671_));
 AOI21x1_ASAP7_75t_SL _30119_ (.A1(_07670_),
    .A2(_07671_),
    .B(_07147_),
    .Y(_07672_));
 AO21x1_ASAP7_75t_SL _30120_ (.A1(_07237_),
    .A2(_07406_),
    .B(_07130_),
    .Y(_07673_));
 AOI21x1_ASAP7_75t_SL _30121_ (.A1(_07367_),
    .A2(_07673_),
    .B(_07146_),
    .Y(_07674_));
 OAI21x1_ASAP7_75t_SL _30122_ (.A1(_07672_),
    .A2(_07674_),
    .B(_07168_),
    .Y(_07675_));
 INVx1_ASAP7_75t_SL _30123_ (.A(_07269_),
    .Y(_07676_));
 AOI21x1_ASAP7_75t_SL _30124_ (.A1(_07676_),
    .A2(_07541_),
    .B(_07146_),
    .Y(_07677_));
 AOI21x1_ASAP7_75t_SL _30125_ (.A1(_07305_),
    .A2(_07409_),
    .B(_07147_),
    .Y(_07678_));
 OAI21x1_ASAP7_75t_SL _30126_ (.A1(_07677_),
    .A2(_07678_),
    .B(_07219_),
    .Y(_07679_));
 NAND3x1_ASAP7_75t_SL _30127_ (.A(_07679_),
    .B(_07250_),
    .C(_07675_),
    .Y(_07680_));
 NAND2x1_ASAP7_75t_SL _30128_ (.A(_07669_),
    .B(_07680_),
    .Y(_07681_));
 NAND2x1_ASAP7_75t_SL _30129_ (.A(_07655_),
    .B(_07681_),
    .Y(_00158_));
 NAND2x1_ASAP7_75t_SL _30130_ (.A(_07130_),
    .B(_07116_),
    .Y(_07682_));
 OAI21x1_ASAP7_75t_SL _30131_ (.A1(_07279_),
    .A2(_07324_),
    .B(_07682_),
    .Y(_07683_));
 AOI21x1_ASAP7_75t_SL _30132_ (.A1(_07147_),
    .A2(_07683_),
    .B(_07219_),
    .Y(_07684_));
 INVx1_ASAP7_75t_SL _30133_ (.A(_07309_),
    .Y(_07685_));
 AO21x1_ASAP7_75t_SL _30134_ (.A1(_07685_),
    .A2(_07398_),
    .B(_07138_),
    .Y(_07686_));
 NAND2x1_ASAP7_75t_SL _30135_ (.A(_07389_),
    .B(_07686_),
    .Y(_07687_));
 NAND2x1_ASAP7_75t_SL _30136_ (.A(_07684_),
    .B(_07687_),
    .Y(_07688_));
 NAND2x1_ASAP7_75t_SL _30137_ (.A(_07138_),
    .B(_07303_),
    .Y(_07689_));
 NOR2x1_ASAP7_75t_SL _30138_ (.A(_07147_),
    .B(_07480_),
    .Y(_07690_));
 AOI21x1_ASAP7_75t_SL _30139_ (.A1(_07689_),
    .A2(_07690_),
    .B(_07168_),
    .Y(_07691_));
 NAND2x1_ASAP7_75t_SL _30140_ (.A(_07493_),
    .B(_07182_),
    .Y(_07692_));
 AOI21x1_ASAP7_75t_SL _30141_ (.A1(_07138_),
    .A2(_07268_),
    .B(_07146_),
    .Y(_07693_));
 NAND2x1_ASAP7_75t_SL _30142_ (.A(_07692_),
    .B(_07693_),
    .Y(_07694_));
 AOI21x1_ASAP7_75t_SL _30143_ (.A1(_07691_),
    .A2(_07694_),
    .B(_07197_),
    .Y(_07695_));
 AOI21x1_ASAP7_75t_SL _30144_ (.A1(_07688_),
    .A2(_07695_),
    .B(_07394_),
    .Y(_07696_));
 AOI21x1_ASAP7_75t_SL _30145_ (.A1(_07327_),
    .A2(_07476_),
    .B(_07146_),
    .Y(_07697_));
 AOI21x1_ASAP7_75t_SL _30146_ (.A1(_07645_),
    .A2(_07443_),
    .B(_07147_),
    .Y(_07698_));
 OAI21x1_ASAP7_75t_SL _30147_ (.A1(_07697_),
    .A2(_07698_),
    .B(_07219_),
    .Y(_07699_));
 NOR2x1_ASAP7_75t_SL _30148_ (.A(_07147_),
    .B(_07361_),
    .Y(_07700_));
 AOI21x1_ASAP7_75t_SL _30149_ (.A1(_07541_),
    .A2(_07700_),
    .B(_07219_),
    .Y(_07701_));
 AO21x1_ASAP7_75t_SL _30150_ (.A1(_07685_),
    .A2(_07136_),
    .B(_07130_),
    .Y(_07702_));
 OA21x2_ASAP7_75t_SL _30151_ (.A1(_07604_),
    .A2(_07349_),
    .B(_07147_),
    .Y(_07703_));
 NAND2x1_ASAP7_75t_SL _30152_ (.A(_07702_),
    .B(_07703_),
    .Y(_07704_));
 AOI21x1_ASAP7_75t_SL _30153_ (.A1(_07701_),
    .A2(_07704_),
    .B(_07198_),
    .Y(_07705_));
 NAND2x1_ASAP7_75t_SL _30154_ (.A(_07699_),
    .B(_07705_),
    .Y(_07706_));
 NAND2x1_ASAP7_75t_SL _30155_ (.A(_07696_),
    .B(_07706_),
    .Y(_07707_));
 INVx1_ASAP7_75t_SL _30156_ (.A(_07523_),
    .Y(_07708_));
 AND3x1_ASAP7_75t_SL _30157_ (.A(_07337_),
    .B(_07152_),
    .C(_07130_),
    .Y(_07709_));
 NAND2x1_ASAP7_75t_SL _30158_ (.A(_01393_),
    .B(_07138_),
    .Y(_07710_));
 AOI21x1_ASAP7_75t_SL _30159_ (.A1(_07710_),
    .A2(_07259_),
    .B(_07219_),
    .Y(_07711_));
 OAI21x1_ASAP7_75t_SL _30160_ (.A1(_07708_),
    .A2(_07709_),
    .B(_07711_),
    .Y(_07712_));
 NAND2x1_ASAP7_75t_SL _30161_ (.A(_07130_),
    .B(_07156_),
    .Y(_07713_));
 OAI21x1_ASAP7_75t_SL _30162_ (.A1(_01402_),
    .A2(_07130_),
    .B(_07146_),
    .Y(_07714_));
 NOR2x1_ASAP7_75t_SL _30163_ (.A(_07714_),
    .B(_07411_),
    .Y(_07715_));
 AOI21x1_ASAP7_75t_SL _30164_ (.A1(_07713_),
    .A2(_07715_),
    .B(_07168_),
    .Y(_07716_));
 AO21x1_ASAP7_75t_SL _30165_ (.A1(_07237_),
    .A2(_07261_),
    .B(_07130_),
    .Y(_07717_));
 AOI21x1_ASAP7_75t_SL _30166_ (.A1(_07305_),
    .A2(_07226_),
    .B(_07146_),
    .Y(_07718_));
 NAND2x1_ASAP7_75t_SL _30167_ (.A(_07717_),
    .B(_07718_),
    .Y(_07719_));
 AOI21x1_ASAP7_75t_SL _30168_ (.A1(_07716_),
    .A2(_07719_),
    .B(_07197_),
    .Y(_07720_));
 AOI21x1_ASAP7_75t_SL _30169_ (.A1(_07712_),
    .A2(_07720_),
    .B(_07250_),
    .Y(_07721_));
 NAND2x1_ASAP7_75t_SL _30170_ (.A(_07305_),
    .B(_07316_),
    .Y(_07722_));
 NOR2x1_ASAP7_75t_SL _30171_ (.A(_01389_),
    .B(_07138_),
    .Y(_07723_));
 AOI21x1_ASAP7_75t_SL _30172_ (.A1(_07138_),
    .A2(_07722_),
    .B(_07723_),
    .Y(_07724_));
 OA21x2_ASAP7_75t_SL _30173_ (.A1(_01385_),
    .A2(_07112_),
    .B(_07146_),
    .Y(_07725_));
 OAI21x1_ASAP7_75t_SL _30174_ (.A1(_07529_),
    .A2(_07565_),
    .B(_07725_),
    .Y(_07726_));
 OAI21x1_ASAP7_75t_SL _30175_ (.A1(_07146_),
    .A2(_07724_),
    .B(_07726_),
    .Y(_07727_));
 AOI21x1_ASAP7_75t_SL _30176_ (.A1(_07219_),
    .A2(_07727_),
    .B(_07198_),
    .Y(_07728_));
 OA21x2_ASAP7_75t_SL _30177_ (.A1(_07280_),
    .A2(_07492_),
    .B(_07146_),
    .Y(_07729_));
 AO21x1_ASAP7_75t_SL _30178_ (.A1(_07685_),
    .A2(_07136_),
    .B(_07138_),
    .Y(_07730_));
 AOI21x1_ASAP7_75t_SL _30179_ (.A1(_07729_),
    .A2(_07730_),
    .B(_07219_),
    .Y(_07731_));
 AO221x1_ASAP7_75t_SL _30180_ (.A1(_07468_),
    .A2(_07274_),
    .B1(_07316_),
    .B2(_07282_),
    .C(_07146_),
    .Y(_07732_));
 NAND2x1_ASAP7_75t_SL _30181_ (.A(_07731_),
    .B(_07732_),
    .Y(_07733_));
 NAND2x1_ASAP7_75t_SL _30182_ (.A(_07728_),
    .B(_07733_),
    .Y(_07734_));
 NAND2x1_ASAP7_75t_SL _30183_ (.A(_07721_),
    .B(_07734_),
    .Y(_07735_));
 NAND2x1_ASAP7_75t_SL _30184_ (.A(_07707_),
    .B(_07735_),
    .Y(_00159_));
 INVx1_ASAP7_75t_R _30185_ (.A(_00488_),
    .Y(text_out[9]));
 INVx1_ASAP7_75t_R _30186_ (.A(_00573_),
    .Y(done));
 INVx1_ASAP7_75t_R _30187_ (.A(_00702_),
    .Y(text_out[0]));
 INVx1_ASAP7_75t_R _30188_ (.A(_00703_),
    .Y(text_out[100]));
 INVx1_ASAP7_75t_R _30189_ (.A(_00704_),
    .Y(text_out[101]));
 INVx1_ASAP7_75t_R _30190_ (.A(_00705_),
    .Y(text_out[102]));
 INVx1_ASAP7_75t_R _30191_ (.A(_00706_),
    .Y(text_out[103]));
 INVx1_ASAP7_75t_R _30192_ (.A(_00707_),
    .Y(text_out[104]));
 INVx1_ASAP7_75t_R _30193_ (.A(_00708_),
    .Y(text_out[105]));
 INVx1_ASAP7_75t_R _30194_ (.A(_00709_),
    .Y(text_out[106]));
 INVx1_ASAP7_75t_R _30195_ (.A(_00710_),
    .Y(text_out[107]));
 INVx1_ASAP7_75t_R _30196_ (.A(_00711_),
    .Y(text_out[108]));
 INVx1_ASAP7_75t_R _30197_ (.A(_00712_),
    .Y(text_out[109]));
 INVx1_ASAP7_75t_R _30198_ (.A(_00713_),
    .Y(text_out[10]));
 INVx1_ASAP7_75t_R _30199_ (.A(_00714_),
    .Y(text_out[110]));
 INVx1_ASAP7_75t_R _30200_ (.A(_00715_),
    .Y(text_out[111]));
 INVx1_ASAP7_75t_R _30201_ (.A(_00716_),
    .Y(text_out[112]));
 INVx1_ASAP7_75t_R _30202_ (.A(_00717_),
    .Y(text_out[113]));
 INVx1_ASAP7_75t_R _30203_ (.A(_00718_),
    .Y(text_out[114]));
 INVx1_ASAP7_75t_R _30204_ (.A(_00719_),
    .Y(text_out[115]));
 INVx1_ASAP7_75t_R _30205_ (.A(_00720_),
    .Y(text_out[116]));
 INVx1_ASAP7_75t_R _30206_ (.A(_00721_),
    .Y(text_out[117]));
 INVx1_ASAP7_75t_R _30207_ (.A(_00722_),
    .Y(text_out[118]));
 INVx1_ASAP7_75t_R _30208_ (.A(_00723_),
    .Y(text_out[119]));
 INVx1_ASAP7_75t_R _30209_ (.A(_00724_),
    .Y(text_out[11]));
 INVx1_ASAP7_75t_R _30210_ (.A(_00725_),
    .Y(text_out[120]));
 INVx1_ASAP7_75t_R _30211_ (.A(_00726_),
    .Y(text_out[121]));
 INVx1_ASAP7_75t_R _30212_ (.A(_00727_),
    .Y(text_out[122]));
 INVx1_ASAP7_75t_R _30213_ (.A(_00728_),
    .Y(text_out[123]));
 INVx1_ASAP7_75t_R _30214_ (.A(_00729_),
    .Y(text_out[124]));
 INVx1_ASAP7_75t_R _30215_ (.A(_00730_),
    .Y(text_out[125]));
 INVx1_ASAP7_75t_R _30216_ (.A(_00731_),
    .Y(text_out[126]));
 INVx1_ASAP7_75t_R _30217_ (.A(_00732_),
    .Y(text_out[127]));
 INVx1_ASAP7_75t_R _30218_ (.A(_00733_),
    .Y(text_out[12]));
 INVx1_ASAP7_75t_R _30219_ (.A(_00734_),
    .Y(text_out[13]));
 INVx1_ASAP7_75t_R _30220_ (.A(_00735_),
    .Y(text_out[14]));
 INVx1_ASAP7_75t_R _30221_ (.A(_00736_),
    .Y(text_out[15]));
 INVx1_ASAP7_75t_R _30222_ (.A(_00737_),
    .Y(text_out[16]));
 INVx1_ASAP7_75t_R _30223_ (.A(_00738_),
    .Y(text_out[17]));
 INVx1_ASAP7_75t_R _30224_ (.A(_00739_),
    .Y(text_out[18]));
 INVx1_ASAP7_75t_R _30225_ (.A(_00740_),
    .Y(text_out[19]));
 INVx1_ASAP7_75t_R _30226_ (.A(_00741_),
    .Y(text_out[1]));
 INVx1_ASAP7_75t_R _30227_ (.A(_00742_),
    .Y(text_out[20]));
 INVx1_ASAP7_75t_R _30228_ (.A(_00743_),
    .Y(text_out[21]));
 INVx1_ASAP7_75t_R _30229_ (.A(_00744_),
    .Y(text_out[22]));
 INVx1_ASAP7_75t_R _30230_ (.A(_00745_),
    .Y(text_out[23]));
 INVx1_ASAP7_75t_R _30231_ (.A(_00746_),
    .Y(text_out[24]));
 INVx1_ASAP7_75t_R _30232_ (.A(_00747_),
    .Y(text_out[25]));
 INVx1_ASAP7_75t_R _30233_ (.A(_00748_),
    .Y(text_out[26]));
 INVx1_ASAP7_75t_R _30234_ (.A(_00749_),
    .Y(text_out[27]));
 INVx1_ASAP7_75t_R _30235_ (.A(_00750_),
    .Y(text_out[28]));
 INVx1_ASAP7_75t_R _30236_ (.A(_00751_),
    .Y(text_out[29]));
 INVx1_ASAP7_75t_R _30237_ (.A(_00752_),
    .Y(text_out[2]));
 INVx1_ASAP7_75t_R _30238_ (.A(_00753_),
    .Y(text_out[30]));
 INVx1_ASAP7_75t_R _30239_ (.A(_00754_),
    .Y(text_out[31]));
 INVx1_ASAP7_75t_R _30240_ (.A(_00755_),
    .Y(text_out[32]));
 INVx1_ASAP7_75t_R _30241_ (.A(_00756_),
    .Y(text_out[33]));
 INVx1_ASAP7_75t_R _30242_ (.A(_00757_),
    .Y(text_out[34]));
 INVx1_ASAP7_75t_R _30243_ (.A(_00758_),
    .Y(text_out[35]));
 INVx1_ASAP7_75t_R _30244_ (.A(_00759_),
    .Y(text_out[36]));
 INVx1_ASAP7_75t_R _30245_ (.A(_00760_),
    .Y(text_out[37]));
 INVx1_ASAP7_75t_R _30246_ (.A(_00761_),
    .Y(text_out[38]));
 INVx1_ASAP7_75t_R _30247_ (.A(_00762_),
    .Y(text_out[39]));
 INVx1_ASAP7_75t_R _30248_ (.A(_00763_),
    .Y(text_out[3]));
 INVx1_ASAP7_75t_R _30249_ (.A(_00764_),
    .Y(text_out[40]));
 INVx1_ASAP7_75t_R _30250_ (.A(_00765_),
    .Y(text_out[41]));
 INVx1_ASAP7_75t_R _30251_ (.A(_00766_),
    .Y(text_out[42]));
 INVx1_ASAP7_75t_R _30252_ (.A(_00767_),
    .Y(text_out[43]));
 INVx1_ASAP7_75t_R _30253_ (.A(_00768_),
    .Y(text_out[44]));
 INVx1_ASAP7_75t_R _30254_ (.A(_00769_),
    .Y(text_out[45]));
 INVx1_ASAP7_75t_R _30255_ (.A(_00770_),
    .Y(text_out[46]));
 INVx1_ASAP7_75t_R _30256_ (.A(_00771_),
    .Y(text_out[47]));
 INVx1_ASAP7_75t_R _30257_ (.A(_00772_),
    .Y(text_out[48]));
 INVx1_ASAP7_75t_R _30258_ (.A(_00773_),
    .Y(text_out[49]));
 INVx1_ASAP7_75t_R _30259_ (.A(_00774_),
    .Y(text_out[4]));
 INVx1_ASAP7_75t_R _30260_ (.A(_00775_),
    .Y(text_out[50]));
 INVx1_ASAP7_75t_R _30261_ (.A(_00776_),
    .Y(text_out[51]));
 INVx1_ASAP7_75t_R _30262_ (.A(_00777_),
    .Y(text_out[52]));
 INVx1_ASAP7_75t_R _30263_ (.A(_00778_),
    .Y(text_out[53]));
 INVx1_ASAP7_75t_R _30264_ (.A(_00779_),
    .Y(text_out[54]));
 INVx1_ASAP7_75t_R _30265_ (.A(_00780_),
    .Y(text_out[55]));
 INVx1_ASAP7_75t_R _30266_ (.A(_00781_),
    .Y(text_out[56]));
 INVx1_ASAP7_75t_R _30267_ (.A(_00782_),
    .Y(text_out[57]));
 INVx1_ASAP7_75t_R _30268_ (.A(_00783_),
    .Y(text_out[58]));
 INVx1_ASAP7_75t_R _30269_ (.A(_00784_),
    .Y(text_out[59]));
 INVx1_ASAP7_75t_R _30270_ (.A(_00785_),
    .Y(text_out[5]));
 INVx1_ASAP7_75t_R _30271_ (.A(_00786_),
    .Y(text_out[60]));
 INVx1_ASAP7_75t_R _30272_ (.A(_00787_),
    .Y(text_out[61]));
 INVx1_ASAP7_75t_R _30273_ (.A(_00788_),
    .Y(text_out[62]));
 INVx1_ASAP7_75t_R _30274_ (.A(_00789_),
    .Y(text_out[63]));
 INVx1_ASAP7_75t_R _30275_ (.A(_00790_),
    .Y(text_out[64]));
 INVx1_ASAP7_75t_R _30276_ (.A(_00791_),
    .Y(text_out[65]));
 INVx1_ASAP7_75t_R _30277_ (.A(_00792_),
    .Y(text_out[66]));
 INVx1_ASAP7_75t_R _30278_ (.A(_00793_),
    .Y(text_out[67]));
 INVx1_ASAP7_75t_R _30279_ (.A(_00794_),
    .Y(text_out[68]));
 INVx1_ASAP7_75t_R _30280_ (.A(_00795_),
    .Y(text_out[69]));
 INVx1_ASAP7_75t_R _30281_ (.A(_00796_),
    .Y(text_out[6]));
 INVx1_ASAP7_75t_R _30282_ (.A(_00797_),
    .Y(text_out[70]));
 INVx1_ASAP7_75t_R _30283_ (.A(_00798_),
    .Y(text_out[71]));
 INVx1_ASAP7_75t_R _30284_ (.A(_00799_),
    .Y(text_out[72]));
 INVx1_ASAP7_75t_R _30285_ (.A(_00800_),
    .Y(text_out[73]));
 INVx1_ASAP7_75t_R _30286_ (.A(_00801_),
    .Y(text_out[74]));
 INVx1_ASAP7_75t_R _30287_ (.A(_00802_),
    .Y(text_out[75]));
 INVx1_ASAP7_75t_R _30288_ (.A(_00803_),
    .Y(text_out[76]));
 INVx1_ASAP7_75t_R _30289_ (.A(_00804_),
    .Y(text_out[77]));
 INVx1_ASAP7_75t_R _30290_ (.A(_00805_),
    .Y(text_out[78]));
 INVx1_ASAP7_75t_R _30291_ (.A(_00806_),
    .Y(text_out[79]));
 INVx1_ASAP7_75t_R _30292_ (.A(_00807_),
    .Y(text_out[7]));
 INVx1_ASAP7_75t_R _30293_ (.A(_00808_),
    .Y(text_out[80]));
 INVx1_ASAP7_75t_R _30294_ (.A(_00809_),
    .Y(text_out[81]));
 INVx1_ASAP7_75t_R _30295_ (.A(_00810_),
    .Y(text_out[82]));
 INVx1_ASAP7_75t_R _30296_ (.A(_00811_),
    .Y(text_out[83]));
 INVx1_ASAP7_75t_R _30297_ (.A(_00812_),
    .Y(text_out[84]));
 INVx1_ASAP7_75t_R _30298_ (.A(_00813_),
    .Y(text_out[85]));
 INVx1_ASAP7_75t_R _30299_ (.A(_00814_),
    .Y(text_out[86]));
 INVx1_ASAP7_75t_R _30300_ (.A(_00815_),
    .Y(text_out[87]));
 INVx1_ASAP7_75t_R _30301_ (.A(_00816_),
    .Y(text_out[88]));
 INVx1_ASAP7_75t_R _30302_ (.A(_00817_),
    .Y(text_out[89]));
 INVx1_ASAP7_75t_R _30303_ (.A(_00818_),
    .Y(text_out[8]));
 INVx1_ASAP7_75t_R _30304_ (.A(_00819_),
    .Y(text_out[90]));
 INVx1_ASAP7_75t_R _30305_ (.A(_00820_),
    .Y(text_out[91]));
 INVx1_ASAP7_75t_R _30306_ (.A(_00821_),
    .Y(text_out[92]));
 INVx1_ASAP7_75t_R _30307_ (.A(_00822_),
    .Y(text_out[93]));
 INVx1_ASAP7_75t_R _30308_ (.A(_00823_),
    .Y(text_out[94]));
 INVx1_ASAP7_75t_R _30309_ (.A(_00824_),
    .Y(text_out[95]));
 INVx1_ASAP7_75t_R _30310_ (.A(_00825_),
    .Y(text_out[96]));
 INVx1_ASAP7_75t_R _30311_ (.A(_00826_),
    .Y(text_out[97]));
 INVx1_ASAP7_75t_R _30312_ (.A(_00827_),
    .Y(text_out[98]));
 INVx1_ASAP7_75t_R _30313_ (.A(_00828_),
    .Y(text_out[99]));
 NOR2x1_ASAP7_75t_R _30315_ (.A(ld),
    .B(_00409_),
    .Y(_07737_));
 AO21x1_ASAP7_75t_R _30316_ (.A1(ld),
    .A2(text_in[0]),
    .B(_07737_),
    .Y(_01408_));
 NOR2x1_ASAP7_75t_R _30317_ (.A(ld),
    .B(_00568_),
    .Y(_07738_));
 AO21x1_ASAP7_75t_R _30318_ (.A1(ld),
    .A2(text_in[100]),
    .B(_07738_),
    .Y(_01409_));
 NOR2x1_ASAP7_75t_R _30320_ (.A(ld),
    .B(_00567_),
    .Y(_07740_));
 AO21x1_ASAP7_75t_R _30321_ (.A1(ld),
    .A2(text_in[101]),
    .B(_07740_),
    .Y(_01410_));
 NOR2x1_ASAP7_75t_R _30322_ (.A(ld),
    .B(_00566_),
    .Y(_07741_));
 AO21x1_ASAP7_75t_R _30323_ (.A1(ld),
    .A2(text_in[102]),
    .B(_07741_),
    .Y(_01411_));
 NOR2x1_ASAP7_75t_R _30324_ (.A(ld),
    .B(_00565_),
    .Y(_07742_));
 AO21x1_ASAP7_75t_R _30325_ (.A1(ld),
    .A2(text_in[103]),
    .B(_07742_),
    .Y(_01412_));
 NOR2x1_ASAP7_75t_R _30326_ (.A(ld),
    .B(_00469_),
    .Y(_07743_));
 AO21x1_ASAP7_75t_R _30327_ (.A1(ld),
    .A2(text_in[104]),
    .B(_07743_),
    .Y(_01413_));
 NOR2x1_ASAP7_75t_R _30328_ (.A(ld),
    .B(_00468_),
    .Y(_07744_));
 AO21x1_ASAP7_75t_R _30329_ (.A1(ld),
    .A2(text_in[105]),
    .B(_07744_),
    .Y(_01414_));
 NOR2x1_ASAP7_75t_R _30330_ (.A(ld),
    .B(_00470_),
    .Y(_07745_));
 AO21x1_ASAP7_75t_R _30331_ (.A1(ld),
    .A2(text_in[106]),
    .B(_07745_),
    .Y(_01415_));
 NOR2x1_ASAP7_75t_R _30332_ (.A(ld),
    .B(_00564_),
    .Y(_07746_));
 AO21x1_ASAP7_75t_R _30333_ (.A1(ld),
    .A2(text_in[107]),
    .B(_07746_),
    .Y(_01416_));
 NOR2x1_ASAP7_75t_R _30334_ (.A(ld),
    .B(_00563_),
    .Y(_07747_));
 AO21x1_ASAP7_75t_R _30335_ (.A1(ld),
    .A2(text_in[108]),
    .B(_07747_),
    .Y(_01417_));
 NOR2x1_ASAP7_75t_R _30337_ (.A(ld),
    .B(_00562_),
    .Y(_07749_));
 AO21x1_ASAP7_75t_R _30338_ (.A1(ld),
    .A2(text_in[109]),
    .B(_07749_),
    .Y(_01418_));
 NOR2x1_ASAP7_75t_R _30339_ (.A(ld),
    .B(_00479_),
    .Y(_07750_));
 AO21x1_ASAP7_75t_R _30340_ (.A1(ld),
    .A2(text_in[10]),
    .B(_07750_),
    .Y(_01419_));
 NOR2x1_ASAP7_75t_R _30342_ (.A(ld),
    .B(_00561_),
    .Y(_07752_));
 AO21x1_ASAP7_75t_R _30343_ (.A1(ld),
    .A2(text_in[110]),
    .B(_07752_),
    .Y(_01420_));
 NOR2x1_ASAP7_75t_R _30344_ (.A(ld),
    .B(_00560_),
    .Y(_07753_));
 AO21x1_ASAP7_75t_R _30345_ (.A1(ld),
    .A2(text_in[111]),
    .B(_07753_),
    .Y(_01421_));
 NOR2x1_ASAP7_75t_R _30346_ (.A(ld),
    .B(_00457_),
    .Y(_07754_));
 AO21x1_ASAP7_75t_R _30347_ (.A1(ld),
    .A2(text_in[112]),
    .B(_07754_),
    .Y(_01422_));
 NOR2x1_ASAP7_75t_R _30348_ (.A(ld),
    .B(_00456_),
    .Y(_07755_));
 AO21x1_ASAP7_75t_R _30349_ (.A1(ld),
    .A2(text_in[113]),
    .B(_07755_),
    .Y(_01423_));
 NOR2x1_ASAP7_75t_R _30350_ (.A(ld),
    .B(_00458_),
    .Y(_07756_));
 AO21x1_ASAP7_75t_R _30351_ (.A1(ld),
    .A2(text_in[114]),
    .B(_07756_),
    .Y(_01424_));
 NOR2x1_ASAP7_75t_R _30352_ (.A(ld),
    .B(_00559_),
    .Y(_07757_));
 AO21x1_ASAP7_75t_R _30353_ (.A1(ld),
    .A2(text_in[115]),
    .B(_07757_),
    .Y(_01425_));
 NOR2x1_ASAP7_75t_R _30354_ (.A(ld),
    .B(_00558_),
    .Y(_07758_));
 AO21x1_ASAP7_75t_R _30355_ (.A1(ld),
    .A2(text_in[116]),
    .B(_07758_),
    .Y(_01426_));
 NOR2x1_ASAP7_75t_R _30356_ (.A(ld),
    .B(_00557_),
    .Y(_07759_));
 AO21x1_ASAP7_75t_R _30357_ (.A1(ld),
    .A2(text_in[117]),
    .B(_07759_),
    .Y(_01427_));
 NOR2x1_ASAP7_75t_R _30359_ (.A(ld),
    .B(_00556_),
    .Y(_07761_));
 AO21x1_ASAP7_75t_R _30360_ (.A1(ld),
    .A2(text_in[118]),
    .B(_07761_),
    .Y(_01428_));
 NOR2x1_ASAP7_75t_R _30361_ (.A(ld),
    .B(_00555_),
    .Y(_07762_));
 AO21x1_ASAP7_75t_R _30362_ (.A1(ld),
    .A2(text_in[119]),
    .B(_07762_),
    .Y(_01429_));
 NOR2x1_ASAP7_75t_R _30364_ (.A(ld),
    .B(_00554_),
    .Y(_07764_));
 AO21x1_ASAP7_75t_R _30365_ (.A1(ld),
    .A2(text_in[11]),
    .B(_07764_),
    .Y(_01430_));
 NOR2x1_ASAP7_75t_R _30366_ (.A(ld),
    .B(_00445_),
    .Y(_07765_));
 AO21x1_ASAP7_75t_R _30367_ (.A1(ld),
    .A2(text_in[120]),
    .B(_07765_),
    .Y(_01431_));
 NOR2x1_ASAP7_75t_R _30368_ (.A(ld),
    .B(_00444_),
    .Y(_07766_));
 AO21x1_ASAP7_75t_R _30369_ (.A1(ld),
    .A2(text_in[121]),
    .B(_07766_),
    .Y(_01432_));
 NOR2x1_ASAP7_75t_R _30370_ (.A(ld),
    .B(_00446_),
    .Y(_07767_));
 AO21x1_ASAP7_75t_R _30371_ (.A1(ld),
    .A2(text_in[122]),
    .B(_07767_),
    .Y(_01433_));
 NOR2x1_ASAP7_75t_R _30372_ (.A(ld),
    .B(_00553_),
    .Y(_07768_));
 AO21x1_ASAP7_75t_R _30373_ (.A1(ld),
    .A2(text_in[123]),
    .B(_07768_),
    .Y(_01434_));
 NOR2x1_ASAP7_75t_R _30374_ (.A(ld),
    .B(_00552_),
    .Y(_07769_));
 AO21x1_ASAP7_75t_R _30375_ (.A1(ld),
    .A2(text_in[124]),
    .B(_07769_),
    .Y(_01435_));
 NOR2x1_ASAP7_75t_R _30376_ (.A(ld),
    .B(_00551_),
    .Y(_07770_));
 AO21x1_ASAP7_75t_R _30377_ (.A1(ld),
    .A2(text_in[125]),
    .B(_07770_),
    .Y(_01436_));
 NOR2x1_ASAP7_75t_R _30378_ (.A(ld),
    .B(_00550_),
    .Y(_07771_));
 AO21x1_ASAP7_75t_R _30379_ (.A1(ld),
    .A2(text_in[126]),
    .B(_07771_),
    .Y(_01437_));
 NOR2x1_ASAP7_75t_R _30381_ (.A(ld),
    .B(_00549_),
    .Y(_07773_));
 AO21x1_ASAP7_75t_R _30382_ (.A1(ld),
    .A2(text_in[127]),
    .B(_07773_),
    .Y(_01438_));
 NOR2x1_ASAP7_75t_R _30383_ (.A(ld),
    .B(_00548_),
    .Y(_07774_));
 AO21x1_ASAP7_75t_R _30384_ (.A1(ld),
    .A2(text_in[12]),
    .B(_07774_),
    .Y(_01439_));
 NOR2x1_ASAP7_75t_R _30386_ (.A(ld),
    .B(_00547_),
    .Y(_07776_));
 AO21x1_ASAP7_75t_R _30387_ (.A1(ld),
    .A2(text_in[13]),
    .B(_07776_),
    .Y(_01440_));
 NOR2x1_ASAP7_75t_R _30388_ (.A(ld),
    .B(_00546_),
    .Y(_07777_));
 AO21x1_ASAP7_75t_R _30389_ (.A1(ld),
    .A2(text_in[14]),
    .B(_07777_),
    .Y(_01441_));
 NOR2x1_ASAP7_75t_R _30390_ (.A(ld),
    .B(_00545_),
    .Y(_07778_));
 AO21x1_ASAP7_75t_R _30391_ (.A1(ld),
    .A2(text_in[15]),
    .B(_07778_),
    .Y(_01442_));
 NOR2x1_ASAP7_75t_R _30392_ (.A(ld),
    .B(_00466_),
    .Y(_07779_));
 AO21x1_ASAP7_75t_R _30393_ (.A1(ld),
    .A2(text_in[16]),
    .B(_07779_),
    .Y(_01443_));
 NOR2x1_ASAP7_75t_R _30394_ (.A(ld),
    .B(_00465_),
    .Y(_07780_));
 AO21x1_ASAP7_75t_R _30395_ (.A1(ld),
    .A2(text_in[17]),
    .B(_07780_),
    .Y(_01444_));
 NOR2x1_ASAP7_75t_R _30396_ (.A(ld),
    .B(_00467_),
    .Y(_07781_));
 AO21x1_ASAP7_75t_R _30397_ (.A1(ld),
    .A2(text_in[18]),
    .B(_07781_),
    .Y(_01445_));
 NOR2x1_ASAP7_75t_R _30398_ (.A(ld),
    .B(_00544_),
    .Y(_07782_));
 AO21x1_ASAP7_75t_R _30399_ (.A1(ld),
    .A2(text_in[19]),
    .B(_07782_),
    .Y(_01446_));
 NOR2x1_ASAP7_75t_R _30400_ (.A(ld),
    .B(_00408_),
    .Y(_07783_));
 AO21x1_ASAP7_75t_R _30401_ (.A1(ld),
    .A2(text_in[1]),
    .B(_07783_),
    .Y(_01447_));
 NOR2x1_ASAP7_75t_R _30403_ (.A(ld),
    .B(_00543_),
    .Y(_07785_));
 AO21x1_ASAP7_75t_R _30404_ (.A1(ld),
    .A2(text_in[20]),
    .B(_07785_),
    .Y(_01448_));
 NOR2x1_ASAP7_75t_R _30405_ (.A(ld),
    .B(_00542_),
    .Y(_07786_));
 AO21x1_ASAP7_75t_R _30406_ (.A1(ld),
    .A2(text_in[21]),
    .B(_07786_),
    .Y(_01449_));
 NOR2x1_ASAP7_75t_R _30408_ (.A(ld),
    .B(_00541_),
    .Y(_07788_));
 AO21x1_ASAP7_75t_R _30409_ (.A1(ld),
    .A2(text_in[22]),
    .B(_07788_),
    .Y(_01450_));
 NOR2x1_ASAP7_75t_R _30410_ (.A(ld),
    .B(_00540_),
    .Y(_07789_));
 AO21x1_ASAP7_75t_R _30411_ (.A1(ld),
    .A2(text_in[23]),
    .B(_07789_),
    .Y(_01451_));
 NOR2x1_ASAP7_75t_R _30412_ (.A(ld),
    .B(_00454_),
    .Y(_07790_));
 AO21x1_ASAP7_75t_R _30413_ (.A1(ld),
    .A2(text_in[24]),
    .B(_07790_),
    .Y(_01452_));
 NOR2x1_ASAP7_75t_R _30414_ (.A(ld),
    .B(_00453_),
    .Y(_07791_));
 AO21x1_ASAP7_75t_R _30415_ (.A1(ld),
    .A2(text_in[25]),
    .B(_07791_),
    .Y(_01453_));
 NOR2x1_ASAP7_75t_R _30416_ (.A(ld),
    .B(_00455_),
    .Y(_07792_));
 AO21x1_ASAP7_75t_R _30417_ (.A1(ld),
    .A2(text_in[26]),
    .B(_07792_),
    .Y(_01454_));
 NOR2x1_ASAP7_75t_R _30418_ (.A(ld),
    .B(_00539_),
    .Y(_07793_));
 AO21x1_ASAP7_75t_R _30419_ (.A1(ld),
    .A2(text_in[27]),
    .B(_07793_),
    .Y(_01455_));
 NOR2x1_ASAP7_75t_R _30420_ (.A(ld),
    .B(_00538_),
    .Y(_07794_));
 AO21x1_ASAP7_75t_R _30421_ (.A1(ld),
    .A2(text_in[28]),
    .B(_07794_),
    .Y(_01456_));
 NOR2x1_ASAP7_75t_R _30422_ (.A(ld),
    .B(_00537_),
    .Y(_07795_));
 AO21x1_ASAP7_75t_R _30423_ (.A1(ld),
    .A2(text_in[29]),
    .B(_07795_),
    .Y(_01457_));
 NOR2x1_ASAP7_75t_R _30425_ (.A(ld),
    .B(_00410_),
    .Y(_07797_));
 AO21x1_ASAP7_75t_R _30426_ (.A1(ld),
    .A2(text_in[2]),
    .B(_07797_),
    .Y(_01458_));
 NOR2x1_ASAP7_75t_R _30427_ (.A(ld),
    .B(_00536_),
    .Y(_07798_));
 AO21x1_ASAP7_75t_R _30428_ (.A1(ld),
    .A2(text_in[30]),
    .B(_07798_),
    .Y(_01459_));
 NOR2x1_ASAP7_75t_R _30430_ (.A(ld),
    .B(_00535_),
    .Y(_07800_));
 AO21x1_ASAP7_75t_R _30431_ (.A1(ld),
    .A2(text_in[31]),
    .B(_07800_),
    .Y(_01460_));
 NOR2x1_ASAP7_75t_R _30432_ (.A(ld),
    .B(_00406_),
    .Y(_07801_));
 AO21x1_ASAP7_75t_R _30433_ (.A1(ld),
    .A2(text_in[32]),
    .B(_07801_),
    .Y(_01461_));
 NOR2x1_ASAP7_75t_R _30434_ (.A(ld),
    .B(_00405_),
    .Y(_07802_));
 AO21x1_ASAP7_75t_R _30435_ (.A1(ld),
    .A2(text_in[33]),
    .B(_07802_),
    .Y(_01462_));
 NOR2x1_ASAP7_75t_R _30436_ (.A(ld),
    .B(_00407_),
    .Y(_07803_));
 AO21x1_ASAP7_75t_R _30437_ (.A1(ld),
    .A2(text_in[34]),
    .B(_07803_),
    .Y(_01463_));
 NOR2x1_ASAP7_75t_R _30438_ (.A(ld),
    .B(_00534_),
    .Y(_07804_));
 AO21x1_ASAP7_75t_R _30439_ (.A1(ld),
    .A2(text_in[35]),
    .B(_07804_),
    .Y(_01464_));
 NOR2x1_ASAP7_75t_R _30440_ (.A(ld),
    .B(_00533_),
    .Y(_07805_));
 AO21x1_ASAP7_75t_R _30441_ (.A1(ld),
    .A2(text_in[36]),
    .B(_07805_),
    .Y(_01465_));
 NOR2x1_ASAP7_75t_R _30442_ (.A(ld),
    .B(_00532_),
    .Y(_07806_));
 AO21x1_ASAP7_75t_R _30443_ (.A1(ld),
    .A2(text_in[37]),
    .B(_07806_),
    .Y(_01466_));
 NOR2x1_ASAP7_75t_R _30444_ (.A(ld),
    .B(_00531_),
    .Y(_07807_));
 AO21x1_ASAP7_75t_R _30445_ (.A1(ld),
    .A2(text_in[38]),
    .B(_07807_),
    .Y(_01467_));
 NOR2x1_ASAP7_75t_R _30447_ (.A(ld),
    .B(_00530_),
    .Y(_07809_));
 AO21x1_ASAP7_75t_R _30448_ (.A1(ld),
    .A2(text_in[39]),
    .B(_07809_),
    .Y(_01468_));
 NOR2x1_ASAP7_75t_R _30449_ (.A(ld),
    .B(_00529_),
    .Y(_07810_));
 AO21x1_ASAP7_75t_R _30450_ (.A1(ld),
    .A2(text_in[3]),
    .B(_07810_),
    .Y(_01469_));
 NOR2x1_ASAP7_75t_R _30452_ (.A(ld),
    .B(_00475_),
    .Y(_07812_));
 AO21x1_ASAP7_75t_R _30453_ (.A1(ld),
    .A2(text_in[40]),
    .B(_07812_),
    .Y(_01470_));
 NOR2x1_ASAP7_75t_R _30454_ (.A(ld),
    .B(_00474_),
    .Y(_07813_));
 AO21x1_ASAP7_75t_R _30455_ (.A1(ld),
    .A2(text_in[41]),
    .B(_07813_),
    .Y(_01471_));
 NOR2x1_ASAP7_75t_R _30456_ (.A(ld),
    .B(_00476_),
    .Y(_07814_));
 AO21x1_ASAP7_75t_R _30457_ (.A1(ld),
    .A2(text_in[42]),
    .B(_07814_),
    .Y(_01472_));
 NOR2x1_ASAP7_75t_R _30458_ (.A(ld),
    .B(_00528_),
    .Y(_07815_));
 AO21x1_ASAP7_75t_R _30459_ (.A1(ld),
    .A2(text_in[43]),
    .B(_07815_),
    .Y(_01473_));
 NOR2x1_ASAP7_75t_R _30460_ (.A(ld),
    .B(_00527_),
    .Y(_07816_));
 AO21x1_ASAP7_75t_R _30461_ (.A1(ld),
    .A2(text_in[44]),
    .B(_07816_),
    .Y(_01474_));
 NOR2x1_ASAP7_75t_R _30462_ (.A(ld),
    .B(_00526_),
    .Y(_07817_));
 AO21x1_ASAP7_75t_R _30463_ (.A1(ld),
    .A2(text_in[45]),
    .B(_07817_),
    .Y(_01475_));
 NOR2x1_ASAP7_75t_R _30464_ (.A(ld),
    .B(_00525_),
    .Y(_07818_));
 AO21x1_ASAP7_75t_R _30465_ (.A1(ld),
    .A2(text_in[46]),
    .B(_07818_),
    .Y(_01476_));
 NOR2x1_ASAP7_75t_R _30466_ (.A(ld),
    .B(_00524_),
    .Y(_07819_));
 AO21x1_ASAP7_75t_R _30467_ (.A1(ld),
    .A2(text_in[47]),
    .B(_07819_),
    .Y(_01477_));
 NOR2x1_ASAP7_75t_R _30469_ (.A(ld),
    .B(_00463_),
    .Y(_07821_));
 AO21x1_ASAP7_75t_R _30470_ (.A1(ld),
    .A2(text_in[48]),
    .B(_07821_),
    .Y(_01478_));
 NOR2x1_ASAP7_75t_R _30471_ (.A(ld),
    .B(_00462_),
    .Y(_07822_));
 AO21x1_ASAP7_75t_R _30472_ (.A1(ld),
    .A2(text_in[49]),
    .B(_07822_),
    .Y(_01479_));
 NOR2x1_ASAP7_75t_R _30474_ (.A(ld),
    .B(_00523_),
    .Y(_07824_));
 AO21x1_ASAP7_75t_R _30475_ (.A1(ld),
    .A2(text_in[4]),
    .B(_07824_),
    .Y(_01480_));
 NOR2x1_ASAP7_75t_R _30476_ (.A(ld),
    .B(_00464_),
    .Y(_07825_));
 AO21x1_ASAP7_75t_R _30477_ (.A1(ld),
    .A2(text_in[50]),
    .B(_07825_),
    .Y(_01481_));
 NOR2x1_ASAP7_75t_R _30478_ (.A(ld),
    .B(_00522_),
    .Y(_07826_));
 AO21x1_ASAP7_75t_R _30479_ (.A1(ld),
    .A2(text_in[51]),
    .B(_07826_),
    .Y(_01482_));
 NOR2x1_ASAP7_75t_R _30480_ (.A(ld),
    .B(_00521_),
    .Y(_07827_));
 AO21x1_ASAP7_75t_R _30481_ (.A1(ld),
    .A2(text_in[52]),
    .B(_07827_),
    .Y(_01483_));
 NOR2x1_ASAP7_75t_R _30482_ (.A(ld),
    .B(_00520_),
    .Y(_07828_));
 AO21x1_ASAP7_75t_R _30483_ (.A1(ld),
    .A2(text_in[53]),
    .B(_07828_),
    .Y(_01484_));
 NOR2x1_ASAP7_75t_R _30484_ (.A(ld),
    .B(_00519_),
    .Y(_07829_));
 AO21x1_ASAP7_75t_R _30485_ (.A1(ld),
    .A2(text_in[54]),
    .B(_07829_),
    .Y(_01485_));
 NOR2x1_ASAP7_75t_R _30486_ (.A(ld),
    .B(_00518_),
    .Y(_07830_));
 AO21x1_ASAP7_75t_R _30487_ (.A1(ld),
    .A2(text_in[55]),
    .B(_07830_),
    .Y(_01486_));
 NOR2x1_ASAP7_75t_R _30488_ (.A(ld),
    .B(_00451_),
    .Y(_07831_));
 AO21x1_ASAP7_75t_R _30489_ (.A1(ld),
    .A2(text_in[56]),
    .B(_07831_),
    .Y(_01487_));
 NOR2x1_ASAP7_75t_R _30491_ (.A(ld),
    .B(_00450_),
    .Y(_07833_));
 AO21x1_ASAP7_75t_R _30492_ (.A1(ld),
    .A2(text_in[57]),
    .B(_07833_),
    .Y(_01488_));
 NOR2x1_ASAP7_75t_R _30493_ (.A(ld),
    .B(_00452_),
    .Y(_07834_));
 AO21x1_ASAP7_75t_R _30494_ (.A1(ld),
    .A2(text_in[58]),
    .B(_07834_),
    .Y(_01489_));
 NOR2x1_ASAP7_75t_R _30496_ (.A(ld),
    .B(_00517_),
    .Y(_07836_));
 AO21x1_ASAP7_75t_R _30497_ (.A1(ld),
    .A2(text_in[59]),
    .B(_07836_),
    .Y(_01490_));
 NOR2x1_ASAP7_75t_R _30498_ (.A(ld),
    .B(_00516_),
    .Y(_07837_));
 AO21x1_ASAP7_75t_R _30499_ (.A1(ld),
    .A2(text_in[5]),
    .B(_07837_),
    .Y(_01491_));
 NOR2x1_ASAP7_75t_R _30500_ (.A(ld),
    .B(_00515_),
    .Y(_07838_));
 AO21x1_ASAP7_75t_R _30501_ (.A1(ld),
    .A2(text_in[60]),
    .B(_07838_),
    .Y(_01492_));
 NOR2x1_ASAP7_75t_R _30502_ (.A(ld),
    .B(_00514_),
    .Y(_07839_));
 AO21x1_ASAP7_75t_R _30503_ (.A1(ld),
    .A2(text_in[61]),
    .B(_07839_),
    .Y(_01493_));
 NOR2x1_ASAP7_75t_R _30504_ (.A(ld),
    .B(_00513_),
    .Y(_07840_));
 AO21x1_ASAP7_75t_R _30505_ (.A1(ld),
    .A2(text_in[62]),
    .B(_07840_),
    .Y(_01494_));
 NOR2x1_ASAP7_75t_R _30506_ (.A(ld),
    .B(_00512_),
    .Y(_07841_));
 AO21x1_ASAP7_75t_R _30507_ (.A1(ld),
    .A2(text_in[63]),
    .B(_07841_),
    .Y(_01495_));
 NOR2x1_ASAP7_75t_R _30508_ (.A(ld),
    .B(_00484_),
    .Y(_07842_));
 AO21x1_ASAP7_75t_R _30509_ (.A1(ld),
    .A2(text_in[64]),
    .B(_07842_),
    .Y(_01496_));
 NOR2x1_ASAP7_75t_R _30510_ (.A(ld),
    .B(_00483_),
    .Y(_07843_));
 AO21x1_ASAP7_75t_R _30511_ (.A1(ld),
    .A2(text_in[65]),
    .B(_07843_),
    .Y(_01497_));
 NOR2x1_ASAP7_75t_R _30513_ (.A(ld),
    .B(_00485_),
    .Y(_07845_));
 AO21x1_ASAP7_75t_R _30514_ (.A1(ld),
    .A2(text_in[66]),
    .B(_07845_),
    .Y(_01498_));
 NOR2x1_ASAP7_75t_R _30515_ (.A(ld),
    .B(_00511_),
    .Y(_07846_));
 AO21x1_ASAP7_75t_R _30516_ (.A1(ld),
    .A2(text_in[67]),
    .B(_07846_),
    .Y(_01499_));
 NOR2x1_ASAP7_75t_R _30518_ (.A(ld),
    .B(_00510_),
    .Y(_07848_));
 AO21x1_ASAP7_75t_R _30519_ (.A1(ld),
    .A2(text_in[68]),
    .B(_07848_),
    .Y(_01500_));
 NOR2x1_ASAP7_75t_R _30520_ (.A(ld),
    .B(_00509_),
    .Y(_07849_));
 AO21x1_ASAP7_75t_R _30521_ (.A1(ld),
    .A2(text_in[69]),
    .B(_07849_),
    .Y(_01501_));
 NOR2x1_ASAP7_75t_R _30522_ (.A(ld),
    .B(_00508_),
    .Y(_07850_));
 AO21x1_ASAP7_75t_R _30523_ (.A1(ld),
    .A2(text_in[6]),
    .B(_07850_),
    .Y(_01502_));
 NOR2x1_ASAP7_75t_R _30524_ (.A(ld),
    .B(_00507_),
    .Y(_07851_));
 AO21x1_ASAP7_75t_R _30525_ (.A1(ld),
    .A2(text_in[70]),
    .B(_07851_),
    .Y(_01503_));
 NOR2x1_ASAP7_75t_R _30526_ (.A(ld),
    .B(_00506_),
    .Y(_07852_));
 AO21x1_ASAP7_75t_R _30527_ (.A1(ld),
    .A2(text_in[71]),
    .B(_07852_),
    .Y(_01504_));
 NOR2x1_ASAP7_75t_R _30528_ (.A(ld),
    .B(_00472_),
    .Y(_07853_));
 AO21x1_ASAP7_75t_R _30529_ (.A1(ld),
    .A2(text_in[72]),
    .B(_07853_),
    .Y(_01505_));
 NOR2x1_ASAP7_75t_R _30530_ (.A(ld),
    .B(_00471_),
    .Y(_07854_));
 AO21x1_ASAP7_75t_R _30531_ (.A1(ld),
    .A2(text_in[73]),
    .B(_07854_),
    .Y(_01506_));
 NOR2x1_ASAP7_75t_R _30532_ (.A(ld),
    .B(_00473_),
    .Y(_07855_));
 AO21x1_ASAP7_75t_R _30533_ (.A1(ld),
    .A2(text_in[74]),
    .B(_07855_),
    .Y(_01507_));
 NOR2x1_ASAP7_75t_R _30535_ (.A(ld),
    .B(_00505_),
    .Y(_07857_));
 AO21x1_ASAP7_75t_R _30536_ (.A1(ld),
    .A2(text_in[75]),
    .B(_07857_),
    .Y(_01508_));
 NOR2x1_ASAP7_75t_R _30537_ (.A(ld),
    .B(_00504_),
    .Y(_07858_));
 AO21x1_ASAP7_75t_R _30538_ (.A1(ld),
    .A2(text_in[76]),
    .B(_07858_),
    .Y(_01509_));
 NOR2x1_ASAP7_75t_R _30540_ (.A(ld),
    .B(_00503_),
    .Y(_07860_));
 AO21x1_ASAP7_75t_R _30541_ (.A1(ld),
    .A2(text_in[77]),
    .B(_07860_),
    .Y(_01510_));
 NOR2x1_ASAP7_75t_R _30542_ (.A(ld),
    .B(_00502_),
    .Y(_07861_));
 AO21x1_ASAP7_75t_R _30543_ (.A1(ld),
    .A2(text_in[78]),
    .B(_07861_),
    .Y(_01511_));
 NOR2x1_ASAP7_75t_R _30544_ (.A(ld),
    .B(_00501_),
    .Y(_07862_));
 AO21x1_ASAP7_75t_R _30545_ (.A1(ld),
    .A2(text_in[79]),
    .B(_07862_),
    .Y(_01512_));
 NOR2x1_ASAP7_75t_R _30546_ (.A(ld),
    .B(_00500_),
    .Y(_07863_));
 AO21x1_ASAP7_75t_R _30547_ (.A1(ld),
    .A2(text_in[7]),
    .B(_07863_),
    .Y(_01513_));
 NOR2x1_ASAP7_75t_R _30548_ (.A(ld),
    .B(_00460_),
    .Y(_07864_));
 AO21x1_ASAP7_75t_R _30549_ (.A1(ld),
    .A2(text_in[80]),
    .B(_07864_),
    .Y(_01514_));
 NOR2x1_ASAP7_75t_R _30550_ (.A(ld),
    .B(_00459_),
    .Y(_07865_));
 AO21x1_ASAP7_75t_R _30551_ (.A1(ld),
    .A2(text_in[81]),
    .B(_07865_),
    .Y(_01515_));
 NOR2x1_ASAP7_75t_R _30552_ (.A(ld),
    .B(_00461_),
    .Y(_07866_));
 AO21x1_ASAP7_75t_R _30553_ (.A1(ld),
    .A2(text_in[82]),
    .B(_07866_),
    .Y(_01516_));
 NOR2x1_ASAP7_75t_R _30554_ (.A(ld),
    .B(_00499_),
    .Y(_07867_));
 AO21x1_ASAP7_75t_R _30555_ (.A1(ld),
    .A2(text_in[83]),
    .B(_07867_),
    .Y(_01517_));
 NOR2x1_ASAP7_75t_R _30557_ (.A(ld),
    .B(_00498_),
    .Y(_07869_));
 AO21x1_ASAP7_75t_R _30558_ (.A1(ld),
    .A2(text_in[84]),
    .B(_07869_),
    .Y(_01518_));
 NOR2x1_ASAP7_75t_R _30559_ (.A(ld),
    .B(_00497_),
    .Y(_07870_));
 AO21x1_ASAP7_75t_R _30560_ (.A1(ld),
    .A2(text_in[85]),
    .B(_07870_),
    .Y(_01519_));
 NOR2x1_ASAP7_75t_R _30562_ (.A(ld),
    .B(_00496_),
    .Y(_07872_));
 AO21x1_ASAP7_75t_R _30563_ (.A1(ld),
    .A2(text_in[86]),
    .B(_07872_),
    .Y(_01520_));
 NOR2x1_ASAP7_75t_R _30564_ (.A(ld),
    .B(_00495_),
    .Y(_07873_));
 AO21x1_ASAP7_75t_R _30565_ (.A1(ld),
    .A2(text_in[87]),
    .B(_07873_),
    .Y(_01521_));
 NOR2x1_ASAP7_75t_R _30566_ (.A(ld),
    .B(_00448_),
    .Y(_07874_));
 AO21x1_ASAP7_75t_R _30567_ (.A1(ld),
    .A2(text_in[88]),
    .B(_07874_),
    .Y(_01522_));
 NOR2x1_ASAP7_75t_R _30568_ (.A(ld),
    .B(_00447_),
    .Y(_07875_));
 AO21x1_ASAP7_75t_R _30569_ (.A1(ld),
    .A2(text_in[89]),
    .B(_07875_),
    .Y(_01523_));
 NOR2x1_ASAP7_75t_R _30570_ (.A(ld),
    .B(_00478_),
    .Y(_07876_));
 AO21x1_ASAP7_75t_R _30571_ (.A1(ld),
    .A2(text_in[8]),
    .B(_07876_),
    .Y(_01524_));
 NOR2x1_ASAP7_75t_R _30572_ (.A(ld),
    .B(_00449_),
    .Y(_07877_));
 AO21x1_ASAP7_75t_R _30573_ (.A1(ld),
    .A2(text_in[90]),
    .B(_07877_),
    .Y(_01525_));
 NOR2x1_ASAP7_75t_R _30574_ (.A(ld),
    .B(_00494_),
    .Y(_07878_));
 AO21x1_ASAP7_75t_R _30575_ (.A1(ld),
    .A2(text_in[91]),
    .B(_07878_),
    .Y(_01526_));
 NOR2x1_ASAP7_75t_R _30576_ (.A(ld),
    .B(_00493_),
    .Y(_07879_));
 AO21x1_ASAP7_75t_R _30577_ (.A1(ld),
    .A2(text_in[92]),
    .B(_07879_),
    .Y(_01527_));
 NOR2x1_ASAP7_75t_R _30578_ (.A(ld),
    .B(_00492_),
    .Y(_07880_));
 AO21x1_ASAP7_75t_R _30579_ (.A1(ld),
    .A2(text_in[93]),
    .B(_07880_),
    .Y(_01528_));
 NOR2x1_ASAP7_75t_R _30580_ (.A(ld),
    .B(_00491_),
    .Y(_07881_));
 AO21x1_ASAP7_75t_R _30581_ (.A1(ld),
    .A2(text_in[94]),
    .B(_07881_),
    .Y(_01529_));
 NOR2x1_ASAP7_75t_R _30582_ (.A(ld),
    .B(_00490_),
    .Y(_07882_));
 AO21x1_ASAP7_75t_R _30583_ (.A1(ld),
    .A2(text_in[95]),
    .B(_07882_),
    .Y(_01530_));
 NOR2x1_ASAP7_75t_R _30584_ (.A(ld),
    .B(_00481_),
    .Y(_07883_));
 AO21x1_ASAP7_75t_R _30585_ (.A1(ld),
    .A2(text_in[96]),
    .B(_07883_),
    .Y(_01531_));
 NOR2x1_ASAP7_75t_R _30586_ (.A(ld),
    .B(_00480_),
    .Y(_07884_));
 AO21x1_ASAP7_75t_R _30587_ (.A1(ld),
    .A2(text_in[97]),
    .B(_07884_),
    .Y(_01532_));
 NOR2x1_ASAP7_75t_R _30588_ (.A(ld),
    .B(_00482_),
    .Y(_07885_));
 AO21x1_ASAP7_75t_R _30589_ (.A1(ld),
    .A2(text_in[98]),
    .B(_07885_),
    .Y(_01533_));
 NOR2x1_ASAP7_75t_R _30590_ (.A(ld),
    .B(_00489_),
    .Y(_07886_));
 AO21x1_ASAP7_75t_R _30591_ (.A1(ld),
    .A2(text_in[99]),
    .B(_07886_),
    .Y(_01534_));
 NOR2x1_ASAP7_75t_R _30592_ (.A(ld),
    .B(_00477_),
    .Y(_07887_));
 AO21x1_ASAP7_75t_R _30593_ (.A1(ld),
    .A2(text_in[9]),
    .B(_07887_),
    .Y(_01535_));
 AND3x1_ASAP7_75t_R _30594_ (.A(_00570_),
    .B(_00571_),
    .C(_00572_),
    .Y(_07888_));
 AOI21x1_ASAP7_75t_R _30595_ (.A1(_00571_),
    .A2(_00572_),
    .B(_00570_),
    .Y(_07889_));
 INVx1_ASAP7_75t_R _30596_ (.A(rst),
    .Y(_07890_));
 AOI21x1_ASAP7_75t_R _30597_ (.A1(_00411_),
    .A2(_07888_),
    .B(_07890_),
    .Y(_07891_));
 OA211x2_ASAP7_75t_R _30598_ (.A1(_07888_),
    .A2(_07889_),
    .B(_07891_),
    .C(_08005_),
    .Y(_01406_));
 XNOR2x2_ASAP7_75t_R _30599_ (.A(_00487_),
    .B(_00971_),
    .Y(_07892_));
 INVx1_ASAP7_75t_R _30600_ (.A(_00970_),
    .Y(_07893_));
 AO21x1_ASAP7_75t_R _30601_ (.A1(_07892_),
    .A2(_07893_),
    .B(ld),
    .Y(_01536_));
 OR3x1_ASAP7_75t_R _30602_ (.A(_00487_),
    .B(_00965_),
    .C(\u0.r0.rcnt_next[0] ),
    .Y(_07894_));
 XOR2x2_ASAP7_75t_R _30603_ (.A(_07894_),
    .B(_00829_),
    .Y(_07895_));
 INVx1_ASAP7_75t_R _30604_ (.A(_07892_),
    .Y(_07896_));
 OR3x1_ASAP7_75t_R _30605_ (.A(_07895_),
    .B(_00966_),
    .C(_07896_),
    .Y(_07897_));
 INVx1_ASAP7_75t_R _30606_ (.A(_07895_),
    .Y(_07898_));
 INVx1_ASAP7_75t_R _30607_ (.A(_00967_),
    .Y(_07899_));
 OR3x1_ASAP7_75t_R _30608_ (.A(_07898_),
    .B(_07899_),
    .C(_07896_),
    .Y(_07900_));
 AOI21x1_ASAP7_75t_R _30609_ (.A1(_07897_),
    .A2(_07900_),
    .B(ld),
    .Y(_01537_));
 OR3x1_ASAP7_75t_R _30610_ (.A(_07895_),
    .B(_00969_),
    .C(_07896_),
    .Y(_07901_));
 OR3x1_ASAP7_75t_R _30611_ (.A(_07898_),
    .B(_00966_),
    .C(_07896_),
    .Y(_07902_));
 AOI21x1_ASAP7_75t_R _30612_ (.A1(_07901_),
    .A2(_07902_),
    .B(ld),
    .Y(_01538_));
 OR3x1_ASAP7_75t_R _30613_ (.A(_07895_),
    .B(_00968_),
    .C(_07896_),
    .Y(_07903_));
 OR3x1_ASAP7_75t_R _30614_ (.A(_07898_),
    .B(_00970_),
    .C(_07896_),
    .Y(_07904_));
 AOI21x1_ASAP7_75t_R _30615_ (.A1(_07903_),
    .A2(_07904_),
    .B(ld),
    .Y(_01539_));
 OR3x1_ASAP7_75t_R _30616_ (.A(_07895_),
    .B(_00970_),
    .C(_07892_),
    .Y(_07905_));
 AOI21x1_ASAP7_75t_R _30617_ (.A1(_07905_),
    .A2(_07900_),
    .B(ld),
    .Y(_01540_));
 OR3x1_ASAP7_75t_R _30618_ (.A(_07895_),
    .B(_00966_),
    .C(_07892_),
    .Y(_07906_));
 AOI21x1_ASAP7_75t_R _30619_ (.A1(_07906_),
    .A2(_07902_),
    .B(ld),
    .Y(_01541_));
 NOR2x1_ASAP7_75t_R _30620_ (.A(ld),
    .B(_07892_),
    .Y(_01546_));
 NAND2x1_ASAP7_75t_R _30621_ (.A(_01546_),
    .B(_07898_),
    .Y(_07907_));
 NOR2x1_ASAP7_75t_R _30622_ (.A(_00969_),
    .B(_07907_),
    .Y(_01542_));
 NOR2x1_ASAP7_75t_R _30623_ (.A(_00968_),
    .B(_07907_),
    .Y(_01543_));
 NOR2x1_ASAP7_75t_R _30624_ (.A(ld),
    .B(\u0.r0.rcnt[0] ),
    .Y(_01544_));
 NOR2x1_ASAP7_75t_R _30625_ (.A(ld),
    .B(_00967_),
    .Y(_01545_));
 AND2x2_ASAP7_75t_R _30626_ (.A(_07895_),
    .B(_08005_),
    .Y(_01547_));
 AO22x1_ASAP7_75t_R _30627_ (.A1(_07891_),
    .A2(_00572_),
    .B1(ld),
    .B2(rst),
    .Y(_01404_));
 OA21x2_ASAP7_75t_R _30628_ (.A1(_00571_),
    .A2(_00572_),
    .B(_08005_),
    .Y(_07908_));
 NAND2x1_ASAP7_75t_R _30629_ (.A(_00571_),
    .B(_00572_),
    .Y(_07909_));
 AO21x1_ASAP7_75t_R _30630_ (.A1(_00411_),
    .A2(_00570_),
    .B(_07909_),
    .Y(_07910_));
 AOI21x1_ASAP7_75t_R _30631_ (.A1(_07908_),
    .A2(_07910_),
    .B(_07890_),
    .Y(_01405_));
 NOR2x1_ASAP7_75t_R _30632_ (.A(_00411_),
    .B(_07888_),
    .Y(_07911_));
 OA21x2_ASAP7_75t_R _30633_ (.A1(_07911_),
    .A2(ld),
    .B(rst),
    .Y(_01407_));
 HAxp5_ASAP7_75t_R _30634_ (.A(\u0.r0.rcnt_next[0] ),
    .B(_00965_),
    .CON(_00966_),
    .SN(_00967_));
 HAxp5_ASAP7_75t_R _30635_ (.A(\u0.r0.rcnt_next[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CON(_00968_),
    .SN(_15573_));
 HAxp5_ASAP7_75t_R _30636_ (.A(\u0.r0.rcnt[0] ),
    .B(_00965_),
    .CON(_00969_),
    .SN(_15574_));
 HAxp5_ASAP7_75t_R _30637_ (.A(\u0.r0.rcnt[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CON(_00970_),
    .SN(_15575_));
 HAxp5_ASAP7_75t_R _30638_ (.A(\u0.r0.rcnt[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CON(_00971_),
    .SN(_15576_));
 HAxp5_ASAP7_75t_SL _30639_ (.A(_00973_),
    .B(_00972_),
    .CON(_00974_),
    .SN(_00975_));
 HAxp5_ASAP7_75t_R _30640_ (.A(_00972_),
    .B(_00973_),
    .CON(_00976_),
    .SN(_15577_));
 HAxp5_ASAP7_75t_SL _30641_ (.A(_00972_),
    .B(_08045_),
    .CON(_00978_),
    .SN(_15578_));
 HAxp5_ASAP7_75t_SL _30642_ (.A(_00972_),
    .B(_08045_),
    .CON(_00979_),
    .SN(_15579_));
 HAxp5_ASAP7_75t_R _30643_ (.A(_08052_),
    .B(_00973_),
    .CON(_00981_),
    .SN(_15580_));
 HAxp5_ASAP7_75t_R _30644_ (.A(_08052_),
    .B(_00973_),
    .CON(_00982_),
    .SN(_15581_));
 HAxp5_ASAP7_75t_R _30645_ (.A(_08052_),
    .B(_08045_),
    .CON(_00983_),
    .SN(_15582_));
 HAxp5_ASAP7_75t_R _30646_ (.A(_08052_),
    .B(_08045_),
    .CON(_00984_),
    .SN(_15583_));
 HAxp5_ASAP7_75t_SL _30647_ (.A(_00972_),
    .B(_08063_),
    .CON(_00986_),
    .SN(_00987_));
 HAxp5_ASAP7_75t_R _30648_ (.A(_00972_),
    .B(_08063_),
    .CON(_00988_),
    .SN(_15584_));
 HAxp5_ASAP7_75t_R _30649_ (.A(_00972_),
    .B(_00989_),
    .CON(_00990_),
    .SN(_15585_));
 HAxp5_ASAP7_75t_SL _30650_ (.A(_00972_),
    .B(_00989_),
    .CON(_00991_),
    .SN(_15586_));
 HAxp5_ASAP7_75t_R _30651_ (.A(_08052_),
    .B(_08063_),
    .CON(_00992_),
    .SN(_15587_));
 HAxp5_ASAP7_75t_R _30652_ (.A(_08052_),
    .B(_08063_),
    .CON(_00993_),
    .SN(_15588_));
 HAxp5_ASAP7_75t_SL _30653_ (.A(_08995_),
    .B(_00994_),
    .CON(_00996_),
    .SN(_00997_));
 HAxp5_ASAP7_75t_SL _30654_ (.A(_00994_),
    .B(_08995_),
    .CON(_00998_),
    .SN(_15589_));
 HAxp5_ASAP7_75t_L _30655_ (.A(_00994_),
    .B(_08907_),
    .CON(_01000_),
    .SN(_15590_));
 HAxp5_ASAP7_75t_L _30656_ (.A(_00994_),
    .B(_08907_),
    .CON(_01001_),
    .SN(_15591_));
 HAxp5_ASAP7_75t_SL _30657_ (.A(_01002_),
    .B(_08995_),
    .CON(_01003_),
    .SN(_15592_));
 HAxp5_ASAP7_75t_R _30658_ (.A(_01002_),
    .B(_08995_),
    .CON(_01004_),
    .SN(_15593_));
 HAxp5_ASAP7_75t_L _30659_ (.A(_01002_),
    .B(_08907_),
    .CON(_01005_),
    .SN(_15594_));
 HAxp5_ASAP7_75t_R _30660_ (.A(_01002_),
    .B(_08907_),
    .CON(_01006_),
    .SN(_15595_));
 HAxp5_ASAP7_75t_R _30661_ (.A(_00994_),
    .B(_08918_),
    .CON(_01008_),
    .SN(_01009_));
 HAxp5_ASAP7_75t_SL _30662_ (.A(_00994_),
    .B(_08918_),
    .CON(_01010_),
    .SN(_15596_));
 HAxp5_ASAP7_75t_R _30663_ (.A(_00994_),
    .B(_08919_),
    .CON(_01012_),
    .SN(_15597_));
 HAxp5_ASAP7_75t_R _30664_ (.A(_00994_),
    .B(_08919_),
    .CON(_01013_),
    .SN(_15598_));
 HAxp5_ASAP7_75t_R _30665_ (.A(_01002_),
    .B(_08918_),
    .CON(_01014_),
    .SN(_15599_));
 HAxp5_ASAP7_75t_R _30666_ (.A(_01002_),
    .B(_08918_),
    .CON(_01015_),
    .SN(_15600_));
 HAxp5_ASAP7_75t_SL _30667_ (.A(_09557_),
    .B(_09554_),
    .CON(_01018_),
    .SN(_01019_));
 HAxp5_ASAP7_75t_L _30668_ (.A(_09554_),
    .B(_09557_),
    .CON(_01020_),
    .SN(_15601_));
 HAxp5_ASAP7_75t_L _30669_ (.A(_09554_),
    .B(_08866_),
    .CON(_01022_),
    .SN(_15602_));
 HAxp5_ASAP7_75t_SL _30670_ (.A(_08866_),
    .B(_09554_),
    .CON(_01023_),
    .SN(_15603_));
 HAxp5_ASAP7_75t_SL _30671_ (.A(_09557_),
    .B(_08871_),
    .CON(_01025_),
    .SN(_15604_));
 HAxp5_ASAP7_75t_L _30672_ (.A(_08871_),
    .B(_09557_),
    .CON(_01026_),
    .SN(_15605_));
 HAxp5_ASAP7_75t_L _30673_ (.A(_08871_),
    .B(_08866_),
    .CON(_01027_),
    .SN(_15606_));
 HAxp5_ASAP7_75t_R _30674_ (.A(_08871_),
    .B(_08866_),
    .CON(_01028_),
    .SN(_15607_));
 HAxp5_ASAP7_75t_SL _30675_ (.A(_09554_),
    .B(_08878_),
    .CON(_01030_),
    .SN(_01031_));
 HAxp5_ASAP7_75t_R _30676_ (.A(_09554_),
    .B(_08878_),
    .CON(_01032_),
    .SN(_15608_));
 HAxp5_ASAP7_75t_R _30677_ (.A(_09554_),
    .B(_08879_),
    .CON(_01034_),
    .SN(_15609_));
 HAxp5_ASAP7_75t_R _30678_ (.A(_09554_),
    .B(_08879_),
    .CON(_01035_),
    .SN(_15610_));
 HAxp5_ASAP7_75t_R _30679_ (.A(_08871_),
    .B(_08878_),
    .CON(_01036_),
    .SN(_15611_));
 HAxp5_ASAP7_75t_R _30680_ (.A(_08871_),
    .B(_08878_),
    .CON(_01037_),
    .SN(_15612_));
 HAxp5_ASAP7_75t_SL _30681_ (.A(_10110_),
    .B(_10103_),
    .CON(_01040_),
    .SN(_01041_));
 HAxp5_ASAP7_75t_L _30682_ (.A(_10103_),
    .B(_10110_),
    .CON(_01042_),
    .SN(_15613_));
 HAxp5_ASAP7_75t_SL _30683_ (.A(_01043_),
    .B(_10103_),
    .CON(_01044_),
    .SN(_15614_));
 HAxp5_ASAP7_75t_L _30684_ (.A(_10103_),
    .B(_01043_),
    .CON(_01045_),
    .SN(_15615_));
 HAxp5_ASAP7_75t_SL _30685_ (.A(_10110_),
    .B(_01046_),
    .CON(_01047_),
    .SN(_15616_));
 HAxp5_ASAP7_75t_SL _30686_ (.A(_10110_),
    .B(_01046_),
    .CON(_01048_),
    .SN(_15617_));
 HAxp5_ASAP7_75t_L _30687_ (.A(_01046_),
    .B(_01043_),
    .CON(_01049_),
    .SN(_15618_));
 HAxp5_ASAP7_75t_L _30688_ (.A(_01046_),
    .B(_01043_),
    .CON(_01050_),
    .SN(_15619_));
 HAxp5_ASAP7_75t_R _30689_ (.A(_10104_),
    .B(_10103_),
    .CON(_01052_),
    .SN(_01053_));
 HAxp5_ASAP7_75t_R _30690_ (.A(_10104_),
    .B(_10103_),
    .CON(_01054_),
    .SN(_15620_));
 HAxp5_ASAP7_75t_R _30691_ (.A(_08958_),
    .B(_10103_),
    .CON(_01056_),
    .SN(_15621_));
 HAxp5_ASAP7_75t_R _30692_ (.A(_08958_),
    .B(_10103_),
    .CON(_01057_),
    .SN(_15622_));
 HAxp5_ASAP7_75t_R _30693_ (.A(_08958_),
    .B(_01046_),
    .CON(_01058_),
    .SN(_15623_));
 HAxp5_ASAP7_75t_R _30694_ (.A(_08958_),
    .B(_01046_),
    .CON(_01059_),
    .SN(_15624_));
 HAxp5_ASAP7_75t_SL _30695_ (.A(_01061_),
    .B(_10723_),
    .CON(_01062_),
    .SN(_01063_));
 HAxp5_ASAP7_75t_SL _30696_ (.A(_10723_),
    .B(_01061_),
    .CON(_01064_),
    .SN(_15625_));
 HAxp5_ASAP7_75t_SL _30697_ (.A(_10687_),
    .B(_10723_),
    .CON(_01066_),
    .SN(_15626_));
 HAxp5_ASAP7_75t_SL _30698_ (.A(_01067_),
    .B(_01061_),
    .CON(_01068_),
    .SN(_15627_));
 HAxp5_ASAP7_75t_R _30699_ (.A(_01067_),
    .B(_01061_),
    .CON(_01069_),
    .SN(_15628_));
 HAxp5_ASAP7_75t_SL _30700_ (.A(_01067_),
    .B(_10687_),
    .CON(_01070_),
    .SN(_15629_));
 HAxp5_ASAP7_75t_L _30701_ (.A(_01067_),
    .B(_10687_),
    .CON(_01071_),
    .SN(_15630_));
 HAxp5_ASAP7_75t_R _30702_ (.A(_10728_),
    .B(_01061_),
    .CON(_01073_),
    .SN(_01074_));
 HAxp5_ASAP7_75t_R _30703_ (.A(_10728_),
    .B(_10687_),
    .CON(_01075_),
    .SN(_15631_));
 HAxp5_ASAP7_75t_R _30704_ (.A(_10728_),
    .B(_10687_),
    .CON(_01076_),
    .SN(_15632_));
 HAxp5_ASAP7_75t_SL _30705_ (.A(_10721_),
    .B(_01061_),
    .CON(_01078_),
    .SN(_15633_));
 HAxp5_ASAP7_75t_SL _30706_ (.A(_10721_),
    .B(_01061_),
    .CON(_01079_),
    .SN(_15634_));
 HAxp5_ASAP7_75t_SL _30707_ (.A(_10721_),
    .B(_10687_),
    .CON(_01080_),
    .SN(_15635_));
 HAxp5_ASAP7_75t_SL _30708_ (.A(_01082_),
    .B(_11449_),
    .CON(_01083_),
    .SN(_01084_));
 HAxp5_ASAP7_75t_L _30709_ (.A(_11449_),
    .B(_01082_),
    .CON(_01085_),
    .SN(_15636_));
 HAxp5_ASAP7_75t_R _30710_ (.A(_11449_),
    .B(_11407_),
    .CON(_01087_),
    .SN(_15637_));
 HAxp5_ASAP7_75t_SL _30711_ (.A(_01088_),
    .B(_01082_),
    .CON(_01089_),
    .SN(_15638_));
 HAxp5_ASAP7_75t_SL _30712_ (.A(_01082_),
    .B(_01088_),
    .CON(_01090_),
    .SN(_15639_));
 HAxp5_ASAP7_75t_SL _30713_ (.A(_01088_),
    .B(_11407_),
    .CON(_01091_),
    .SN(_15640_));
 HAxp5_ASAP7_75t_L _30714_ (.A(_01088_),
    .B(_11407_),
    .CON(_01092_),
    .SN(_15641_));
 HAxp5_ASAP7_75t_R _30715_ (.A(_11452_),
    .B(_01082_),
    .CON(_01094_),
    .SN(_01095_));
 HAxp5_ASAP7_75t_R _30716_ (.A(_11452_),
    .B(_11407_),
    .CON(_01096_),
    .SN(_15642_));
 HAxp5_ASAP7_75t_R _30717_ (.A(_11452_),
    .B(_11407_),
    .CON(_01097_),
    .SN(_15643_));
 HAxp5_ASAP7_75t_SL _30718_ (.A(_11446_),
    .B(_01082_),
    .CON(_01099_),
    .SN(_15644_));
 HAxp5_ASAP7_75t_R _30719_ (.A(_11446_),
    .B(_01082_),
    .CON(_01100_),
    .SN(_15645_));
 HAxp5_ASAP7_75t_R _30720_ (.A(_11446_),
    .B(_11407_),
    .CON(_01101_),
    .SN(_15646_));
 HAxp5_ASAP7_75t_SL _30721_ (.A(_01103_),
    .B(_12136_),
    .CON(_01104_),
    .SN(_01105_));
 HAxp5_ASAP7_75t_R _30722_ (.A(_12136_),
    .B(_01103_),
    .CON(_01106_),
    .SN(_15647_));
 HAxp5_ASAP7_75t_R _30723_ (.A(_12136_),
    .B(_12096_),
    .CON(_01108_),
    .SN(_15648_));
 HAxp5_ASAP7_75t_SL _30724_ (.A(_12114_),
    .B(_01103_),
    .CON(_01110_),
    .SN(_15649_));
 HAxp5_ASAP7_75t_SL _30725_ (.A(_12114_),
    .B(_01103_),
    .CON(_01111_),
    .SN(_15650_));
 HAxp5_ASAP7_75t_SL _30726_ (.A(_12114_),
    .B(_12096_),
    .CON(_01112_),
    .SN(_15651_));
 HAxp5_ASAP7_75t_SL _30727_ (.A(_12114_),
    .B(_12096_),
    .CON(_01113_),
    .SN(_15652_));
 HAxp5_ASAP7_75t_SL _30728_ (.A(_12140_),
    .B(_01103_),
    .CON(_01115_),
    .SN(_01116_));
 HAxp5_ASAP7_75t_R _30729_ (.A(_12140_),
    .B(_12096_),
    .CON(_01117_),
    .SN(_15653_));
 HAxp5_ASAP7_75t_SL _30730_ (.A(_12140_),
    .B(_12096_),
    .CON(_01118_),
    .SN(_15654_));
 HAxp5_ASAP7_75t_SL _30731_ (.A(_12132_),
    .B(_01103_),
    .CON(_01120_),
    .SN(_15655_));
 HAxp5_ASAP7_75t_SL _30732_ (.A(_12132_),
    .B(_01103_),
    .CON(_01121_),
    .SN(_15656_));
 HAxp5_ASAP7_75t_R _30733_ (.A(_12132_),
    .B(_12096_),
    .CON(_01122_),
    .SN(_15657_));
 HAxp5_ASAP7_75t_SL _30734_ (.A(_01124_),
    .B(_01123_),
    .CON(_01125_),
    .SN(_01126_));
 HAxp5_ASAP7_75t_L _30735_ (.A(_01123_),
    .B(_01124_),
    .CON(_01127_),
    .SN(_15658_));
 HAxp5_ASAP7_75t_SL _30736_ (.A(_12785_),
    .B(_01123_),
    .CON(_01129_),
    .SN(_15659_));
 HAxp5_ASAP7_75t_SL _30737_ (.A(_01124_),
    .B(_12803_),
    .CON(_01131_),
    .SN(_15660_));
 HAxp5_ASAP7_75t_L _30738_ (.A(_12803_),
    .B(_01124_),
    .CON(_01132_),
    .SN(_15661_));
 HAxp5_ASAP7_75t_R _30739_ (.A(_12803_),
    .B(_12785_),
    .CON(_01133_),
    .SN(_15662_));
 HAxp5_ASAP7_75t_SL _30740_ (.A(_12785_),
    .B(_12803_),
    .CON(_01134_),
    .SN(_15663_));
 HAxp5_ASAP7_75t_R _30741_ (.A(_12826_),
    .B(_01124_),
    .CON(_01136_),
    .SN(_01137_));
 HAxp5_ASAP7_75t_R _30742_ (.A(_12826_),
    .B(_12785_),
    .CON(_01138_),
    .SN(_15664_));
 HAxp5_ASAP7_75t_R _30743_ (.A(_12826_),
    .B(_12785_),
    .CON(_01139_),
    .SN(_15665_));
 HAxp5_ASAP7_75t_SL _30744_ (.A(_12821_),
    .B(_01124_),
    .CON(_01141_),
    .SN(_15666_));
 HAxp5_ASAP7_75t_R _30745_ (.A(_12821_),
    .B(_01124_),
    .CON(_01142_),
    .SN(_15667_));
 HAxp5_ASAP7_75t_R _30746_ (.A(_12821_),
    .B(_12785_),
    .CON(_01143_),
    .SN(_15668_));
 HAxp5_ASAP7_75t_SL _30747_ (.A(_13537_),
    .B(_13510_),
    .CON(_01146_),
    .SN(_01147_));
 HAxp5_ASAP7_75t_R _30748_ (.A(_13510_),
    .B(_13537_),
    .CON(_01148_),
    .SN(_15669_));
 HAxp5_ASAP7_75t_R _30749_ (.A(_13510_),
    .B(_13471_),
    .CON(_01150_),
    .SN(_15670_));
 HAxp5_ASAP7_75t_SL _30750_ (.A(_13489_),
    .B(_13537_),
    .CON(_01152_),
    .SN(_15671_));
 HAxp5_ASAP7_75t_R _30751_ (.A(_13489_),
    .B(_13537_),
    .CON(_01153_),
    .SN(_15672_));
 HAxp5_ASAP7_75t_SL _30752_ (.A(_13489_),
    .B(_13471_),
    .CON(_01154_),
    .SN(_15673_));
 HAxp5_ASAP7_75t_SL _30753_ (.A(_13471_),
    .B(_13489_),
    .CON(_01155_),
    .SN(_15674_));
 HAxp5_ASAP7_75t_SL _30754_ (.A(_13513_),
    .B(_13537_),
    .CON(_01157_),
    .SN(_01158_));
 HAxp5_ASAP7_75t_SL _30755_ (.A(_13513_),
    .B(_13471_),
    .CON(_01159_),
    .SN(_15675_));
 HAxp5_ASAP7_75t_R _30756_ (.A(_13513_),
    .B(_13471_),
    .CON(_01160_),
    .SN(_15676_));
 HAxp5_ASAP7_75t_R _30757_ (.A(_13507_),
    .B(_13537_),
    .CON(_01162_),
    .SN(_15677_));
 HAxp5_ASAP7_75t_SL _30758_ (.A(_13507_),
    .B(_13537_),
    .CON(_01163_),
    .SN(_15678_));
 HAxp5_ASAP7_75t_SL _30759_ (.A(_13507_),
    .B(_13471_),
    .CON(_01164_),
    .SN(_15679_));
 HAxp5_ASAP7_75t_SL _30760_ (.A(_14308_),
    .B(_14227_),
    .CON(_01167_),
    .SN(_01168_));
 HAxp5_ASAP7_75t_SL _30761_ (.A(_14227_),
    .B(_14308_),
    .CON(_01169_),
    .SN(_15680_));
 HAxp5_ASAP7_75t_L _30762_ (.A(_14227_),
    .B(_14188_),
    .CON(_01171_),
    .SN(_15681_));
 HAxp5_ASAP7_75t_R _30763_ (.A(_14205_),
    .B(_14308_),
    .CON(_01173_),
    .SN(_15682_));
 HAxp5_ASAP7_75t_R _30764_ (.A(_14205_),
    .B(_14308_),
    .CON(_01174_),
    .SN(_15683_));
 HAxp5_ASAP7_75t_R _30765_ (.A(_14205_),
    .B(_14188_),
    .CON(_01175_),
    .SN(_15684_));
 HAxp5_ASAP7_75t_L _30766_ (.A(_14205_),
    .B(_14188_),
    .CON(_01176_),
    .SN(_15685_));
 HAxp5_ASAP7_75t_SL _30767_ (.A(_14230_),
    .B(_14308_),
    .CON(_01178_),
    .SN(_01179_));
 HAxp5_ASAP7_75t_SL _30768_ (.A(_14230_),
    .B(_14188_),
    .CON(_01180_),
    .SN(_15686_));
 HAxp5_ASAP7_75t_SL _30769_ (.A(_14230_),
    .B(_14188_),
    .CON(_01181_),
    .SN(_15687_));
 HAxp5_ASAP7_75t_SL _30770_ (.A(_14222_),
    .B(_14308_),
    .CON(_01183_),
    .SN(_15688_));
 HAxp5_ASAP7_75t_R _30771_ (.A(_14222_),
    .B(_14308_),
    .CON(_01184_),
    .SN(_15689_));
 HAxp5_ASAP7_75t_SL _30772_ (.A(_14222_),
    .B(_14188_),
    .CON(_01185_),
    .SN(_15690_));
 HAxp5_ASAP7_75t_SL _30773_ (.A(_01187_),
    .B(_01186_),
    .CON(_01188_),
    .SN(_01189_));
 HAxp5_ASAP7_75t_R _30774_ (.A(_01186_),
    .B(_01187_),
    .CON(_01190_),
    .SN(_15691_));
 HAxp5_ASAP7_75t_R _30775_ (.A(_01186_),
    .B(_14903_),
    .CON(_01192_),
    .SN(_15692_));
 HAxp5_ASAP7_75t_L _30776_ (.A(_01193_),
    .B(_01187_),
    .CON(_01194_),
    .SN(_15693_));
 HAxp5_ASAP7_75t_SL _30777_ (.A(_01193_),
    .B(_01187_),
    .CON(_01195_),
    .SN(_15694_));
 HAxp5_ASAP7_75t_R _30778_ (.A(_01193_),
    .B(_14903_),
    .CON(_01196_),
    .SN(_15695_));
 HAxp5_ASAP7_75t_SL _30779_ (.A(_14903_),
    .B(_01193_),
    .CON(_01197_),
    .SN(_15696_));
 HAxp5_ASAP7_75t_R _30780_ (.A(_14942_),
    .B(_01187_),
    .CON(_01199_),
    .SN(_01200_));
 HAxp5_ASAP7_75t_R _30781_ (.A(_14942_),
    .B(_14903_),
    .CON(_01201_),
    .SN(_15697_));
 HAxp5_ASAP7_75t_SL _30782_ (.A(_14942_),
    .B(_14903_),
    .CON(_01202_),
    .SN(_15698_));
 HAxp5_ASAP7_75t_R _30783_ (.A(_14937_),
    .B(_01187_),
    .CON(_01204_),
    .SN(_15699_));
 HAxp5_ASAP7_75t_R _30784_ (.A(_14937_),
    .B(_01187_),
    .CON(_01205_),
    .SN(_15700_));
 HAxp5_ASAP7_75t_R _30785_ (.A(_14937_),
    .B(_14903_),
    .CON(_01206_),
    .SN(_15701_));
 HAxp5_ASAP7_75t_SL _30786_ (.A(_01208_),
    .B(_01635_),
    .CON(_01209_),
    .SN(_01210_));
 HAxp5_ASAP7_75t_SL _30787_ (.A(_01635_),
    .B(_01208_),
    .CON(_01211_),
    .SN(_15702_));
 HAxp5_ASAP7_75t_SL _30788_ (.A(_01595_),
    .B(_01635_),
    .CON(_01213_),
    .SN(_15703_));
 HAxp5_ASAP7_75t_R _30789_ (.A(_01611_),
    .B(_01208_),
    .CON(_01215_),
    .SN(_15704_));
 HAxp5_ASAP7_75t_SL _30790_ (.A(_01611_),
    .B(_01208_),
    .CON(_01216_),
    .SN(_15705_));
 HAxp5_ASAP7_75t_SL _30791_ (.A(_01611_),
    .B(_01595_),
    .CON(_01217_),
    .SN(_15706_));
 HAxp5_ASAP7_75t_L _30792_ (.A(_01611_),
    .B(_01595_),
    .CON(_01218_),
    .SN(_15707_));
 HAxp5_ASAP7_75t_R _30793_ (.A(_01638_),
    .B(_01208_),
    .CON(_01220_),
    .SN(_01221_));
 HAxp5_ASAP7_75t_R _30794_ (.A(_01638_),
    .B(_01595_),
    .CON(_01222_),
    .SN(_15708_));
 HAxp5_ASAP7_75t_SL _30795_ (.A(_01638_),
    .B(_01595_),
    .CON(_01223_),
    .SN(_15709_));
 HAxp5_ASAP7_75t_R _30796_ (.A(_01633_),
    .B(_01208_),
    .CON(_01225_),
    .SN(_15710_));
 HAxp5_ASAP7_75t_R _30797_ (.A(_01633_),
    .B(_01208_),
    .CON(_01226_),
    .SN(_15711_));
 HAxp5_ASAP7_75t_R _30798_ (.A(_01633_),
    .B(_01595_),
    .CON(_01227_),
    .SN(_15712_));
 HAxp5_ASAP7_75t_SL _30799_ (.A(_02357_),
    .B(_02426_),
    .CON(_01230_),
    .SN(_01231_));
 HAxp5_ASAP7_75t_L _30800_ (.A(_02426_),
    .B(_02357_),
    .CON(_01232_),
    .SN(_15713_));
 HAxp5_ASAP7_75t_SL _30801_ (.A(_01233_),
    .B(_02426_),
    .CON(_01234_),
    .SN(_15714_));
 HAxp5_ASAP7_75t_SL _30802_ (.A(_02426_),
    .B(_01233_),
    .CON(_01235_),
    .SN(_15715_));
 HAxp5_ASAP7_75t_R _30803_ (.A(_01236_),
    .B(_02357_),
    .CON(_01237_),
    .SN(_15716_));
 HAxp5_ASAP7_75t_SL _30804_ (.A(_01236_),
    .B(_02357_),
    .CON(_01238_),
    .SN(_15717_));
 HAxp5_ASAP7_75t_SL _30805_ (.A(_01233_),
    .B(_01236_),
    .CON(_01239_),
    .SN(_15718_));
 HAxp5_ASAP7_75t_R _30806_ (.A(_01236_),
    .B(_01233_),
    .CON(_01240_),
    .SN(_15719_));
 HAxp5_ASAP7_75t_R _30807_ (.A(_02360_),
    .B(_02357_),
    .CON(_01242_),
    .SN(_01243_));
 HAxp5_ASAP7_75t_R _30808_ (.A(_02360_),
    .B(_01233_),
    .CON(_01244_),
    .SN(_15720_));
 HAxp5_ASAP7_75t_R _30809_ (.A(_02360_),
    .B(_01233_),
    .CON(_01245_),
    .SN(_15721_));
 HAxp5_ASAP7_75t_R _30810_ (.A(_02354_),
    .B(_02357_),
    .CON(_01247_),
    .SN(_15722_));
 HAxp5_ASAP7_75t_R _30811_ (.A(_02354_),
    .B(_02357_),
    .CON(_01248_),
    .SN(_15723_));
 HAxp5_ASAP7_75t_R _30812_ (.A(_02354_),
    .B(_01233_),
    .CON(_01249_),
    .SN(_15724_));
 HAxp5_ASAP7_75t_R _30813_ (.A(_02354_),
    .B(_01233_),
    .CON(_01250_),
    .SN(_15725_));
 HAxp5_ASAP7_75t_SL _30814_ (.A(_03043_),
    .B(_03052_),
    .CON(_01253_),
    .SN(_01254_));
 HAxp5_ASAP7_75t_R _30815_ (.A(_03052_),
    .B(_03043_),
    .CON(_01255_),
    .SN(_15726_));
 HAxp5_ASAP7_75t_R _30816_ (.A(_03052_),
    .B(_01256_),
    .CON(_01257_),
    .SN(_15727_));
 HAxp5_ASAP7_75t_L _30817_ (.A(_03052_),
    .B(_01256_),
    .CON(_01258_),
    .SN(_15728_));
 HAxp5_ASAP7_75t_R _30818_ (.A(_01259_),
    .B(_03043_),
    .CON(_01260_),
    .SN(_15729_));
 HAxp5_ASAP7_75t_L _30819_ (.A(_01259_),
    .B(_03043_),
    .CON(_01261_),
    .SN(_15730_));
 HAxp5_ASAP7_75t_L _30820_ (.A(_01256_),
    .B(_01259_),
    .CON(_01262_),
    .SN(_15731_));
 HAxp5_ASAP7_75t_SL _30821_ (.A(_01256_),
    .B(_01259_),
    .CON(_01263_),
    .SN(_15732_));
 HAxp5_ASAP7_75t_R _30822_ (.A(_03048_),
    .B(_03043_),
    .CON(_01265_),
    .SN(_01266_));
 HAxp5_ASAP7_75t_R _30823_ (.A(_03048_),
    .B(_01256_),
    .CON(_01267_),
    .SN(_15733_));
 HAxp5_ASAP7_75t_R _30824_ (.A(_03048_),
    .B(_01256_),
    .CON(_01268_),
    .SN(_15734_));
 HAxp5_ASAP7_75t_R _30825_ (.A(_03040_),
    .B(_03043_),
    .CON(_01270_),
    .SN(_15735_));
 HAxp5_ASAP7_75t_R _30826_ (.A(_03040_),
    .B(_03043_),
    .CON(_01271_),
    .SN(_15736_));
 HAxp5_ASAP7_75t_R _30827_ (.A(_03040_),
    .B(_01256_),
    .CON(_01272_),
    .SN(_15737_));
 HAxp5_ASAP7_75t_R _30828_ (.A(_03040_),
    .B(_01256_),
    .CON(_01273_),
    .SN(_15738_));
 HAxp5_ASAP7_75t_SL _30829_ (.A(_01275_),
    .B(_01274_),
    .CON(_01276_),
    .SN(_01277_));
 HAxp5_ASAP7_75t_L _30830_ (.A(_01274_),
    .B(_01275_),
    .CON(_01278_),
    .SN(_15739_));
 HAxp5_ASAP7_75t_L _30831_ (.A(_01274_),
    .B(_01279_),
    .CON(_01280_),
    .SN(_15740_));
 HAxp5_ASAP7_75t_L _30832_ (.A(_01274_),
    .B(_01279_),
    .CON(_01281_),
    .SN(_15741_));
 HAxp5_ASAP7_75t_R _30833_ (.A(_01282_),
    .B(_01275_),
    .CON(_01283_),
    .SN(_15742_));
 HAxp5_ASAP7_75t_R _30834_ (.A(_01282_),
    .B(_01275_),
    .CON(_01284_),
    .SN(_15743_));
 HAxp5_ASAP7_75t_L _30835_ (.A(_01282_),
    .B(_01279_),
    .CON(_01285_),
    .SN(_15744_));
 HAxp5_ASAP7_75t_SL _30836_ (.A(_01282_),
    .B(_01279_),
    .CON(_01286_),
    .SN(_15745_));
 HAxp5_ASAP7_75t_SL _30837_ (.A(_03731_),
    .B(_01275_),
    .CON(_01288_),
    .SN(_01289_));
 HAxp5_ASAP7_75t_SL _30838_ (.A(_03731_),
    .B(_01279_),
    .CON(_01290_),
    .SN(_15746_));
 HAxp5_ASAP7_75t_SL _30839_ (.A(_03731_),
    .B(_01279_),
    .CON(_01291_),
    .SN(_15747_));
 HAxp5_ASAP7_75t_SL _30840_ (.A(_03721_),
    .B(_01275_),
    .CON(_01293_),
    .SN(_15748_));
 HAxp5_ASAP7_75t_R _30841_ (.A(_03721_),
    .B(_01275_),
    .CON(_01294_),
    .SN(_15749_));
 HAxp5_ASAP7_75t_SL _30842_ (.A(_03721_),
    .B(_01279_),
    .CON(_01295_),
    .SN(_15750_));
 HAxp5_ASAP7_75t_SL _30843_ (.A(_03721_),
    .B(_01279_),
    .CON(_01296_),
    .SN(_15751_));
 HAxp5_ASAP7_75t_SL _30844_ (.A(_01298_),
    .B(_04448_),
    .CON(_01299_),
    .SN(_01300_));
 HAxp5_ASAP7_75t_SL _30845_ (.A(_04448_),
    .B(_01298_),
    .CON(_01301_),
    .SN(_15752_));
 HAxp5_ASAP7_75t_L _30846_ (.A(_04448_),
    .B(_01302_),
    .CON(_01303_),
    .SN(_15753_));
 HAxp5_ASAP7_75t_SL _30847_ (.A(_01302_),
    .B(_04448_),
    .CON(_01304_),
    .SN(_15754_));
 HAxp5_ASAP7_75t_R _30848_ (.A(_01305_),
    .B(_01298_),
    .CON(_01306_),
    .SN(_15755_));
 HAxp5_ASAP7_75t_SL _30849_ (.A(_01305_),
    .B(_01298_),
    .CON(_01307_),
    .SN(_15756_));
 HAxp5_ASAP7_75t_L _30850_ (.A(_01305_),
    .B(_01302_),
    .CON(_01308_),
    .SN(_15757_));
 HAxp5_ASAP7_75t_R _30851_ (.A(_01305_),
    .B(_01302_),
    .CON(_01309_),
    .SN(_15758_));
 HAxp5_ASAP7_75t_SL _30852_ (.A(_04408_),
    .B(_01298_),
    .CON(_01311_),
    .SN(_01312_));
 HAxp5_ASAP7_75t_R _30853_ (.A(_04408_),
    .B(_01302_),
    .CON(_01313_),
    .SN(_15759_));
 HAxp5_ASAP7_75t_SL _30854_ (.A(_04408_),
    .B(_01302_),
    .CON(_01314_),
    .SN(_15760_));
 HAxp5_ASAP7_75t_R _30855_ (.A(_04402_),
    .B(_01298_),
    .CON(_01316_),
    .SN(_15761_));
 HAxp5_ASAP7_75t_SL _30856_ (.A(_04402_),
    .B(_01298_),
    .CON(_01317_),
    .SN(_15762_));
 HAxp5_ASAP7_75t_R _30857_ (.A(_04402_),
    .B(_01302_),
    .CON(_01318_),
    .SN(_15763_));
 HAxp5_ASAP7_75t_SL _30858_ (.A(_04402_),
    .B(_01302_),
    .CON(_01319_),
    .SN(_15764_));
 HAxp5_ASAP7_75t_SL _30859_ (.A(_01321_),
    .B(_05071_),
    .CON(_01322_),
    .SN(_01323_));
 HAxp5_ASAP7_75t_L _30860_ (.A(_05071_),
    .B(_01321_),
    .CON(_01324_),
    .SN(_15765_));
 HAxp5_ASAP7_75t_R _30861_ (.A(_05071_),
    .B(_05040_),
    .CON(_01326_),
    .SN(_15766_));
 HAxp5_ASAP7_75t_R _30862_ (.A(_05051_),
    .B(_01321_),
    .CON(_01328_),
    .SN(_15767_));
 HAxp5_ASAP7_75t_SL _30863_ (.A(_05051_),
    .B(_01321_),
    .CON(_01329_),
    .SN(_15768_));
 HAxp5_ASAP7_75t_R _30864_ (.A(_05051_),
    .B(_05040_),
    .CON(_01330_),
    .SN(_15769_));
 HAxp5_ASAP7_75t_SL _30865_ (.A(_05040_),
    .B(_05051_),
    .CON(_01331_),
    .SN(_15770_));
 HAxp5_ASAP7_75t_R _30866_ (.A(_05074_),
    .B(_01321_),
    .CON(_01333_),
    .SN(_01334_));
 HAxp5_ASAP7_75t_R _30867_ (.A(_05074_),
    .B(_05040_),
    .CON(_01335_),
    .SN(_15771_));
 HAxp5_ASAP7_75t_R _30868_ (.A(_05074_),
    .B(_05040_),
    .CON(_01336_),
    .SN(_15772_));
 HAxp5_ASAP7_75t_R _30869_ (.A(_05068_),
    .B(_01321_),
    .CON(_01338_),
    .SN(_15773_));
 HAxp5_ASAP7_75t_R _30870_ (.A(_05068_),
    .B(_01321_),
    .CON(_01339_),
    .SN(_15774_));
 HAxp5_ASAP7_75t_R _30871_ (.A(_05068_),
    .B(_05040_),
    .CON(_01340_),
    .SN(_15775_));
 HAxp5_ASAP7_75t_SL _30872_ (.A(_01342_),
    .B(_05761_),
    .CON(_01343_),
    .SN(_01344_));
 HAxp5_ASAP7_75t_L _30873_ (.A(_05761_),
    .B(_01342_),
    .CON(_01345_),
    .SN(_15776_));
 HAxp5_ASAP7_75t_R _30874_ (.A(_05761_),
    .B(_05722_),
    .CON(_01347_),
    .SN(_15777_));
 HAxp5_ASAP7_75t_R _30875_ (.A(_05737_),
    .B(_01342_),
    .CON(_01349_),
    .SN(_15778_));
 HAxp5_ASAP7_75t_SL _30876_ (.A(_01342_),
    .B(_05737_),
    .CON(_01350_),
    .SN(_15779_));
 HAxp5_ASAP7_75t_R _30877_ (.A(_05737_),
    .B(_05722_),
    .CON(_01351_),
    .SN(_15780_));
 HAxp5_ASAP7_75t_L _30878_ (.A(_05737_),
    .B(_05722_),
    .CON(_01352_),
    .SN(_15781_));
 HAxp5_ASAP7_75t_R _30879_ (.A(_05764_),
    .B(_01342_),
    .CON(_01354_),
    .SN(_01355_));
 HAxp5_ASAP7_75t_SL _30880_ (.A(_05764_),
    .B(_05722_),
    .CON(_01356_),
    .SN(_15782_));
 HAxp5_ASAP7_75t_SL _30881_ (.A(_05764_),
    .B(_05722_),
    .CON(_01357_),
    .SN(_15783_));
 HAxp5_ASAP7_75t_SL _30882_ (.A(_05757_),
    .B(_01342_),
    .CON(_01359_),
    .SN(_15784_));
 HAxp5_ASAP7_75t_R _30883_ (.A(_05757_),
    .B(_01342_),
    .CON(_01360_),
    .SN(_15785_));
 HAxp5_ASAP7_75t_R _30884_ (.A(_05757_),
    .B(_05722_),
    .CON(_01361_),
    .SN(_15786_));
 HAxp5_ASAP7_75t_SL _30885_ (.A(_06439_),
    .B(_06424_),
    .CON(_01364_),
    .SN(_01365_));
 HAxp5_ASAP7_75t_R _30886_ (.A(_06424_),
    .B(_06439_),
    .CON(_01366_),
    .SN(_15787_));
 HAxp5_ASAP7_75t_L _30887_ (.A(_06424_),
    .B(_06392_),
    .CON(_01368_),
    .SN(_15788_));
 HAxp5_ASAP7_75t_SL _30888_ (.A(_06439_),
    .B(_06405_),
    .CON(_01370_),
    .SN(_15789_));
 HAxp5_ASAP7_75t_R _30889_ (.A(_06405_),
    .B(_06439_),
    .CON(_01371_),
    .SN(_15790_));
 HAxp5_ASAP7_75t_R _30890_ (.A(_06405_),
    .B(_06392_),
    .CON(_01372_),
    .SN(_15791_));
 HAxp5_ASAP7_75t_R _30891_ (.A(_06405_),
    .B(_06392_),
    .CON(_01373_),
    .SN(_15792_));
 HAxp5_ASAP7_75t_R _30892_ (.A(_06428_),
    .B(_06439_),
    .CON(_01375_),
    .SN(_01376_));
 HAxp5_ASAP7_75t_R _30893_ (.A(_06428_),
    .B(_06392_),
    .CON(_01377_),
    .SN(_15793_));
 HAxp5_ASAP7_75t_SL _30894_ (.A(_06428_),
    .B(_06392_),
    .CON(_01378_),
    .SN(_15794_));
 HAxp5_ASAP7_75t_R _30895_ (.A(_06421_),
    .B(_06439_),
    .CON(_01380_),
    .SN(_15795_));
 HAxp5_ASAP7_75t_R _30896_ (.A(_06421_),
    .B(_06439_),
    .CON(_01381_),
    .SN(_15796_));
 HAxp5_ASAP7_75t_R _30897_ (.A(_06421_),
    .B(_06392_),
    .CON(_01382_),
    .SN(_15797_));
 HAxp5_ASAP7_75t_SL _30898_ (.A(_01384_),
    .B(_07116_),
    .CON(_01385_),
    .SN(_01386_));
 HAxp5_ASAP7_75t_SL _30899_ (.A(_07116_),
    .B(_01384_),
    .CON(_01387_),
    .SN(_15798_));
 HAxp5_ASAP7_75t_SL _30900_ (.A(_07116_),
    .B(_07081_),
    .CON(_01389_),
    .SN(_15799_));
 HAxp5_ASAP7_75t_R _30901_ (.A(_07094_),
    .B(_01384_),
    .CON(_01391_),
    .SN(_15800_));
 HAxp5_ASAP7_75t_SL _30902_ (.A(_07094_),
    .B(_01384_),
    .CON(_01392_),
    .SN(_15801_));
 HAxp5_ASAP7_75t_SL _30903_ (.A(_07094_),
    .B(_07081_),
    .CON(_01393_),
    .SN(_15802_));
 HAxp5_ASAP7_75t_R _30904_ (.A(_07094_),
    .B(_07081_),
    .CON(_01394_),
    .SN(_15803_));
 HAxp5_ASAP7_75t_SL _30905_ (.A(_07119_),
    .B(_01384_),
    .CON(_01396_),
    .SN(_01397_));
 HAxp5_ASAP7_75t_SL _30906_ (.A(_07119_),
    .B(_07081_),
    .CON(_01398_),
    .SN(_15804_));
 HAxp5_ASAP7_75t_SL _30907_ (.A(_07119_),
    .B(_07081_),
    .CON(_01399_),
    .SN(_15805_));
 HAxp5_ASAP7_75t_SL _30908_ (.A(_07112_),
    .B(_01384_),
    .CON(_01401_),
    .SN(_15806_));
 HAxp5_ASAP7_75t_SL _30909_ (.A(_07112_),
    .B(_01384_),
    .CON(_01402_),
    .SN(_15807_));
 HAxp5_ASAP7_75t_R _30910_ (.A(_07112_),
    .B(_07081_),
    .CON(_01403_),
    .SN(_15808_));
 DFFHQNx1_ASAP7_75t_SL \dcnt[0]$_SDFFE_PN0P_  (.CLK(clk),
    .D(_01404_),
    .QN(_00572_));
 DFFHQNx1_ASAP7_75t_SL \dcnt[1]$_SDFFE_PN0P_  (.CLK(clk),
    .D(_01405_),
    .QN(_00571_));
 DFFHQNx1_ASAP7_75t_SL \dcnt[2]$_SDFFE_PP0P_  (.CLK(clk),
    .D(_01406_),
    .QN(_00570_));
 DFFHQNx1_ASAP7_75t_SL \dcnt[3]$_SDFFE_PN0P_  (.CLK(clk),
    .D(_01407_),
    .QN(_00411_));
 DFFHQNx1_ASAP7_75t_SL \done$_DFF_P_  (.CLK(clk),
    .D(_00160_),
    .QN(_00573_));
 DFFHQNx2_ASAP7_75t_SL \ld_r$_DFF_P_  (.CLK(clk),
    .D(ld),
    .QN(_00574_));
 DFFHQNx1_ASAP7_75t_SL \sa00_sr[0]$_DFF_P_  (.CLK(clk),
    .D(_00032_),
    .QN(_00575_));
 DFFHQNx1_ASAP7_75t_SL \sa00_sr[1]$_DFF_P_  (.CLK(clk),
    .D(_00033_),
    .QN(_00576_));
 DFFHQNx1_ASAP7_75t_SL \sa00_sr[2]$_DFF_P_  (.CLK(clk),
    .D(_00034_),
    .QN(_00577_));
 DFFHQNx1_ASAP7_75t_SL \sa00_sr[3]$_DFF_P_  (.CLK(clk),
    .D(_00035_),
    .QN(_00578_));
 DFFHQNx1_ASAP7_75t_SL \sa00_sr[4]$_DFF_P_  (.CLK(clk),
    .D(_00036_),
    .QN(_00579_));
 DFFHQNx1_ASAP7_75t_SL \sa00_sr[5]$_DFF_P_  (.CLK(clk),
    .D(_00037_),
    .QN(_00580_));
 DFFHQNx1_ASAP7_75t_SL \sa00_sr[6]$_DFF_P_  (.CLK(clk),
    .D(_00038_),
    .QN(_00581_));
 DFFHQNx1_ASAP7_75t_SL \sa00_sr[7]$_DFF_P_  (.CLK(clk),
    .D(_00039_),
    .QN(_00582_));
 DFFHQNx1_ASAP7_75t_SL \sa01_sr[0]$_DFF_P_  (.CLK(clk),
    .D(_00040_),
    .QN(_00583_));
 DFFHQNx1_ASAP7_75t_SL \sa01_sr[1]$_DFF_P_  (.CLK(clk),
    .D(_00041_),
    .QN(_00584_));
 DFFHQNx1_ASAP7_75t_SL \sa01_sr[2]$_DFF_P_  (.CLK(clk),
    .D(_00042_),
    .QN(_00585_));
 DFFHQNx1_ASAP7_75t_SL \sa01_sr[3]$_DFF_P_  (.CLK(clk),
    .D(_00043_),
    .QN(_00586_));
 DFFHQNx1_ASAP7_75t_SL \sa01_sr[4]$_DFF_P_  (.CLK(clk),
    .D(_00044_),
    .QN(_00587_));
 DFFHQNx1_ASAP7_75t_SL \sa01_sr[5]$_DFF_P_  (.CLK(clk),
    .D(_00045_),
    .QN(_00588_));
 DFFHQNx1_ASAP7_75t_SL \sa01_sr[6]$_DFF_P_  (.CLK(clk),
    .D(_00046_),
    .QN(_00589_));
 DFFHQNx1_ASAP7_75t_SL \sa01_sr[7]$_DFF_P_  (.CLK(clk),
    .D(_00047_),
    .QN(_00590_));
 DFFHQNx1_ASAP7_75t_SL \sa02_sr[0]$_DFF_P_  (.CLK(clk),
    .D(_00048_),
    .QN(_00591_));
 DFFHQNx1_ASAP7_75t_SL \sa02_sr[1]$_DFF_P_  (.CLK(clk),
    .D(_00049_),
    .QN(_00592_));
 DFFHQNx1_ASAP7_75t_SL \sa02_sr[2]$_DFF_P_  (.CLK(clk),
    .D(_00050_),
    .QN(_00593_));
 DFFHQNx1_ASAP7_75t_SL \sa02_sr[3]$_DFF_P_  (.CLK(clk),
    .D(_00051_),
    .QN(_00594_));
 DFFHQNx1_ASAP7_75t_SL \sa02_sr[4]$_DFF_P_  (.CLK(clk),
    .D(_00052_),
    .QN(_00595_));
 DFFHQNx1_ASAP7_75t_SL \sa02_sr[5]$_DFF_P_  (.CLK(clk),
    .D(_00053_),
    .QN(_00596_));
 DFFHQNx1_ASAP7_75t_SL \sa02_sr[6]$_DFF_P_  (.CLK(clk),
    .D(_00054_),
    .QN(_00597_));
 DFFHQNx1_ASAP7_75t_SL \sa02_sr[7]$_DFF_P_  (.CLK(clk),
    .D(_00055_),
    .QN(_00598_));
 DFFHQNx1_ASAP7_75t_SL \sa03_sr[0]$_DFF_P_  (.CLK(clk),
    .D(_00056_),
    .QN(_00599_));
 DFFHQNx1_ASAP7_75t_SL \sa03_sr[1]$_DFF_P_  (.CLK(clk),
    .D(_00057_),
    .QN(_00600_));
 DFFHQNx1_ASAP7_75t_SL \sa03_sr[2]$_DFF_P_  (.CLK(clk),
    .D(_00058_),
    .QN(_00601_));
 DFFHQNx1_ASAP7_75t_SL \sa03_sr[3]$_DFF_P_  (.CLK(clk),
    .D(_00059_),
    .QN(_00602_));
 DFFHQNx1_ASAP7_75t_SL \sa03_sr[4]$_DFF_P_  (.CLK(clk),
    .D(_00060_),
    .QN(_00603_));
 DFFHQNx1_ASAP7_75t_SL \sa03_sr[5]$_DFF_P_  (.CLK(clk),
    .D(_00061_),
    .QN(_00604_));
 DFFHQNx1_ASAP7_75t_SL \sa03_sr[6]$_DFF_P_  (.CLK(clk),
    .D(_00062_),
    .QN(_00605_));
 DFFHQNx1_ASAP7_75t_SL \sa03_sr[7]$_DFF_P_  (.CLK(clk),
    .D(_00063_),
    .QN(_00606_));
 DFFHQNx2_ASAP7_75t_SL \sa10_sr[0]$_DFF_P_  (.CLK(clk),
    .D(_00072_),
    .QN(_00607_));
 DFFHQNx1_ASAP7_75t_SL \sa10_sr[1]$_DFF_P_  (.CLK(clk),
    .D(_00073_),
    .QN(_00608_));
 DFFHQNx1_ASAP7_75t_SL \sa10_sr[2]$_DFF_P_  (.CLK(clk),
    .D(_00074_),
    .QN(_00609_));
 DFFHQNx1_ASAP7_75t_SL \sa10_sr[3]$_DFF_P_  (.CLK(clk),
    .D(_00075_),
    .QN(_00610_));
 DFFHQNx1_ASAP7_75t_SL \sa10_sr[4]$_DFF_P_  (.CLK(clk),
    .D(_00076_),
    .QN(_00611_));
 DFFHQNx1_ASAP7_75t_SL \sa10_sr[5]$_DFF_P_  (.CLK(clk),
    .D(_00077_),
    .QN(_00612_));
 DFFHQNx1_ASAP7_75t_SL \sa10_sr[6]$_DFF_P_  (.CLK(clk),
    .D(_00078_),
    .QN(_00613_));
 DFFHQNx1_ASAP7_75t_SL \sa10_sr[7]$_DFF_P_  (.CLK(clk),
    .D(_00079_),
    .QN(_00614_));
 DFFHQNx2_ASAP7_75t_SL \sa11_sr[0]$_DFF_P_  (.CLK(clk),
    .D(_00080_),
    .QN(_00615_));
 DFFHQNx1_ASAP7_75t_SL \sa11_sr[1]$_DFF_P_  (.CLK(clk),
    .D(_00081_),
    .QN(_00616_));
 DFFHQNx1_ASAP7_75t_SL \sa11_sr[2]$_DFF_P_  (.CLK(clk),
    .D(_00082_),
    .QN(_00617_));
 DFFHQNx1_ASAP7_75t_SL \sa11_sr[3]$_DFF_P_  (.CLK(clk),
    .D(_00083_),
    .QN(_00618_));
 DFFHQNx1_ASAP7_75t_SL \sa11_sr[4]$_DFF_P_  (.CLK(clk),
    .D(_00084_),
    .QN(_00619_));
 DFFHQNx1_ASAP7_75t_SL \sa11_sr[5]$_DFF_P_  (.CLK(clk),
    .D(_00085_),
    .QN(_00620_));
 DFFHQNx1_ASAP7_75t_SL \sa11_sr[6]$_DFF_P_  (.CLK(clk),
    .D(_00086_),
    .QN(_00621_));
 DFFHQNx1_ASAP7_75t_SL \sa11_sr[7]$_DFF_P_  (.CLK(clk),
    .D(_00087_),
    .QN(_00622_));
 DFFHQNx2_ASAP7_75t_SL \sa12_sr[0]$_DFF_P_  (.CLK(clk),
    .D(_00088_),
    .QN(_00623_));
 DFFHQNx1_ASAP7_75t_SL \sa12_sr[1]$_DFF_P_  (.CLK(clk),
    .D(_00089_),
    .QN(_00624_));
 DFFHQNx1_ASAP7_75t_SL \sa12_sr[2]$_DFF_P_  (.CLK(clk),
    .D(_00090_),
    .QN(_00625_));
 DFFHQNx1_ASAP7_75t_SL \sa12_sr[3]$_DFF_P_  (.CLK(clk),
    .D(_00091_),
    .QN(_00626_));
 DFFHQNx1_ASAP7_75t_SL \sa12_sr[4]$_DFF_P_  (.CLK(clk),
    .D(_00092_),
    .QN(_00627_));
 DFFHQNx1_ASAP7_75t_SL \sa12_sr[5]$_DFF_P_  (.CLK(clk),
    .D(_00093_),
    .QN(_00628_));
 DFFHQNx1_ASAP7_75t_SL \sa12_sr[6]$_DFF_P_  (.CLK(clk),
    .D(_00094_),
    .QN(_00629_));
 DFFHQNx1_ASAP7_75t_SL \sa12_sr[7]$_DFF_P_  (.CLK(clk),
    .D(_00095_),
    .QN(_00630_));
 DFFHQNx2_ASAP7_75t_SL \sa13_sr[0]$_DFF_P_  (.CLK(clk),
    .D(_00064_),
    .QN(_00631_));
 DFFHQNx1_ASAP7_75t_SL \sa13_sr[1]$_DFF_P_  (.CLK(clk),
    .D(_00065_),
    .QN(_00632_));
 DFFHQNx1_ASAP7_75t_SL \sa13_sr[2]$_DFF_P_  (.CLK(clk),
    .D(_00066_),
    .QN(_00633_));
 DFFHQNx1_ASAP7_75t_SL \sa13_sr[3]$_DFF_P_  (.CLK(clk),
    .D(_00067_),
    .QN(_00634_));
 DFFHQNx1_ASAP7_75t_SL \sa13_sr[4]$_DFF_P_  (.CLK(clk),
    .D(_00068_),
    .QN(_00635_));
 DFFHQNx1_ASAP7_75t_SL \sa13_sr[5]$_DFF_P_  (.CLK(clk),
    .D(_00069_),
    .QN(_00636_));
 DFFHQNx1_ASAP7_75t_SL \sa13_sr[6]$_DFF_P_  (.CLK(clk),
    .D(_00070_),
    .QN(_00637_));
 DFFHQNx1_ASAP7_75t_SL \sa13_sr[7]$_DFF_P_  (.CLK(clk),
    .D(_00071_),
    .QN(_00638_));
 DFFHQNx1_ASAP7_75t_SL \sa20_sr[0]$_DFF_P_  (.CLK(clk),
    .D(_00112_),
    .QN(_00639_));
 DFFHQNx2_ASAP7_75t_SL \sa20_sr[1]$_DFF_P_  (.CLK(clk),
    .D(_00113_),
    .QN(_00640_));
 DFFHQNx1_ASAP7_75t_SL \sa20_sr[2]$_DFF_P_  (.CLK(clk),
    .D(_00114_),
    .QN(_00641_));
 DFFHQNx1_ASAP7_75t_SL \sa20_sr[3]$_DFF_P_  (.CLK(clk),
    .D(_00115_),
    .QN(_00642_));
 DFFHQNx1_ASAP7_75t_SL \sa20_sr[4]$_DFF_P_  (.CLK(clk),
    .D(_00116_),
    .QN(_00643_));
 DFFHQNx1_ASAP7_75t_SL \sa20_sr[5]$_DFF_P_  (.CLK(clk),
    .D(_00117_),
    .QN(_00644_));
 DFFHQNx1_ASAP7_75t_SL \sa20_sr[6]$_DFF_P_  (.CLK(clk),
    .D(_00118_),
    .QN(_00645_));
 DFFHQNx1_ASAP7_75t_SL \sa20_sr[7]$_DFF_P_  (.CLK(clk),
    .D(_00119_),
    .QN(_00646_));
 DFFHQNx1_ASAP7_75t_SL \sa21_sr[0]$_DFF_P_  (.CLK(clk),
    .D(_00120_),
    .QN(_00647_));
 DFFHQNx1_ASAP7_75t_SL \sa21_sr[1]$_DFF_P_  (.CLK(clk),
    .D(_00121_),
    .QN(_00648_));
 DFFHQNx1_ASAP7_75t_SL \sa21_sr[2]$_DFF_P_  (.CLK(clk),
    .D(_00122_),
    .QN(_00649_));
 DFFHQNx1_ASAP7_75t_SL \sa21_sr[3]$_DFF_P_  (.CLK(clk),
    .D(_00123_),
    .QN(_00650_));
 DFFHQNx1_ASAP7_75t_SL \sa21_sr[4]$_DFF_P_  (.CLK(clk),
    .D(_00124_),
    .QN(_00651_));
 DFFHQNx1_ASAP7_75t_SL \sa21_sr[5]$_DFF_P_  (.CLK(clk),
    .D(_00125_),
    .QN(_00652_));
 DFFHQNx1_ASAP7_75t_SL \sa21_sr[6]$_DFF_P_  (.CLK(clk),
    .D(_00126_),
    .QN(_00653_));
 DFFHQNx1_ASAP7_75t_SL \sa21_sr[7]$_DFF_P_  (.CLK(clk),
    .D(_00127_),
    .QN(_00654_));
 DFFHQNx1_ASAP7_75t_SL \sa22_sr[0]$_DFF_P_  (.CLK(clk),
    .D(_00096_),
    .QN(_00655_));
 DFFHQNx2_ASAP7_75t_SL \sa22_sr[1]$_DFF_P_  (.CLK(clk),
    .D(_00097_),
    .QN(_00656_));
 DFFHQNx1_ASAP7_75t_SL \sa22_sr[2]$_DFF_P_  (.CLK(clk),
    .D(_00098_),
    .QN(_00657_));
 DFFHQNx1_ASAP7_75t_SL \sa22_sr[3]$_DFF_P_  (.CLK(clk),
    .D(_00099_),
    .QN(_00658_));
 DFFHQNx1_ASAP7_75t_SL \sa22_sr[4]$_DFF_P_  (.CLK(clk),
    .D(_00100_),
    .QN(_00659_));
 DFFHQNx1_ASAP7_75t_SL \sa22_sr[5]$_DFF_P_  (.CLK(clk),
    .D(_00101_),
    .QN(_00660_));
 DFFHQNx1_ASAP7_75t_SL \sa22_sr[6]$_DFF_P_  (.CLK(clk),
    .D(_00102_),
    .QN(_00661_));
 DFFHQNx1_ASAP7_75t_SL \sa22_sr[7]$_DFF_P_  (.CLK(clk),
    .D(_00103_),
    .QN(_00662_));
 DFFHQNx1_ASAP7_75t_SL \sa23_sr[0]$_DFF_P_  (.CLK(clk),
    .D(_00104_),
    .QN(_00663_));
 DFFHQNx2_ASAP7_75t_SL \sa23_sr[1]$_DFF_P_  (.CLK(clk),
    .D(_00105_),
    .QN(_00664_));
 DFFHQNx1_ASAP7_75t_SL \sa23_sr[2]$_DFF_P_  (.CLK(clk),
    .D(_00106_),
    .QN(_00665_));
 DFFHQNx1_ASAP7_75t_SL \sa23_sr[3]$_DFF_P_  (.CLK(clk),
    .D(_00107_),
    .QN(_00666_));
 DFFHQNx1_ASAP7_75t_SL \sa23_sr[4]$_DFF_P_  (.CLK(clk),
    .D(_00108_),
    .QN(_00667_));
 DFFHQNx1_ASAP7_75t_SL \sa23_sr[5]$_DFF_P_  (.CLK(clk),
    .D(_00109_),
    .QN(_00668_));
 DFFHQNx1_ASAP7_75t_SL \sa23_sr[6]$_DFF_P_  (.CLK(clk),
    .D(_00110_),
    .QN(_00669_));
 DFFHQNx1_ASAP7_75t_SL \sa23_sr[7]$_DFF_P_  (.CLK(clk),
    .D(_00111_),
    .QN(_00670_));
 DFFHQNx1_ASAP7_75t_SL \sa30_sr[0]$_DFF_P_  (.CLK(clk),
    .D(_00152_),
    .QN(_00671_));
 DFFHQNx1_ASAP7_75t_SL \sa30_sr[1]$_DFF_P_  (.CLK(clk),
    .D(_00153_),
    .QN(_00672_));
 DFFHQNx1_ASAP7_75t_SL \sa30_sr[2]$_DFF_P_  (.CLK(clk),
    .D(_00154_),
    .QN(_00673_));
 DFFHQNx1_ASAP7_75t_SL \sa30_sr[3]$_DFF_P_  (.CLK(clk),
    .D(_00155_),
    .QN(_00674_));
 DFFHQNx1_ASAP7_75t_SL \sa30_sr[4]$_DFF_P_  (.CLK(clk),
    .D(_00156_),
    .QN(_00675_));
 DFFHQNx1_ASAP7_75t_SL \sa30_sr[5]$_DFF_P_  (.CLK(clk),
    .D(_00157_),
    .QN(_00676_));
 DFFHQNx1_ASAP7_75t_SL \sa30_sr[6]$_DFF_P_  (.CLK(clk),
    .D(_00158_),
    .QN(_00677_));
 DFFHQNx2_ASAP7_75t_SL \sa30_sr[7]$_DFF_P_  (.CLK(clk),
    .D(_00159_),
    .QN(_00678_));
 DFFHQNx1_ASAP7_75t_SL \sa31_sr[0]$_DFF_P_  (.CLK(clk),
    .D(_00128_),
    .QN(_00679_));
 DFFHQNx1_ASAP7_75t_SL \sa31_sr[1]$_DFF_P_  (.CLK(clk),
    .D(_00129_),
    .QN(_00680_));
 DFFHQNx1_ASAP7_75t_SL \sa31_sr[2]$_DFF_P_  (.CLK(clk),
    .D(_00130_),
    .QN(_00681_));
 DFFHQNx1_ASAP7_75t_SL \sa31_sr[3]$_DFF_P_  (.CLK(clk),
    .D(_00131_),
    .QN(_00682_));
 DFFHQNx1_ASAP7_75t_SL \sa31_sr[4]$_DFF_P_  (.CLK(clk),
    .D(_00132_),
    .QN(_00683_));
 DFFHQNx1_ASAP7_75t_SL \sa31_sr[5]$_DFF_P_  (.CLK(clk),
    .D(_00133_),
    .QN(_00684_));
 DFFHQNx1_ASAP7_75t_SL \sa31_sr[6]$_DFF_P_  (.CLK(clk),
    .D(_00134_),
    .QN(_00685_));
 DFFHQNx1_ASAP7_75t_SL \sa31_sr[7]$_DFF_P_  (.CLK(clk),
    .D(_00135_),
    .QN(_00686_));
 DFFHQNx1_ASAP7_75t_SL \sa32_sr[0]$_DFF_P_  (.CLK(clk),
    .D(_00136_),
    .QN(_00687_));
 DFFHQNx1_ASAP7_75t_SL \sa32_sr[1]$_DFF_P_  (.CLK(clk),
    .D(_00137_),
    .QN(_00688_));
 DFFHQNx1_ASAP7_75t_SL \sa32_sr[2]$_DFF_P_  (.CLK(clk),
    .D(_00138_),
    .QN(_00689_));
 DFFHQNx1_ASAP7_75t_SL \sa32_sr[3]$_DFF_P_  (.CLK(clk),
    .D(_00139_),
    .QN(_00690_));
 DFFHQNx1_ASAP7_75t_SL \sa32_sr[4]$_DFF_P_  (.CLK(clk),
    .D(_00140_),
    .QN(_00691_));
 DFFHQNx1_ASAP7_75t_SL \sa32_sr[5]$_DFF_P_  (.CLK(clk),
    .D(_00141_),
    .QN(_00692_));
 DFFHQNx1_ASAP7_75t_SL \sa32_sr[6]$_DFF_P_  (.CLK(clk),
    .D(_00142_),
    .QN(_00693_));
 DFFHQNx2_ASAP7_75t_SL \sa32_sr[7]$_DFF_P_  (.CLK(clk),
    .D(_00143_),
    .QN(_00694_));
 DFFHQNx1_ASAP7_75t_SL \sa33_sr[0]$_DFF_P_  (.CLK(clk),
    .D(_00144_),
    .QN(_00695_));
 DFFHQNx1_ASAP7_75t_SL \sa33_sr[1]$_DFF_P_  (.CLK(clk),
    .D(_00145_),
    .QN(_00696_));
 DFFHQNx1_ASAP7_75t_SL \sa33_sr[2]$_DFF_P_  (.CLK(clk),
    .D(_00146_),
    .QN(_00697_));
 DFFHQNx1_ASAP7_75t_SL \sa33_sr[3]$_DFF_P_  (.CLK(clk),
    .D(_00147_),
    .QN(_00698_));
 DFFHQNx1_ASAP7_75t_SL \sa33_sr[4]$_DFF_P_  (.CLK(clk),
    .D(_00148_),
    .QN(_00699_));
 DFFHQNx1_ASAP7_75t_SL \sa33_sr[5]$_DFF_P_  (.CLK(clk),
    .D(_00149_),
    .QN(_00700_));
 DFFHQNx1_ASAP7_75t_SL \sa33_sr[6]$_DFF_P_  (.CLK(clk),
    .D(_00150_),
    .QN(_00701_));
 DFFHQNx1_ASAP7_75t_SL \sa33_sr[7]$_DFF_P_  (.CLK(clk),
    .D(_00151_),
    .QN(_00569_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[0]$_DFFE_PP_  (.CLK(clk),
    .D(_01408_),
    .QN(_00409_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[100]$_DFFE_PP_  (.CLK(clk),
    .D(_01409_),
    .QN(_00568_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[101]$_DFFE_PP_  (.CLK(clk),
    .D(_01410_),
    .QN(_00567_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[102]$_DFFE_PP_  (.CLK(clk),
    .D(_01411_),
    .QN(_00566_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[103]$_DFFE_PP_  (.CLK(clk),
    .D(_01412_),
    .QN(_00565_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[104]$_DFFE_PP_  (.CLK(clk),
    .D(_01413_),
    .QN(_00469_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[105]$_DFFE_PP_  (.CLK(clk),
    .D(_01414_),
    .QN(_00468_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[106]$_DFFE_PP_  (.CLK(clk),
    .D(_01415_),
    .QN(_00470_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[107]$_DFFE_PP_  (.CLK(clk),
    .D(_01416_),
    .QN(_00564_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[108]$_DFFE_PP_  (.CLK(clk),
    .D(_01417_),
    .QN(_00563_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[109]$_DFFE_PP_  (.CLK(clk),
    .D(_01418_),
    .QN(_00562_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[10]$_DFFE_PP_  (.CLK(clk),
    .D(_01419_),
    .QN(_00479_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[110]$_DFFE_PP_  (.CLK(clk),
    .D(_01420_),
    .QN(_00561_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[111]$_DFFE_PP_  (.CLK(clk),
    .D(_01421_),
    .QN(_00560_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[112]$_DFFE_PP_  (.CLK(clk),
    .D(_01422_),
    .QN(_00457_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[113]$_DFFE_PP_  (.CLK(clk),
    .D(_01423_),
    .QN(_00456_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[114]$_DFFE_PP_  (.CLK(clk),
    .D(_01424_),
    .QN(_00458_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[115]$_DFFE_PP_  (.CLK(clk),
    .D(_01425_),
    .QN(_00559_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[116]$_DFFE_PP_  (.CLK(clk),
    .D(_01426_),
    .QN(_00558_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[117]$_DFFE_PP_  (.CLK(clk),
    .D(_01427_),
    .QN(_00557_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[118]$_DFFE_PP_  (.CLK(clk),
    .D(_01428_),
    .QN(_00556_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[119]$_DFFE_PP_  (.CLK(clk),
    .D(_01429_),
    .QN(_00555_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[11]$_DFFE_PP_  (.CLK(clk),
    .D(_01430_),
    .QN(_00554_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[120]$_DFFE_PP_  (.CLK(clk),
    .D(_01431_),
    .QN(_00445_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[121]$_DFFE_PP_  (.CLK(clk),
    .D(_01432_),
    .QN(_00444_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[122]$_DFFE_PP_  (.CLK(clk),
    .D(_01433_),
    .QN(_00446_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[123]$_DFFE_PP_  (.CLK(clk),
    .D(_01434_),
    .QN(_00553_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[124]$_DFFE_PP_  (.CLK(clk),
    .D(_01435_),
    .QN(_00552_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[125]$_DFFE_PP_  (.CLK(clk),
    .D(_01436_),
    .QN(_00551_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[126]$_DFFE_PP_  (.CLK(clk),
    .D(_01437_),
    .QN(_00550_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[127]$_DFFE_PP_  (.CLK(clk),
    .D(_01438_),
    .QN(_00549_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[12]$_DFFE_PP_  (.CLK(clk),
    .D(_01439_),
    .QN(_00548_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[13]$_DFFE_PP_  (.CLK(clk),
    .D(_01440_),
    .QN(_00547_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[14]$_DFFE_PP_  (.CLK(clk),
    .D(_01441_),
    .QN(_00546_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[15]$_DFFE_PP_  (.CLK(clk),
    .D(_01442_),
    .QN(_00545_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[16]$_DFFE_PP_  (.CLK(clk),
    .D(_01443_),
    .QN(_00466_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[17]$_DFFE_PP_  (.CLK(clk),
    .D(_01444_),
    .QN(_00465_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[18]$_DFFE_PP_  (.CLK(clk),
    .D(_01445_),
    .QN(_00467_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[19]$_DFFE_PP_  (.CLK(clk),
    .D(_01446_),
    .QN(_00544_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[1]$_DFFE_PP_  (.CLK(clk),
    .D(_01447_),
    .QN(_00408_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[20]$_DFFE_PP_  (.CLK(clk),
    .D(_01448_),
    .QN(_00543_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[21]$_DFFE_PP_  (.CLK(clk),
    .D(_01449_),
    .QN(_00542_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[22]$_DFFE_PP_  (.CLK(clk),
    .D(_01450_),
    .QN(_00541_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[23]$_DFFE_PP_  (.CLK(clk),
    .D(_01451_),
    .QN(_00540_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[24]$_DFFE_PP_  (.CLK(clk),
    .D(_01452_),
    .QN(_00454_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[25]$_DFFE_PP_  (.CLK(clk),
    .D(_01453_),
    .QN(_00453_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[26]$_DFFE_PP_  (.CLK(clk),
    .D(_01454_),
    .QN(_00455_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[27]$_DFFE_PP_  (.CLK(clk),
    .D(_01455_),
    .QN(_00539_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[28]$_DFFE_PP_  (.CLK(clk),
    .D(_01456_),
    .QN(_00538_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[29]$_DFFE_PP_  (.CLK(clk),
    .D(_01457_),
    .QN(_00537_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[2]$_DFFE_PP_  (.CLK(clk),
    .D(_01458_),
    .QN(_00410_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[30]$_DFFE_PP_  (.CLK(clk),
    .D(_01459_),
    .QN(_00536_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[31]$_DFFE_PP_  (.CLK(clk),
    .D(_01460_),
    .QN(_00535_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[32]$_DFFE_PP_  (.CLK(clk),
    .D(_01461_),
    .QN(_00406_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[33]$_DFFE_PP_  (.CLK(clk),
    .D(_01462_),
    .QN(_00405_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[34]$_DFFE_PP_  (.CLK(clk),
    .D(_01463_),
    .QN(_00407_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[35]$_DFFE_PP_  (.CLK(clk),
    .D(_01464_),
    .QN(_00534_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[36]$_DFFE_PP_  (.CLK(clk),
    .D(_01465_),
    .QN(_00533_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[37]$_DFFE_PP_  (.CLK(clk),
    .D(_01466_),
    .QN(_00532_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[38]$_DFFE_PP_  (.CLK(clk),
    .D(_01467_),
    .QN(_00531_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[39]$_DFFE_PP_  (.CLK(clk),
    .D(_01468_),
    .QN(_00530_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[3]$_DFFE_PP_  (.CLK(clk),
    .D(_01469_),
    .QN(_00529_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[40]$_DFFE_PP_  (.CLK(clk),
    .D(_01470_),
    .QN(_00475_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[41]$_DFFE_PP_  (.CLK(clk),
    .D(_01471_),
    .QN(_00474_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[42]$_DFFE_PP_  (.CLK(clk),
    .D(_01472_),
    .QN(_00476_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[43]$_DFFE_PP_  (.CLK(clk),
    .D(_01473_),
    .QN(_00528_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[44]$_DFFE_PP_  (.CLK(clk),
    .D(_01474_),
    .QN(_00527_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[45]$_DFFE_PP_  (.CLK(clk),
    .D(_01475_),
    .QN(_00526_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[46]$_DFFE_PP_  (.CLK(clk),
    .D(_01476_),
    .QN(_00525_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[47]$_DFFE_PP_  (.CLK(clk),
    .D(_01477_),
    .QN(_00524_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[48]$_DFFE_PP_  (.CLK(clk),
    .D(_01478_),
    .QN(_00463_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[49]$_DFFE_PP_  (.CLK(clk),
    .D(_01479_),
    .QN(_00462_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[4]$_DFFE_PP_  (.CLK(clk),
    .D(_01480_),
    .QN(_00523_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[50]$_DFFE_PP_  (.CLK(clk),
    .D(_01481_),
    .QN(_00464_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[51]$_DFFE_PP_  (.CLK(clk),
    .D(_01482_),
    .QN(_00522_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[52]$_DFFE_PP_  (.CLK(clk),
    .D(_01483_),
    .QN(_00521_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[53]$_DFFE_PP_  (.CLK(clk),
    .D(_01484_),
    .QN(_00520_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[54]$_DFFE_PP_  (.CLK(clk),
    .D(_01485_),
    .QN(_00519_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[55]$_DFFE_PP_  (.CLK(clk),
    .D(_01486_),
    .QN(_00518_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[56]$_DFFE_PP_  (.CLK(clk),
    .D(_01487_),
    .QN(_00451_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[57]$_DFFE_PP_  (.CLK(clk),
    .D(_01488_),
    .QN(_00450_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[58]$_DFFE_PP_  (.CLK(clk),
    .D(_01489_),
    .QN(_00452_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[59]$_DFFE_PP_  (.CLK(clk),
    .D(_01490_),
    .QN(_00517_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[5]$_DFFE_PP_  (.CLK(clk),
    .D(_01491_),
    .QN(_00516_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[60]$_DFFE_PP_  (.CLK(clk),
    .D(_01492_),
    .QN(_00515_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[61]$_DFFE_PP_  (.CLK(clk),
    .D(_01493_),
    .QN(_00514_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[62]$_DFFE_PP_  (.CLK(clk),
    .D(_01494_),
    .QN(_00513_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[63]$_DFFE_PP_  (.CLK(clk),
    .D(_01495_),
    .QN(_00512_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[64]$_DFFE_PP_  (.CLK(clk),
    .D(_01496_),
    .QN(_00484_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[65]$_DFFE_PP_  (.CLK(clk),
    .D(_01497_),
    .QN(_00483_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[66]$_DFFE_PP_  (.CLK(clk),
    .D(_01498_),
    .QN(_00485_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[67]$_DFFE_PP_  (.CLK(clk),
    .D(_01499_),
    .QN(_00511_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[68]$_DFFE_PP_  (.CLK(clk),
    .D(_01500_),
    .QN(_00510_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[69]$_DFFE_PP_  (.CLK(clk),
    .D(_01501_),
    .QN(_00509_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[6]$_DFFE_PP_  (.CLK(clk),
    .D(_01502_),
    .QN(_00508_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[70]$_DFFE_PP_  (.CLK(clk),
    .D(_01503_),
    .QN(_00507_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[71]$_DFFE_PP_  (.CLK(clk),
    .D(_01504_),
    .QN(_00506_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[72]$_DFFE_PP_  (.CLK(clk),
    .D(_01505_),
    .QN(_00472_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[73]$_DFFE_PP_  (.CLK(clk),
    .D(_01506_),
    .QN(_00471_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[74]$_DFFE_PP_  (.CLK(clk),
    .D(_01507_),
    .QN(_00473_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[75]$_DFFE_PP_  (.CLK(clk),
    .D(_01508_),
    .QN(_00505_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[76]$_DFFE_PP_  (.CLK(clk),
    .D(_01509_),
    .QN(_00504_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[77]$_DFFE_PP_  (.CLK(clk),
    .D(_01510_),
    .QN(_00503_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[78]$_DFFE_PP_  (.CLK(clk),
    .D(_01511_),
    .QN(_00502_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[79]$_DFFE_PP_  (.CLK(clk),
    .D(_01512_),
    .QN(_00501_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[7]$_DFFE_PP_  (.CLK(clk),
    .D(_01513_),
    .QN(_00500_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[80]$_DFFE_PP_  (.CLK(clk),
    .D(_01514_),
    .QN(_00460_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[81]$_DFFE_PP_  (.CLK(clk),
    .D(_01515_),
    .QN(_00459_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[82]$_DFFE_PP_  (.CLK(clk),
    .D(_01516_),
    .QN(_00461_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[83]$_DFFE_PP_  (.CLK(clk),
    .D(_01517_),
    .QN(_00499_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[84]$_DFFE_PP_  (.CLK(clk),
    .D(_01518_),
    .QN(_00498_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[85]$_DFFE_PP_  (.CLK(clk),
    .D(_01519_),
    .QN(_00497_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[86]$_DFFE_PP_  (.CLK(clk),
    .D(_01520_),
    .QN(_00496_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[87]$_DFFE_PP_  (.CLK(clk),
    .D(_01521_),
    .QN(_00495_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[88]$_DFFE_PP_  (.CLK(clk),
    .D(_01522_),
    .QN(_00448_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[89]$_DFFE_PP_  (.CLK(clk),
    .D(_01523_),
    .QN(_00447_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[8]$_DFFE_PP_  (.CLK(clk),
    .D(_01524_),
    .QN(_00478_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[90]$_DFFE_PP_  (.CLK(clk),
    .D(_01525_),
    .QN(_00449_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[91]$_DFFE_PP_  (.CLK(clk),
    .D(_01526_),
    .QN(_00494_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[92]$_DFFE_PP_  (.CLK(clk),
    .D(_01527_),
    .QN(_00493_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[93]$_DFFE_PP_  (.CLK(clk),
    .D(_01528_),
    .QN(_00492_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[94]$_DFFE_PP_  (.CLK(clk),
    .D(_01529_),
    .QN(_00491_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[95]$_DFFE_PP_  (.CLK(clk),
    .D(_01530_),
    .QN(_00490_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[96]$_DFFE_PP_  (.CLK(clk),
    .D(_01531_),
    .QN(_00481_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[97]$_DFFE_PP_  (.CLK(clk),
    .D(_01532_),
    .QN(_00480_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[98]$_DFFE_PP_  (.CLK(clk),
    .D(_01533_),
    .QN(_00482_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[99]$_DFFE_PP_  (.CLK(clk),
    .D(_01534_),
    .QN(_00489_));
 DFFHQNx1_ASAP7_75t_SL \text_in_r[9]$_DFFE_PP_  (.CLK(clk),
    .D(_01535_),
    .QN(_00477_));
 DFFHQNx1_ASAP7_75t_SL \text_out[0]$_DFF_P_  (.CLK(clk),
    .D(_00265_),
    .QN(_00702_));
 DFFHQNx1_ASAP7_75t_SL \text_out[100]$_DFF_P_  (.CLK(clk),
    .D(_00165_),
    .QN(_00703_));
 DFFHQNx1_ASAP7_75t_SL \text_out[101]$_DFF_P_  (.CLK(clk),
    .D(_00166_),
    .QN(_00704_));
 DFFHQNx1_ASAP7_75t_SL \text_out[102]$_DFF_P_  (.CLK(clk),
    .D(_00167_),
    .QN(_00705_));
 DFFHQNx1_ASAP7_75t_SL \text_out[103]$_DFF_P_  (.CLK(clk),
    .D(_00168_),
    .QN(_00706_));
 DFFHQNx1_ASAP7_75t_SL \text_out[104]$_DFF_P_  (.CLK(clk),
    .D(_00169_),
    .QN(_00707_));
 DFFHQNx1_ASAP7_75t_SL \text_out[105]$_DFF_P_  (.CLK(clk),
    .D(_00170_),
    .QN(_00708_));
 DFFHQNx1_ASAP7_75t_SL \text_out[106]$_DFF_P_  (.CLK(clk),
    .D(_00171_),
    .QN(_00709_));
 DFFHQNx1_ASAP7_75t_SL \text_out[107]$_DFF_P_  (.CLK(clk),
    .D(_00172_),
    .QN(_00710_));
 DFFHQNx1_ASAP7_75t_SL \text_out[108]$_DFF_P_  (.CLK(clk),
    .D(_00173_),
    .QN(_00711_));
 DFFHQNx1_ASAP7_75t_SL \text_out[109]$_DFF_P_  (.CLK(clk),
    .D(_00174_),
    .QN(_00712_));
 DFFHQNx1_ASAP7_75t_SL \text_out[10]$_DFF_P_  (.CLK(clk),
    .D(_00195_),
    .QN(_00713_));
 DFFHQNx1_ASAP7_75t_SL \text_out[110]$_DFF_P_  (.CLK(clk),
    .D(_00175_),
    .QN(_00714_));
 DFFHQNx1_ASAP7_75t_SL \text_out[111]$_DFF_P_  (.CLK(clk),
    .D(_00176_),
    .QN(_00715_));
 DFFHQNx1_ASAP7_75t_SL \text_out[112]$_DFF_P_  (.CLK(clk),
    .D(_00177_),
    .QN(_00716_));
 DFFHQNx1_ASAP7_75t_SL \text_out[113]$_DFF_P_  (.CLK(clk),
    .D(_00178_),
    .QN(_00717_));
 DFFHQNx1_ASAP7_75t_SL \text_out[114]$_DFF_P_  (.CLK(clk),
    .D(_00179_),
    .QN(_00718_));
 DFFHQNx1_ASAP7_75t_SL \text_out[115]$_DFF_P_  (.CLK(clk),
    .D(_00180_),
    .QN(_00719_));
 DFFHQNx1_ASAP7_75t_SL \text_out[116]$_DFF_P_  (.CLK(clk),
    .D(_00181_),
    .QN(_00720_));
 DFFHQNx1_ASAP7_75t_SL \text_out[117]$_DFF_P_  (.CLK(clk),
    .D(_00182_),
    .QN(_00721_));
 DFFHQNx1_ASAP7_75t_SL \text_out[118]$_DFF_P_  (.CLK(clk),
    .D(_00183_),
    .QN(_00722_));
 DFFHQNx1_ASAP7_75t_SL \text_out[119]$_DFF_P_  (.CLK(clk),
    .D(_00184_),
    .QN(_00723_));
 DFFHQNx1_ASAP7_75t_SL \text_out[11]$_DFF_P_  (.CLK(clk),
    .D(_00196_),
    .QN(_00724_));
 DFFHQNx1_ASAP7_75t_SL \text_out[120]$_DFF_P_  (.CLK(clk),
    .D(_00185_),
    .QN(_00725_));
 DFFHQNx1_ASAP7_75t_SL \text_out[121]$_DFF_P_  (.CLK(clk),
    .D(_00186_),
    .QN(_00726_));
 DFFHQNx1_ASAP7_75t_SL \text_out[122]$_DFF_P_  (.CLK(clk),
    .D(_00187_),
    .QN(_00727_));
 DFFHQNx1_ASAP7_75t_SL \text_out[123]$_DFF_P_  (.CLK(clk),
    .D(_00188_),
    .QN(_00728_));
 DFFHQNx1_ASAP7_75t_SL \text_out[124]$_DFF_P_  (.CLK(clk),
    .D(_00189_),
    .QN(_00729_));
 DFFHQNx1_ASAP7_75t_SL \text_out[125]$_DFF_P_  (.CLK(clk),
    .D(_00190_),
    .QN(_00730_));
 DFFHQNx1_ASAP7_75t_SL \text_out[126]$_DFF_P_  (.CLK(clk),
    .D(_00191_),
    .QN(_00731_));
 DFFHQNx1_ASAP7_75t_SL \text_out[127]$_DFF_P_  (.CLK(clk),
    .D(_00192_),
    .QN(_00732_));
 DFFHQNx1_ASAP7_75t_SL \text_out[12]$_DFF_P_  (.CLK(clk),
    .D(_00197_),
    .QN(_00733_));
 DFFHQNx1_ASAP7_75t_SL \text_out[13]$_DFF_P_  (.CLK(clk),
    .D(_00198_),
    .QN(_00734_));
 DFFHQNx1_ASAP7_75t_SL \text_out[14]$_DFF_P_  (.CLK(clk),
    .D(_00199_),
    .QN(_00735_));
 DFFHQNx1_ASAP7_75t_SL \text_out[15]$_DFF_P_  (.CLK(clk),
    .D(_00200_),
    .QN(_00736_));
 DFFHQNx1_ASAP7_75t_SL \text_out[16]$_DFF_P_  (.CLK(clk),
    .D(_00201_),
    .QN(_00737_));
 DFFHQNx1_ASAP7_75t_SL \text_out[17]$_DFF_P_  (.CLK(clk),
    .D(_00202_),
    .QN(_00738_));
 DFFHQNx1_ASAP7_75t_SL \text_out[18]$_DFF_P_  (.CLK(clk),
    .D(_00203_),
    .QN(_00739_));
 DFFHQNx1_ASAP7_75t_SL \text_out[19]$_DFF_P_  (.CLK(clk),
    .D(_00204_),
    .QN(_00740_));
 DFFHQNx1_ASAP7_75t_SL \text_out[1]$_DFF_P_  (.CLK(clk),
    .D(_00266_),
    .QN(_00741_));
 DFFHQNx1_ASAP7_75t_SL \text_out[20]$_DFF_P_  (.CLK(clk),
    .D(_00205_),
    .QN(_00742_));
 DFFHQNx1_ASAP7_75t_SL \text_out[21]$_DFF_P_  (.CLK(clk),
    .D(_00206_),
    .QN(_00743_));
 DFFHQNx1_ASAP7_75t_SL \text_out[22]$_DFF_P_  (.CLK(clk),
    .D(_00207_),
    .QN(_00744_));
 DFFHQNx1_ASAP7_75t_SL \text_out[23]$_DFF_P_  (.CLK(clk),
    .D(_00208_),
    .QN(_00745_));
 DFFHQNx1_ASAP7_75t_SL \text_out[24]$_DFF_P_  (.CLK(clk),
    .D(_00209_),
    .QN(_00746_));
 DFFHQNx1_ASAP7_75t_SL \text_out[25]$_DFF_P_  (.CLK(clk),
    .D(_00210_),
    .QN(_00747_));
 DFFHQNx1_ASAP7_75t_SL \text_out[26]$_DFF_P_  (.CLK(clk),
    .D(_00211_),
    .QN(_00748_));
 DFFHQNx1_ASAP7_75t_SL \text_out[27]$_DFF_P_  (.CLK(clk),
    .D(_00212_),
    .QN(_00749_));
 DFFHQNx1_ASAP7_75t_SL \text_out[28]$_DFF_P_  (.CLK(clk),
    .D(_00213_),
    .QN(_00750_));
 DFFHQNx1_ASAP7_75t_SL \text_out[29]$_DFF_P_  (.CLK(clk),
    .D(_00214_),
    .QN(_00751_));
 DFFHQNx1_ASAP7_75t_SL \text_out[2]$_DFF_P_  (.CLK(clk),
    .D(_00267_),
    .QN(_00752_));
 DFFHQNx1_ASAP7_75t_SL \text_out[30]$_DFF_P_  (.CLK(clk),
    .D(_00215_),
    .QN(_00753_));
 DFFHQNx1_ASAP7_75t_SL \text_out[31]$_DFF_P_  (.CLK(clk),
    .D(_00216_),
    .QN(_00754_));
 DFFHQNx1_ASAP7_75t_SL \text_out[32]$_DFF_P_  (.CLK(clk),
    .D(_00217_),
    .QN(_00755_));
 DFFHQNx1_ASAP7_75t_SL \text_out[33]$_DFF_P_  (.CLK(clk),
    .D(_00218_),
    .QN(_00756_));
 DFFHQNx1_ASAP7_75t_SL \text_out[34]$_DFF_P_  (.CLK(clk),
    .D(_00219_),
    .QN(_00757_));
 DFFHQNx1_ASAP7_75t_SL \text_out[35]$_DFF_P_  (.CLK(clk),
    .D(_00220_),
    .QN(_00758_));
 DFFHQNx1_ASAP7_75t_SL \text_out[36]$_DFF_P_  (.CLK(clk),
    .D(_00221_),
    .QN(_00759_));
 DFFHQNx1_ASAP7_75t_SL \text_out[37]$_DFF_P_  (.CLK(clk),
    .D(_00222_),
    .QN(_00760_));
 DFFHQNx1_ASAP7_75t_SL \text_out[38]$_DFF_P_  (.CLK(clk),
    .D(_00223_),
    .QN(_00761_));
 DFFHQNx1_ASAP7_75t_SL \text_out[39]$_DFF_P_  (.CLK(clk),
    .D(_00224_),
    .QN(_00762_));
 DFFHQNx1_ASAP7_75t_SL \text_out[3]$_DFF_P_  (.CLK(clk),
    .D(_00268_),
    .QN(_00763_));
 DFFHQNx1_ASAP7_75t_SL \text_out[40]$_DFF_P_  (.CLK(clk),
    .D(_00225_),
    .QN(_00764_));
 DFFHQNx1_ASAP7_75t_SL \text_out[41]$_DFF_P_  (.CLK(clk),
    .D(_00226_),
    .QN(_00765_));
 DFFHQNx1_ASAP7_75t_SL \text_out[42]$_DFF_P_  (.CLK(clk),
    .D(_00227_),
    .QN(_00766_));
 DFFHQNx1_ASAP7_75t_SL \text_out[43]$_DFF_P_  (.CLK(clk),
    .D(_00228_),
    .QN(_00767_));
 DFFHQNx1_ASAP7_75t_SL \text_out[44]$_DFF_P_  (.CLK(clk),
    .D(_00229_),
    .QN(_00768_));
 DFFHQNx1_ASAP7_75t_SL \text_out[45]$_DFF_P_  (.CLK(clk),
    .D(_00230_),
    .QN(_00769_));
 DFFHQNx1_ASAP7_75t_SL \text_out[46]$_DFF_P_  (.CLK(clk),
    .D(_00231_),
    .QN(_00770_));
 DFFHQNx1_ASAP7_75t_SL \text_out[47]$_DFF_P_  (.CLK(clk),
    .D(_00232_),
    .QN(_00771_));
 DFFHQNx1_ASAP7_75t_SL \text_out[48]$_DFF_P_  (.CLK(clk),
    .D(_00233_),
    .QN(_00772_));
 DFFHQNx1_ASAP7_75t_SL \text_out[49]$_DFF_P_  (.CLK(clk),
    .D(_00234_),
    .QN(_00773_));
 DFFHQNx1_ASAP7_75t_SL \text_out[4]$_DFF_P_  (.CLK(clk),
    .D(_00269_),
    .QN(_00774_));
 DFFHQNx1_ASAP7_75t_SL \text_out[50]$_DFF_P_  (.CLK(clk),
    .D(_00235_),
    .QN(_00775_));
 DFFHQNx1_ASAP7_75t_SL \text_out[51]$_DFF_P_  (.CLK(clk),
    .D(_00236_),
    .QN(_00776_));
 DFFHQNx1_ASAP7_75t_SL \text_out[52]$_DFF_P_  (.CLK(clk),
    .D(_00237_),
    .QN(_00777_));
 DFFHQNx1_ASAP7_75t_SL \text_out[53]$_DFF_P_  (.CLK(clk),
    .D(_00238_),
    .QN(_00778_));
 DFFHQNx1_ASAP7_75t_SL \text_out[54]$_DFF_P_  (.CLK(clk),
    .D(_00239_),
    .QN(_00779_));
 DFFHQNx1_ASAP7_75t_SL \text_out[55]$_DFF_P_  (.CLK(clk),
    .D(_00240_),
    .QN(_00780_));
 DFFHQNx1_ASAP7_75t_SL \text_out[56]$_DFF_P_  (.CLK(clk),
    .D(_00241_),
    .QN(_00781_));
 DFFHQNx1_ASAP7_75t_SL \text_out[57]$_DFF_P_  (.CLK(clk),
    .D(_00242_),
    .QN(_00782_));
 DFFHQNx1_ASAP7_75t_SL \text_out[58]$_DFF_P_  (.CLK(clk),
    .D(_00243_),
    .QN(_00783_));
 DFFHQNx1_ASAP7_75t_SL \text_out[59]$_DFF_P_  (.CLK(clk),
    .D(_00244_),
    .QN(_00784_));
 DFFHQNx1_ASAP7_75t_SL \text_out[5]$_DFF_P_  (.CLK(clk),
    .D(_00270_),
    .QN(_00785_));
 DFFHQNx1_ASAP7_75t_SL \text_out[60]$_DFF_P_  (.CLK(clk),
    .D(_00245_),
    .QN(_00786_));
 DFFHQNx1_ASAP7_75t_SL \text_out[61]$_DFF_P_  (.CLK(clk),
    .D(_00246_),
    .QN(_00787_));
 DFFHQNx1_ASAP7_75t_SL \text_out[62]$_DFF_P_  (.CLK(clk),
    .D(_00247_),
    .QN(_00788_));
 DFFHQNx1_ASAP7_75t_SL \text_out[63]$_DFF_P_  (.CLK(clk),
    .D(_00248_),
    .QN(_00789_));
 DFFHQNx1_ASAP7_75t_SL \text_out[64]$_DFF_P_  (.CLK(clk),
    .D(_00249_),
    .QN(_00790_));
 DFFHQNx1_ASAP7_75t_SL \text_out[65]$_DFF_P_  (.CLK(clk),
    .D(_00250_),
    .QN(_00791_));
 DFFHQNx1_ASAP7_75t_SL \text_out[66]$_DFF_P_  (.CLK(clk),
    .D(_00251_),
    .QN(_00792_));
 DFFHQNx1_ASAP7_75t_SL \text_out[67]$_DFF_P_  (.CLK(clk),
    .D(_00252_),
    .QN(_00793_));
 DFFHQNx1_ASAP7_75t_SL \text_out[68]$_DFF_P_  (.CLK(clk),
    .D(_00253_),
    .QN(_00794_));
 DFFHQNx1_ASAP7_75t_SL \text_out[69]$_DFF_P_  (.CLK(clk),
    .D(_00254_),
    .QN(_00795_));
 DFFHQNx1_ASAP7_75t_SL \text_out[6]$_DFF_P_  (.CLK(clk),
    .D(_00271_),
    .QN(_00796_));
 DFFHQNx1_ASAP7_75t_SL \text_out[70]$_DFF_P_  (.CLK(clk),
    .D(_00255_),
    .QN(_00797_));
 DFFHQNx1_ASAP7_75t_SL \text_out[71]$_DFF_P_  (.CLK(clk),
    .D(_00256_),
    .QN(_00798_));
 DFFHQNx1_ASAP7_75t_SL \text_out[72]$_DFF_P_  (.CLK(clk),
    .D(_00257_),
    .QN(_00799_));
 DFFHQNx1_ASAP7_75t_SL \text_out[73]$_DFF_P_  (.CLK(clk),
    .D(_00258_),
    .QN(_00800_));
 DFFHQNx1_ASAP7_75t_SL \text_out[74]$_DFF_P_  (.CLK(clk),
    .D(_00259_),
    .QN(_00801_));
 DFFHQNx1_ASAP7_75t_SL \text_out[75]$_DFF_P_  (.CLK(clk),
    .D(_00260_),
    .QN(_00802_));
 DFFHQNx1_ASAP7_75t_SL \text_out[76]$_DFF_P_  (.CLK(clk),
    .D(_00261_),
    .QN(_00803_));
 DFFHQNx1_ASAP7_75t_SL \text_out[77]$_DFF_P_  (.CLK(clk),
    .D(_00262_),
    .QN(_00804_));
 DFFHQNx1_ASAP7_75t_SL \text_out[78]$_DFF_P_  (.CLK(clk),
    .D(_00263_),
    .QN(_00805_));
 DFFHQNx1_ASAP7_75t_SL \text_out[79]$_DFF_P_  (.CLK(clk),
    .D(_00264_),
    .QN(_00806_));
 DFFHQNx1_ASAP7_75t_SL \text_out[7]$_DFF_P_  (.CLK(clk),
    .D(_00272_),
    .QN(_00807_));
 DFFHQNx1_ASAP7_75t_SL \text_out[80]$_DFF_P_  (.CLK(clk),
    .D(_00273_),
    .QN(_00808_));
 DFFHQNx1_ASAP7_75t_SL \text_out[81]$_DFF_P_  (.CLK(clk),
    .D(_00274_),
    .QN(_00809_));
 DFFHQNx1_ASAP7_75t_SL \text_out[82]$_DFF_P_  (.CLK(clk),
    .D(_00275_),
    .QN(_00810_));
 DFFHQNx1_ASAP7_75t_SL \text_out[83]$_DFF_P_  (.CLK(clk),
    .D(_00276_),
    .QN(_00811_));
 DFFHQNx1_ASAP7_75t_SL \text_out[84]$_DFF_P_  (.CLK(clk),
    .D(_00277_),
    .QN(_00812_));
 DFFHQNx1_ASAP7_75t_SL \text_out[85]$_DFF_P_  (.CLK(clk),
    .D(_00278_),
    .QN(_00813_));
 DFFHQNx1_ASAP7_75t_SL \text_out[86]$_DFF_P_  (.CLK(clk),
    .D(_00279_),
    .QN(_00814_));
 DFFHQNx1_ASAP7_75t_SL \text_out[87]$_DFF_P_  (.CLK(clk),
    .D(_00280_),
    .QN(_00815_));
 DFFHQNx1_ASAP7_75t_SL \text_out[88]$_DFF_P_  (.CLK(clk),
    .D(_00281_),
    .QN(_00816_));
 DFFHQNx1_ASAP7_75t_SL \text_out[89]$_DFF_P_  (.CLK(clk),
    .D(_00282_),
    .QN(_00817_));
 DFFHQNx1_ASAP7_75t_SL \text_out[8]$_DFF_P_  (.CLK(clk),
    .D(_00193_),
    .QN(_00818_));
 DFFHQNx1_ASAP7_75t_SL \text_out[90]$_DFF_P_  (.CLK(clk),
    .D(_00283_),
    .QN(_00819_));
 DFFHQNx1_ASAP7_75t_SL \text_out[91]$_DFF_P_  (.CLK(clk),
    .D(_00284_),
    .QN(_00820_));
 DFFHQNx1_ASAP7_75t_SL \text_out[92]$_DFF_P_  (.CLK(clk),
    .D(_00285_),
    .QN(_00821_));
 DFFHQNx1_ASAP7_75t_SL \text_out[93]$_DFF_P_  (.CLK(clk),
    .D(_00286_),
    .QN(_00822_));
 DFFHQNx1_ASAP7_75t_SL \text_out[94]$_DFF_P_  (.CLK(clk),
    .D(_00287_),
    .QN(_00823_));
 DFFHQNx1_ASAP7_75t_SL \text_out[95]$_DFF_P_  (.CLK(clk),
    .D(_00288_),
    .QN(_00824_));
 DFFHQNx1_ASAP7_75t_SL \text_out[96]$_DFF_P_  (.CLK(clk),
    .D(_00161_),
    .QN(_00825_));
 DFFHQNx1_ASAP7_75t_SL \text_out[97]$_DFF_P_  (.CLK(clk),
    .D(_00162_),
    .QN(_00826_));
 DFFHQNx1_ASAP7_75t_SL \text_out[98]$_DFF_P_  (.CLK(clk),
    .D(_00163_),
    .QN(_00827_));
 DFFHQNx1_ASAP7_75t_SL \text_out[99]$_DFF_P_  (.CLK(clk),
    .D(_00164_),
    .QN(_00828_));
 DFFHQNx1_ASAP7_75t_SL \text_out[9]$_DFF_P_  (.CLK(clk),
    .D(_00194_),
    .QN(_00488_));
 DFFHQNx1_ASAP7_75t_SL \u0.r0.out[24]$_SDFF_PP1_  (.CLK(clk),
    .D(_01536_),
    .QN(_00413_));
 DFFHQNx1_ASAP7_75t_SL \u0.r0.out[25]$_SDFF_PP0_  (.CLK(clk),
    .D(_01537_),
    .QN(_00414_));
 DFFHQNx1_ASAP7_75t_SL \u0.r0.out[26]$_SDFF_PP0_  (.CLK(clk),
    .D(_01538_),
    .QN(_00415_));
 DFFHQNx1_ASAP7_75t_SL \u0.r0.out[27]$_SDFF_PP0_  (.CLK(clk),
    .D(_01539_),
    .QN(_00416_));
 DFFHQNx1_ASAP7_75t_SL \u0.r0.out[28]$_SDFF_PP0_  (.CLK(clk),
    .D(_01540_),
    .QN(_00417_));
 DFFHQNx1_ASAP7_75t_SL \u0.r0.out[29]$_SDFF_PP0_  (.CLK(clk),
    .D(_01541_),
    .QN(_00418_));
 DFFHQNx1_ASAP7_75t_SL \u0.r0.out[30]$_SDFF_PP0_  (.CLK(clk),
    .D(_01542_),
    .QN(_00419_));
 DFFHQNx1_ASAP7_75t_SL \u0.r0.out[31]$_SDFF_PP0_  (.CLK(clk),
    .D(_01543_),
    .QN(_00420_));
 DFFHQNx1_ASAP7_75t_SL \u0.r0.rcnt[0]$_SDFF_PP0_  (.CLK(clk),
    .D(_01544_),
    .QN(\u0.r0.rcnt_next[0] ));
 DFFHQNx1_ASAP7_75t_SL \u0.r0.rcnt[1]$_SDFF_PP0_  (.CLK(clk),
    .D(_01545_),
    .QN(_00965_));
 DFFHQNx1_ASAP7_75t_SL \u0.r0.rcnt[2]$_SDFF_PP0_  (.CLK(clk),
    .D(_01546_),
    .QN(_00487_));
 DFFHQNx1_ASAP7_75t_SL \u0.r0.rcnt[3]$_SDFF_PP0_  (.CLK(clk),
    .D(_01547_),
    .QN(_00829_));
 DFFHQNx1_ASAP7_75t_SL \u0.u0.d[0]$_DFF_P_  (.CLK(clk),
    .D(_00000_),
    .QN(_00830_));
 DFFHQNx1_ASAP7_75t_SL \u0.u0.d[1]$_DFF_P_  (.CLK(clk),
    .D(_00001_),
    .QN(_00831_));
 DFFHQNx1_ASAP7_75t_SL \u0.u0.d[2]$_DFF_P_  (.CLK(clk),
    .D(_00002_),
    .QN(_00832_));
 DFFHQNx1_ASAP7_75t_SL \u0.u0.d[3]$_DFF_P_  (.CLK(clk),
    .D(_00003_),
    .QN(_00833_));
 DFFHQNx1_ASAP7_75t_SL \u0.u0.d[4]$_DFF_P_  (.CLK(clk),
    .D(_00004_),
    .QN(_00834_));
 DFFHQNx1_ASAP7_75t_SL \u0.u0.d[5]$_DFF_P_  (.CLK(clk),
    .D(_00005_),
    .QN(_00835_));
 DFFHQNx1_ASAP7_75t_SL \u0.u0.d[6]$_DFF_P_  (.CLK(clk),
    .D(_00006_),
    .QN(_00836_));
 DFFHQNx1_ASAP7_75t_SL \u0.u0.d[7]$_DFF_P_  (.CLK(clk),
    .D(_00007_),
    .QN(_00837_));
 DFFHQNx1_ASAP7_75t_SL \u0.u1.d[0]$_DFF_P_  (.CLK(clk),
    .D(_00008_),
    .QN(_00437_));
 DFFHQNx1_ASAP7_75t_SL \u0.u1.d[1]$_DFF_P_  (.CLK(clk),
    .D(_00009_),
    .QN(_00438_));
 DFFHQNx1_ASAP7_75t_SL \u0.u1.d[2]$_DFF_P_  (.CLK(clk),
    .D(_00010_),
    .QN(_00412_));
 DFFHQNx1_ASAP7_75t_SL \u0.u1.d[3]$_DFF_P_  (.CLK(clk),
    .D(_00011_),
    .QN(_00439_));
 DFFHQNx1_ASAP7_75t_SL \u0.u1.d[4]$_DFF_P_  (.CLK(clk),
    .D(_00012_),
    .QN(_00440_));
 DFFHQNx1_ASAP7_75t_SL \u0.u1.d[5]$_DFF_P_  (.CLK(clk),
    .D(_00013_),
    .QN(_00441_));
 DFFHQNx1_ASAP7_75t_SL \u0.u1.d[6]$_DFF_P_  (.CLK(clk),
    .D(_00014_),
    .QN(_00442_));
 DFFHQNx1_ASAP7_75t_SL \u0.u1.d[7]$_DFF_P_  (.CLK(clk),
    .D(_00015_),
    .QN(_00443_));
 DFFHQNx1_ASAP7_75t_SL \u0.u2.d[0]$_DFF_P_  (.CLK(clk),
    .D(_00016_),
    .QN(_00429_));
 DFFHQNx1_ASAP7_75t_SL \u0.u2.d[1]$_DFF_P_  (.CLK(clk),
    .D(_00017_),
    .QN(_00430_));
 DFFHQNx1_ASAP7_75t_SL \u0.u2.d[2]$_DFF_P_  (.CLK(clk),
    .D(_00018_),
    .QN(_00431_));
 DFFHQNx1_ASAP7_75t_SL \u0.u2.d[3]$_DFF_P_  (.CLK(clk),
    .D(_00019_),
    .QN(_00432_));
 DFFHQNx1_ASAP7_75t_SL \u0.u2.d[4]$_DFF_P_  (.CLK(clk),
    .D(_00020_),
    .QN(_00433_));
 DFFHQNx1_ASAP7_75t_SL \u0.u2.d[5]$_DFF_P_  (.CLK(clk),
    .D(_00021_),
    .QN(_00434_));
 DFFHQNx1_ASAP7_75t_SL \u0.u2.d[6]$_DFF_P_  (.CLK(clk),
    .D(_00022_),
    .QN(_00435_));
 DFFHQNx1_ASAP7_75t_SL \u0.u2.d[7]$_DFF_P_  (.CLK(clk),
    .D(_00023_),
    .QN(_00436_));
 DFFHQNx1_ASAP7_75t_SL \u0.u3.d[0]$_DFF_P_  (.CLK(clk),
    .D(_00024_),
    .QN(_00421_));
 DFFHQNx1_ASAP7_75t_SL \u0.u3.d[1]$_DFF_P_  (.CLK(clk),
    .D(_00025_),
    .QN(_00422_));
 DFFHQNx1_ASAP7_75t_SL \u0.u3.d[2]$_DFF_P_  (.CLK(clk),
    .D(_00026_),
    .QN(_00423_));
 DFFHQNx1_ASAP7_75t_SL \u0.u3.d[3]$_DFF_P_  (.CLK(clk),
    .D(_00027_),
    .QN(_00424_));
 DFFHQNx1_ASAP7_75t_SL \u0.u3.d[4]$_DFF_P_  (.CLK(clk),
    .D(_00028_),
    .QN(_00425_));
 DFFHQNx1_ASAP7_75t_SL \u0.u3.d[5]$_DFF_P_  (.CLK(clk),
    .D(_00029_),
    .QN(_00426_));
 DFFHQNx1_ASAP7_75t_SL \u0.u3.d[6]$_DFF_P_  (.CLK(clk),
    .D(_00030_),
    .QN(_00427_));
 DFFHQNx1_ASAP7_75t_SL \u0.u3.d[7]$_DFF_P_  (.CLK(clk),
    .D(_00031_),
    .QN(_00428_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][0]$_DFF_P_  (.CLK(clk),
    .D(_00289_),
    .QN(_00838_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][10]$_DFF_P_  (.CLK(clk),
    .D(_00290_),
    .QN(_00839_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][11]$_DFF_P_  (.CLK(clk),
    .D(_00291_),
    .QN(_00840_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][12]$_DFF_P_  (.CLK(clk),
    .D(_00292_),
    .QN(_00841_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][13]$_DFF_P_  (.CLK(clk),
    .D(_00293_),
    .QN(_00842_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][14]$_DFF_P_  (.CLK(clk),
    .D(_00294_),
    .QN(_00843_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][15]$_DFF_P_  (.CLK(clk),
    .D(_00295_),
    .QN(_00844_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][16]$_DFF_P_  (.CLK(clk),
    .D(_00296_),
    .QN(_00845_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][17]$_DFF_P_  (.CLK(clk),
    .D(_00297_),
    .QN(_00846_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][18]$_DFF_P_  (.CLK(clk),
    .D(_00298_),
    .QN(_00847_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][19]$_DFF_P_  (.CLK(clk),
    .D(_00299_),
    .QN(_00848_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][1]$_DFF_P_  (.CLK(clk),
    .D(_00300_),
    .QN(_00849_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][20]$_DFF_P_  (.CLK(clk),
    .D(_00301_),
    .QN(_00850_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][21]$_DFF_P_  (.CLK(clk),
    .D(_00302_),
    .QN(_00851_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][22]$_DFF_P_  (.CLK(clk),
    .D(_00303_),
    .QN(_00852_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][23]$_DFF_P_  (.CLK(clk),
    .D(_00304_),
    .QN(_00853_));
 DFFHQNx2_ASAP7_75t_SL \u0.w[0][24]$_DFF_P_  (.CLK(clk),
    .D(_00305_),
    .QN(_00854_));
 DFFHQNx2_ASAP7_75t_SL \u0.w[0][25]$_DFF_P_  (.CLK(clk),
    .D(_00306_),
    .QN(_00855_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][26]$_DFF_P_  (.CLK(clk),
    .D(_00307_),
    .QN(_00856_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][27]$_DFF_P_  (.CLK(clk),
    .D(_00308_),
    .QN(_00857_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][28]$_DFF_P_  (.CLK(clk),
    .D(_00309_),
    .QN(_00858_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][29]$_DFF_P_  (.CLK(clk),
    .D(_00310_),
    .QN(_00859_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][2]$_DFF_P_  (.CLK(clk),
    .D(_00311_),
    .QN(_00860_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][30]$_DFF_P_  (.CLK(clk),
    .D(_00312_),
    .QN(_00861_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][31]$_DFF_P_  (.CLK(clk),
    .D(_00313_),
    .QN(_00862_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][3]$_DFF_P_  (.CLK(clk),
    .D(_00314_),
    .QN(_00863_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][4]$_DFF_P_  (.CLK(clk),
    .D(_00315_),
    .QN(_00864_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][5]$_DFF_P_  (.CLK(clk),
    .D(_00316_),
    .QN(_00865_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][6]$_DFF_P_  (.CLK(clk),
    .D(_00317_),
    .QN(_00866_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][7]$_DFF_P_  (.CLK(clk),
    .D(_00318_),
    .QN(_00867_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][8]$_DFF_P_  (.CLK(clk),
    .D(_00319_),
    .QN(_00868_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[0][9]$_DFF_P_  (.CLK(clk),
    .D(_00320_),
    .QN(_00869_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][0]$_DFF_P_  (.CLK(clk),
    .D(_00321_),
    .QN(_00870_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][10]$_DFF_P_  (.CLK(clk),
    .D(_00322_),
    .QN(_00871_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][11]$_DFF_P_  (.CLK(clk),
    .D(_00323_),
    .QN(_00872_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][12]$_DFF_P_  (.CLK(clk),
    .D(_00324_),
    .QN(_00873_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][13]$_DFF_P_  (.CLK(clk),
    .D(_00325_),
    .QN(_00874_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][14]$_DFF_P_  (.CLK(clk),
    .D(_00326_),
    .QN(_00875_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][15]$_DFF_P_  (.CLK(clk),
    .D(_00327_),
    .QN(_00876_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][16]$_DFF_P_  (.CLK(clk),
    .D(_00328_),
    .QN(_00877_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][17]$_DFF_P_  (.CLK(clk),
    .D(_00329_),
    .QN(_00878_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][18]$_DFF_P_  (.CLK(clk),
    .D(_00330_),
    .QN(_00879_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][19]$_DFF_P_  (.CLK(clk),
    .D(_00331_),
    .QN(_00880_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][1]$_DFF_P_  (.CLK(clk),
    .D(_00332_),
    .QN(_00881_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][20]$_DFF_P_  (.CLK(clk),
    .D(_00333_),
    .QN(_00882_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][21]$_DFF_P_  (.CLK(clk),
    .D(_00334_),
    .QN(_00883_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][22]$_DFF_P_  (.CLK(clk),
    .D(_00335_),
    .QN(_00884_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][23]$_DFF_P_  (.CLK(clk),
    .D(_00336_),
    .QN(_00885_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][24]$_DFF_P_  (.CLK(clk),
    .D(_00337_),
    .QN(_00886_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][25]$_DFF_P_  (.CLK(clk),
    .D(_00338_),
    .QN(_00887_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][26]$_DFF_P_  (.CLK(clk),
    .D(_00339_),
    .QN(_00888_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][27]$_DFF_P_  (.CLK(clk),
    .D(_00340_),
    .QN(_00889_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][28]$_DFF_P_  (.CLK(clk),
    .D(_00341_),
    .QN(_00890_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][29]$_DFF_P_  (.CLK(clk),
    .D(_00342_),
    .QN(_00891_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][2]$_DFF_P_  (.CLK(clk),
    .D(_00343_),
    .QN(_00892_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][30]$_DFF_P_  (.CLK(clk),
    .D(_00344_),
    .QN(_00893_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][31]$_DFF_P_  (.CLK(clk),
    .D(_00345_),
    .QN(_00894_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][3]$_DFF_P_  (.CLK(clk),
    .D(_00346_),
    .QN(_00895_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][4]$_DFF_P_  (.CLK(clk),
    .D(_00347_),
    .QN(_00896_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][5]$_DFF_P_  (.CLK(clk),
    .D(_00348_),
    .QN(_00897_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][6]$_DFF_P_  (.CLK(clk),
    .D(_00349_),
    .QN(_00898_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][7]$_DFF_P_  (.CLK(clk),
    .D(_00350_),
    .QN(_00899_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][8]$_DFF_P_  (.CLK(clk),
    .D(_00351_),
    .QN(_00900_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[1][9]$_DFF_P_  (.CLK(clk),
    .D(_00352_),
    .QN(_00901_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][0]$_DFF_P_  (.CLK(clk),
    .D(_00353_),
    .QN(_00902_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][10]$_DFF_P_  (.CLK(clk),
    .D(_00354_),
    .QN(_00903_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][11]$_DFF_P_  (.CLK(clk),
    .D(_00355_),
    .QN(_00904_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][12]$_DFF_P_  (.CLK(clk),
    .D(_00356_),
    .QN(_00905_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][13]$_DFF_P_  (.CLK(clk),
    .D(_00357_),
    .QN(_00906_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][14]$_DFF_P_  (.CLK(clk),
    .D(_00358_),
    .QN(_00907_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][15]$_DFF_P_  (.CLK(clk),
    .D(_00359_),
    .QN(_00908_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][16]$_DFF_P_  (.CLK(clk),
    .D(_00360_),
    .QN(_00909_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][17]$_DFF_P_  (.CLK(clk),
    .D(_00361_),
    .QN(_00910_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][18]$_DFF_P_  (.CLK(clk),
    .D(_00362_),
    .QN(_00911_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][19]$_DFF_P_  (.CLK(clk),
    .D(_00363_),
    .QN(_00912_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][1]$_DFF_P_  (.CLK(clk),
    .D(_00364_),
    .QN(_00913_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][20]$_DFF_P_  (.CLK(clk),
    .D(_00365_),
    .QN(_00914_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][21]$_DFF_P_  (.CLK(clk),
    .D(_00366_),
    .QN(_00915_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][22]$_DFF_P_  (.CLK(clk),
    .D(_00367_),
    .QN(_00916_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][23]$_DFF_P_  (.CLK(clk),
    .D(_00368_),
    .QN(_00917_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][24]$_DFF_P_  (.CLK(clk),
    .D(_00369_),
    .QN(_00918_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][25]$_DFF_P_  (.CLK(clk),
    .D(_00370_),
    .QN(_00919_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][26]$_DFF_P_  (.CLK(clk),
    .D(_00371_),
    .QN(_00920_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][27]$_DFF_P_  (.CLK(clk),
    .D(_00372_),
    .QN(_00921_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][28]$_DFF_P_  (.CLK(clk),
    .D(_00373_),
    .QN(_00922_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][29]$_DFF_P_  (.CLK(clk),
    .D(_00374_),
    .QN(_00923_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][2]$_DFF_P_  (.CLK(clk),
    .D(_00375_),
    .QN(_00924_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][30]$_DFF_P_  (.CLK(clk),
    .D(_00376_),
    .QN(_00925_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][31]$_DFF_P_  (.CLK(clk),
    .D(_00377_),
    .QN(_00926_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][3]$_DFF_P_  (.CLK(clk),
    .D(_00378_),
    .QN(_00927_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][4]$_DFF_P_  (.CLK(clk),
    .D(_00379_),
    .QN(_00928_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][5]$_DFF_P_  (.CLK(clk),
    .D(_00380_),
    .QN(_00929_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][6]$_DFF_P_  (.CLK(clk),
    .D(_00381_),
    .QN(_00930_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][7]$_DFF_P_  (.CLK(clk),
    .D(_00382_),
    .QN(_00931_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][8]$_DFF_P_  (.CLK(clk),
    .D(_00383_),
    .QN(_00932_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[2][9]$_DFF_P_  (.CLK(clk),
    .D(_00384_),
    .QN(_00933_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][0]$_DFF_P_  (.CLK(clk),
    .D(_09557_),
    .QN(_00934_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][10]$_DFF_P_  (.CLK(clk),
    .D(_08919_),
    .QN(_00935_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][11]$_DFF_P_  (.CLK(clk),
    .D(_08925_),
    .QN(_00936_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][12]$_DFF_P_  (.CLK(clk),
    .D(_08929_),
    .QN(_00937_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][13]$_DFF_P_  (.CLK(clk),
    .D(_08934_),
    .QN(_00938_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][14]$_DFF_P_  (.CLK(clk),
    .D(_08938_),
    .QN(_00939_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][15]$_DFF_P_  (.CLK(clk),
    .D(_08941_),
    .QN(_00940_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][16]$_DFF_P_  (.CLK(clk),
    .D(_00973_),
    .QN(_00941_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][17]$_DFF_P_  (.CLK(clk),
    .D(_00972_),
    .QN(_00942_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][18]$_DFF_P_  (.CLK(clk),
    .D(_00989_),
    .QN(_00943_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][19]$_DFF_P_  (.CLK(clk),
    .D(_08037_),
    .QN(_00944_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][1]$_DFF_P_  (.CLK(clk),
    .D(_09554_),
    .QN(_00945_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][20]$_DFF_P_  (.CLK(clk),
    .D(_08020_),
    .QN(_00946_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][21]$_DFF_P_  (.CLK(clk),
    .D(_08028_),
    .QN(_00947_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][22]$_DFF_P_  (.CLK(clk),
    .D(_08071_),
    .QN(_00948_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][23]$_DFF_P_  (.CLK(clk),
    .D(_08078_),
    .QN(_00949_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][24]$_DFF_P_  (.CLK(clk),
    .D(_10110_),
    .QN(_00950_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][25]$_DFF_P_  (.CLK(clk),
    .D(_10103_),
    .QN(_00951_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][26]$_DFF_P_  (.CLK(clk),
    .D(_10104_),
    .QN(_00952_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][27]$_DFF_P_  (.CLK(clk),
    .D(_08968_),
    .QN(_00953_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][28]$_DFF_P_  (.CLK(clk),
    .D(_08976_),
    .QN(_00954_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][29]$_DFF_P_  (.CLK(clk),
    .D(_08982_),
    .QN(_00955_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][2]$_DFF_P_  (.CLK(clk),
    .D(_08879_),
    .QN(_00956_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][30]$_DFF_P_  (.CLK(clk),
    .D(_08988_),
    .QN(_00957_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][31]$_DFF_P_  (.CLK(clk),
    .D(_08992_),
    .QN(_00958_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][3]$_DFF_P_  (.CLK(clk),
    .D(_08885_),
    .QN(_00959_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][4]$_DFF_P_  (.CLK(clk),
    .D(_08890_),
    .QN(_00960_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][5]$_DFF_P_  (.CLK(clk),
    .D(_08894_),
    .QN(_00961_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][6]$_DFF_P_  (.CLK(clk),
    .D(_08899_),
    .QN(_00962_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][7]$_DFF_P_  (.CLK(clk),
    .D(_08902_),
    .QN(_00963_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][8]$_DFF_P_  (.CLK(clk),
    .D(_08995_),
    .QN(_00964_));
 DFFHQNx1_ASAP7_75t_SL \u0.w[3][9]$_DFF_P_  (.CLK(clk),
    .D(_00994_),
    .QN(_00486_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_Right_170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_Right_171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_Right_172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_Right_173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_Right_174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_Right_175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_Right_176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_Right_177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_Right_178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_Right_179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_Right_180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_Right_181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_Right_182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_Right_183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_Right_184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_Right_185 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_Right_186 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_Right_187 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_Right_188 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_Right_189 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_Right_190 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_Right_191 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_Right_192 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_Right_193 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_Right_194 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_Right_195 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_Right_196 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_Right_197 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_Right_198 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_Right_199 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_Right_200 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_Right_201 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_Right_202 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_Right_203 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_Right_204 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_Right_205 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_Right_206 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_Right_207 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_Right_208 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_Right_209 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_Right_210 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_Right_211 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_Right_212 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_Right_213 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_Right_214 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_Right_215 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_Right_216 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_Right_217 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_Right_218 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_Right_219 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_Right_220 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_Right_221 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_Right_222 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_Right_223 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_Right_224 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_Right_225 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_Right_226 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_Right_227 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_Right_228 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_Right_229 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_Right_230 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_Right_231 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_Right_232 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_Right_233 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_Right_234 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_Right_235 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_Right_236 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_Right_237 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_Right_238 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_Right_239 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_240 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_241 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_242 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_243 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_244 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_245 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_246 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_247 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_248 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_249 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_250 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_251 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_252 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_253 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_254 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_255 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_256 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_257 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_258 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_259 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_260 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_261 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_262 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_263 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_264 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_265 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_266 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_267 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_268 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_269 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_270 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_271 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_272 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_273 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_274 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_275 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_276 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_277 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_278 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_279 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_280 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_281 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_282 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_283 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_284 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_285 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_286 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_287 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Left_288 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Left_289 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Left_290 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Left_291 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Left_292 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Left_293 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Left_294 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Left_295 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Left_296 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Left_297 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Left_298 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Left_299 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Left_300 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Left_301 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_Left_302 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_Left_303 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_Left_304 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_Left_305 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_Left_306 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_Left_307 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_Left_308 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_Left_309 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_Left_310 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_Left_311 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_Left_312 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_Left_313 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_Left_314 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_Left_315 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_Left_316 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_Left_317 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_Left_318 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_Left_319 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_Left_320 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_Left_321 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_Left_322 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_Left_323 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_Left_324 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_Left_325 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_Left_326 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_Left_327 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_Left_328 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_Left_329 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_Left_330 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_Left_331 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_Left_332 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_Left_333 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_Left_334 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_Left_335 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_Left_336 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_Left_337 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_Left_338 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_Left_339 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_Left_340 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_Left_341 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_Left_342 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_Left_343 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_Left_344 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_Left_345 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_Left_346 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_Left_347 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_Left_348 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_Left_349 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_Left_350 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_Left_351 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_Left_352 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_Left_353 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_Left_354 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_Left_355 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_Left_356 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_Left_357 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_Left_358 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_Left_359 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_Left_360 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_Left_361 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_Left_362 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_Left_363 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_Left_364 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_Left_365 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_Left_366 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_Left_367 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_Left_368 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_Left_369 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_Left_370 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_Left_371 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_Left_372 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_Left_373 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_Left_374 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_Left_375 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_Left_376 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_Left_377 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_Left_378 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_Left_379 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_Left_380 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_Left_381 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_Left_382 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_Left_383 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_Left_384 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_Left_385 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_Left_386 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_Left_387 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_Left_388 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_Left_389 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_Left_390 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_Left_391 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_Left_392 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_Left_393 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_Left_394 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_Left_395 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_Left_396 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_Left_397 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_Left_398 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_Left_399 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_Left_400 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_Left_401 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_Left_402 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_Left_403 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_Left_404 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_Left_405 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_Left_406 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_Left_407 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_Left_408 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_Left_409 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_Left_410 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_Left_411 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_Left_412 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_Left_413 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_Left_414 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_Left_415 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_Left_416 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_Left_417 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_Left_418 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_Left_419 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_Left_420 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_Left_421 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_Left_422 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_Left_423 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_Left_424 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_Left_425 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_Left_426 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_Left_427 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_Left_428 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_Left_429 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_Left_430 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_Left_431 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_Left_432 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_Left_433 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_Left_434 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_Left_435 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_Left_436 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_Left_437 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_Left_438 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_Left_439 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_Left_440 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_Left_441 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_Left_442 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_Left_443 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_Left_444 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_Left_445 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_Left_446 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_Left_447 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_Left_448 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_Left_449 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_Left_450 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_Left_451 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_Left_452 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_Left_453 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_Left_454 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_Left_455 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_Left_456 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_Left_457 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_Left_458 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_Left_459 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_Left_460 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_Left_461 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_Left_462 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_Left_463 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_Left_464 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_Left_465 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_Left_466 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_Left_467 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_Left_468 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_Left_469 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_Left_470 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_Left_471 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_Left_472 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_Left_473 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_Left_474 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_Left_475 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_Left_476 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_Left_477 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_Left_478 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_Left_479 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_480 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_481 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1_482 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_483 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_3_484 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_485 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_5_486 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_487 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_7_488 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_489 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_9_490 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_491 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_11_492 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_493 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_494 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_14_495 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_15_496 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_16_497 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_17_498 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_18_499 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_19_500 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_20_501 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_21_502 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_22_503 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_23_504 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_24_505 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_25_506 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_26_507 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_27_508 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_28_509 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_29_510 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_30_511 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_31_512 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_32_513 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_33_514 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_34_515 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_35_516 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_36_517 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_37_518 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_38_519 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_39_520 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_40_521 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_41_522 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_42_523 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_43_524 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_44_525 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_45_526 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_46_527 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_47_528 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_48_529 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_49_530 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_50_531 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_51_532 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_52_533 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_53_534 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_54_535 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_55_536 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_56_537 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_57_538 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_58_539 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_59_540 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_60_541 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_61_542 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_62_543 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_63_544 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_64_545 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_65_546 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_66_547 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_67_548 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_68_549 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_69_550 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_70_551 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_71_552 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_72_553 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_73_554 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_74_555 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_75_556 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_76_557 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_77_558 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_78_559 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_79_560 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_80_561 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_81_562 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_82_563 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_83_564 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_84_565 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_85_566 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_86_567 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_87_568 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_88_569 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_89_570 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_90_571 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_91_572 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_92_573 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_93_574 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_94_575 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_95_576 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_96_577 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_97_578 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_98_579 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_99_580 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_100_581 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_101_582 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_102_583 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_103_584 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_104_585 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_105_586 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_106_587 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_107_588 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_108_589 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_109_590 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_110_591 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_111_592 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_112_593 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_113_594 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_114_595 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_115_596 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_116_597 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_117_598 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_118_599 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_119_600 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_120_601 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_121_602 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_122_603 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_123_604 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_124_605 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_125_606 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_126_607 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_127_608 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_128_609 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_129_610 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_130_611 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_131_612 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_132_613 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_133_614 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_134_615 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_135_616 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_136_617 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_137_618 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_138_619 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_139_620 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_140_621 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_141_622 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_142_623 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_143_624 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_144_625 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_145_626 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_146_627 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_147_628 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_148_629 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_149_630 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_150_631 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_151_632 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_152_633 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_153_634 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_154_635 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_155_636 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_156_637 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_157_638 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_158_639 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_159_640 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_160_641 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_161_642 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_162_643 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_163_644 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_164_645 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_165_646 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_166_647 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_167_648 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_168_649 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_169_650 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_170_651 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_171_652 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_172_653 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_173_654 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_174_655 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_175_656 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_176_657 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_177_658 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_659 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_179_660 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_180_661 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_181_662 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_182_663 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_183_664 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_184_665 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_185_666 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_186_667 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_187_668 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_188_669 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_670 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_190_671 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_191_672 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_192_673 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_193_674 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_194_675 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_195_676 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_196_677 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_197_678 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_198_679 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_199_680 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_200_681 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_201_682 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_202_683 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_203_684 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_204_685 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_205_686 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_206_687 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_207_688 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_208_689 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_209_690 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_210_691 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_211_692 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_212_693 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_213_694 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_214_695 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_215_696 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_216_697 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_217_698 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_218_699 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_219_700 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_220_701 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_221_702 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_222_703 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_223_704 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_224_705 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_225_706 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_226_707 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_227_708 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_228_709 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_229_710 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_230_711 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_231_712 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_232_713 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_233_714 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_234_715 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_235_716 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_236_717 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_237_718 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_238_719 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_239_720 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_239_721 ();
endmodule
